

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
p0avYmdVO1CjpRDP5Bh7BvOEbTLrShAbzJj48OCdmdROF1tR/WnkAB/64d0hrOzRzcSLHtzBC0tK
07WonAQXnMqJrU5Dkow0am9i4vaJ7ptJ//gHTV83ytfBbX7aKpJ0DV04NVhGtIYErVto7dZYBcVg
FfG+/URXXTfe7bLe+YxZA1Vg5RKOU9aihZv+zpadDdqhQrY4J5mJZG9L+F6eYoQg+NMTSXhX+oPL
CDgPCzbgbKZu9BeXKemOgCiiGhmtn6EyB78/HUBc/WAZTfY9mTg9Err1GVDgfFCEXBXHL+lrbZXw
dkUXx0UAXLXmu8yE27+f8jmKiO5qMZ3OkHgjp2PhXr2INZh0TXocuuALIg4+hrP+o8zPjKT+p5bC
I7kFvcB/doQRPvl+WH+23FIk3jdqqcai8KBhr5brT1XofoLpyQfq1lMv7iuNcs3dkpsESgU4+Tdd
2C1Dn1YqW5skqfMWJtZdiwoOrqc5IKV4Php54UFijOrWxSZZ18HAcaL0EU+IKcNGt+aenqanIAEs
oglUshzJVT4YhlQOX+PoeiXU45n9vU18a1R32LKE8axMC/EoOeyKud9efeHBcnwzk87uFWWG7WzI
DGtTXXqN5wWw1tro/TuXCBKfO0cugQRooTbvetUuJTfWAvOJuDa/AbgK6kGXsiIjyAgYzhSSfHqj
Ja2dlFL03DuP1REgOBENl0bP98wIuNHDvPuc9xW1Y6/eX9ZbzlBGdqMohmZaCXj5R1RzlsRn5HNk
tO4wyk/paWOjK0fCrp6eWYK44nuRS8L4+m6k4sPhyPpdWzosn6oslGyitenTlV02RuCWsKggrUNe
MXMX2Kk5YYsrkgs0zxfCWciZNIopMByMisbwvRQUr4nquLSRwqwiU6ROeE4Ex+mu19N07k4kvZQB
u6rMqJBIoTOXnZ3QWcYftXXQHCER3AB7iwAsouw5KxLIX9jZcXRwb9OXggDsVKebgcp/KRqcnMfF
TFGreOkEC4j2yQWRjQuyiCQvC2d7QpDud1KVfcicUheGptR4FNU6LwoOewuPygc2u7lQwcFi0byM
yb3ZKMRS18aSL5jysauLNky+my8HrQo+zHWg0zRoyg7vjH0fnxqpUSSMQRgpPA0o1mTbKaF86Gsi
f82/14dMNG078FBDy5bXEo2Ud1xAW1h8XGY0uL4ZKXE9QZ5u6WAM2A1M38IsyHiK2bjnkNyi3xGF
/EWcYQHZTJhK0a6hqe7IYBhwVGcHsSr0qcOVjnsFZZEZJGgOuS4FgOTTWKXTy6BQPOpxoh77fHsH
2Y76FKF01S/eGMMrmVagXd4MqoUe4oDmmzIm8Zf1TLpY56+sd7CJ19OJqoUGQCjyS+fGjdzdTZs1
wOopzTCRXy0u3C1sXB+5UH7Dqd1jRqoxO06wSsHjcXite0FabqXFS5tc+V8v6Od3Mgimj0a1VgSj
JvjbtT4cjrWodNvRrTjNTp4I+kHVtFhv9SWIUTIvtJfON9C+ohL9sPoFHZticnlfdv2u4/rmS9DU
lJcbvvay8YKcSql4QzWYwGf5F+Vt0M8BZ0UKdDdw9vPl4M6NcXGNF9255twipLV4hkOpCOvyqmh+
jZxy8SgZ3RZfgEkeYm1XyV3xlBNDTB63MBKAiaYM9E1G5JA0mfoUXvWx594Mj7SNM4gG47uLucyB
oRm3YVV1YEoKpIJaSTvtY0C0Z8hQdS0OM6h+Qo+3CBb3DERtie4T8zI+iDpjptu4uoTKX3MeCWWh
Rik6D8DMU+GeWhABuRgL+Wq6udpkLvcCTQWsrc0RbKZziuVyGArCrp1coq7PnVoOA/IYXebaBEeo
vLeIAxUSuEfgcEzdVsMzDTuzzYiufMJcINngJEdTHU02BnZ1eureg2FGdYrm8XNYDsXR2GOfh11G
zY8V+QWuBAddYLUPhgMr0ZgmQkvNroysGMqn5J4l3oniCc9QwXMwu2Y44sK67VoQ0YURrq+vM0+4
2QY+uas/NuND2CUabKQYdTAZD5DW59aW04AbdMZHK61u0FhRPV+v4LpCfAdRqHUvJ9jG+8trjDqV
uiXSAlvNOuQcnLXCTagoUBaTnSM74eBJPxonXSYArVqXxQl2A0v6Fvhm6FQXgmO9fc4Fn+wl2QDz
dzvc/bUfNcDkB3MJ3Mb6r8HChp+GMKOr6XLnbN4BZmgB9fOXHOv+CNDoaKUPVypskWTd+UsHkRIG
GlXQZR1Av2b8YTLPbaUBx6oKHwGGT2uwvR0sDgycqIFqgPg1C4s9OsWv2SCvM3/2bCyGjWtXJ2nm
e+EwqknvrXOIrhdBlRY6f+nbZjbMFHmBgsnNzVwhVAKjRFp4nDkuLSrC3sZcC1a+4aftP/U9itwz
luV+PrEVoIvLXXJGSVsFbgUxZe7Jr1osNleaYBeBzX1mczrxU2KbZWh5gJZx6djQIXMD3YDdQxKh
IFMPw1MxIUqjUUIYySCo+029SlrUMaDUb8vL3PN5eokjHheh+erAldfbCCTBj657TidUWPAqMlpl
iS85xPAsT0RcEvR7frT1sUEiQ71MLJDXjwHokJsLatwAx/gjU9qqkGCFasboyLlEM/Se5zcrFINQ
oJag9A5OhMNazYYf65V9BRw0z8eUFWRcbNV9SRiUC0vsTKr7MWp4LfNsK624Yml6sfbYuO6RBpyv
sUL1c1ZG3HKmYSK8G2FIvPNHhwnwzIYNdL7pBR2Sc7dd7sMZ/p49SKZi5+Ie5KY64ICa8QUqdWNO
jtvBZ3hr1ef7OP2IsauPEzBY5StfrnA2FN2TlThadwmaBqZfC2RiZiGisXI8ogEcDApEf5qBz2W+
NF5MQJ4JsMQ3whfepEEFICVEekS+oumFernFdyvAq2Wv85Kny7nu2W+cCFWOzyqmyZTuEWgtBbcx
kJWJlfDdoc0lphtwBcRyB37hoxfPZhoi/+NFM2TUTGVCOr9I1dIrzFYIHqRzfTrVbD6+kYzGBi7h
vege0uB0ltNi0MlgWxOdHvLu/qs8qFoas1DSTuliLyZpxvxLYRWtZzjTk02g1EXGadFKj8koBgb/
DabNs12QWeZ18qvgnnv5/Q2x0z6fH1CZBbk09nLXJovDdHRKo9Qs6tU/e9N3G88HPutZPoeXiMcM
VjwO9NuPmOReOxivadtyi7eUTc8DGYgRluDgdKTYtqGoa+v4XuiimFsDYMmVV87gPPilsceH6dzQ
SyOgS7ierYRJ9p789rRamzU219mR2Q02T4SsI8LY67uy5q0fn5zkxm31cf0ShXwqm6NMKnTXUsq9
T5YWms31ZCDq+h70lBdXQmKf9805HnGelu8dB5U4A6fCSzgqlth+BZ73a171mCiQ0q4JRwUBhpHe
M8OumWvi/jZ2EJyXMX17D+uYFHXhREOcd7ta0DtSp0LPu2tTzAhASbifQ7EK1YWrajt3ZJry9tAr
Sdmwip99VPwYaa1c2myFWbBSAPgIMjHR91AyIqkqzwlex5P1Sf3i9mHDdshcsAW7xP965l1lJYN+
l2KIvpMp5IsuGEvW+IlsycCvkONs5hH6hO885OvBsw1Jf2uidCpwml7t/zBs2EyrrzlvBbyzlD/Q
vkngED/VQ10akpLkIiwjQ5acej9YNBrJHUw82ixTxg2ovxxu4luKx4dvUo+LUo7wR65zl5gLUGt7
I/ARbYVCVoy0pIAXM7Xonc/jaFdrqOdWIMhdte5QSJT8O7bVEt4Jpn1kyvHeVf0rOHQyjQTz1WBC
x9q0g/rJUfK9a7iH7VtylU28x0fb3CPrfNlAuGXv0Y8UkR5gM99Kq2Jnt4xr+CRX/jDIFYkfeWBD
VCcoTBMsaJMT+9+v9mqmEn84nYmsvuwenf0NavhRBNK5dyuDiXHg2LmwnJQcYPs/DrXYWapacuMK
rR5ddIpFUbSiPkuv1jTnnUx5SfyRXN16jekH0n4yeGA0kiJAUyvDp4YYzS1Uh67Cb1nUqKGvb/2A
Es15+Bd4k8HUeNOcO7S6x/7Paw1wZcbVV5sT9aGjxpP15y0Lmc3X3QJSyEqsHbeiC45JRxT4GdCp
TecIWkA6sgA829LbP/YalvQVmMfkm1vEPbXJLkceSwIzX21EObE61GgIrXLyPW1dTytlc6kN3QIz
JIMpPuCD9JzFKDppRInHErvL0aIVJ/RE7jvrcPC5UePwwG8OlqU+lgtOpkvF8ux+zsjOukirlb6n
Qbpl5WWTRn982HMouBA96gf9FSAZFZnGdUXB2NRsDYi1Xk8pYWSq2IIVpJMKkD55pqNcoi6sKehC
wYFpr2ICvO47p1bnMsJQrSWAasYhiealWT13pzDrIiVkjdeuPAUiScBUKPyf+NZCjVnowu1cRtcM
b98UQQDaRZcKJUCuv/yiyFBVWLnRr5aGI7FeY5zoxqoKMoyuEblNMeveg8SJ6gDqep6PVExJteCf
6D+Ps9Cf/Tmy+1OjzLi6G8GM1fkj/Ohvf2evoWP5Y30hMJ7SPGJSKV7XLxXlHin9lXeqvcIO+AtY
pFSaw8ne9B1QR2C09a/5ujA1blVhBYGfDIVd5njqM3alblcV6eJEbPqmCnsijroeBc5efOVqiabA
yR2nJYaUc+cjNOsxnqXzGrY+iRlPHPFS9kAIPGbD7WtAnPbQpXaGiXW8B198o/92M9x801EyWJPo
NkN3ZRjYEFvNAmxXg9T5GRAbrx4YUuNwqZCOd6G7kadOX/mk2R/BNz/bU8jRuGU7E1sT3T3shEu8
MhtI2l0+cXSAxAmTIan7H5nHGKH+qAOitxkDbDeYjID1z6sa/LESs6vm8Dvxg8P6bTflTfmH+8qw
b1ylyXYFJ/VGE4idGPmpXcN/uCSSyZMYMZSSGhi3tTRG1VQoomMakhLwDwdpqWOK3BYkcrE1VEMg
JymbysRJ9cnDUKXE5h9AN+2E0kYS/yWCg8W5jJC55m5Tv4G7P3oZwXeToS0yFLQARNDgBmPrLVM6
pO815yP3Rx6n659FiF4iv0qrdMsGPVznTf5MC2fsf7AgsDkKsvEGg5ojzBQ55Gaj8IWfxTsdAH4d
W9pVNTRaoe7NvoN/fTGYnC6PjgyuvoYvPbk/YdVNaXgDv4kWGQJakoxGBsutEUZUYQ+srhF5p5jQ
aQY6snjmqBiripjAtO3CVKTeHVawy1TUc2oAiDOezPxasJi8jpoCq6k3UUNXU4hbnyFYmq7catzI
UlxBXky3+pfBpm6fQZQQy6B88nN6Zcp9/NMBJDoXek8lzfvvZKKqVxxdO1mDxRE0Fyg3UVb37jXb
xwbIcJ5MmGQpQ4GIzRiVLV82CQVdc8kgjbMPqEG/P69lOFuX7vvDnjL4C1k0so1/rMcbHkIVnlIj
+0fGnaS51i3pMgTI+dtTmICTncsLVaNRKHAxvyxSHybw8nhulYiBdUaXkE/4xTCM4nHWeLQJXZjb
4dbxNNy9BXUIaaer8JD4KRYtGG6tnmJTWXzoZ+EY1UZ3AgNs0vhw2JiuGRd5Abu9KnFrvqhJXP8h
1hP5OwfGLdEMXGhHM05TgWoYCc9nSpJCJC7ohbohMJl+wheiyDne2ExU4VLPqK0AFYJRAynxeWST
OICXYpWacpvFPbCr1/m7sco425OqmHJpVzlKMhNg4mK0uLQWJ2bqyl3Xw8bN4E3006sp8iPhNJKS
d5pkZuqPcyd/RkoQJWRSbxmQ6QnVK24M6GmgB9BRf+aHSqwXxIelRrTL7zkD8VdivI7tCj8bluHQ
epi882x2uGlLpPQWkIE8TfCSqPkl9VbHT0CVSA51f4bXABOXKIhUpfqbywTUoI1kFuDVR+Jzje7w
TUcfgghPmBb5SQ8JUDrfo/0x6XKrh4ASBtWIjB21S7LDKmnmaCUH0p7HDI8qopQudMD0md66OIPz
KKZiQnvEGILkxHwfg2nHjhPqjHz5DamitMnWabUJDHWlalEpoT84lr0Cf0Xr9uUIb4cCd4hxQtCW
IPcW70k4jLW1Zhk/UF++cq0deZOF/nLX/ROAfHekUdJuL8BRO6h6kQZ2wyX2WmIzH/TP/3E2mobA
t/BwDRbBmLBP9jd3xuKHZUHpGVZNKXyfJoJhnGVg6c1mOHpGlPiCR5lc7841HWf1CMJwbWLjCJJy
CaOJMrSjCFmVtI2tSczDHF/d1iGWQ3332pMaXz8r6Xbn9XG7oXNqZlmLtfsyCDt75sfmgX7OeHhK
c8L6oP0uZtyKyWJgunyJtjy4wCejcduQA2qvfkofIJAEv5kATm+eB+GR5weVzs18tplj124xqvnf
ZcoIorjto8WFaTHt7ehz1u+yvN+sWRckpGfpj/telRK6zJgtLyuk2hu/DqjEF8zC71K3yWnx5+qb
MJoqG/AA8uMn5OGrU5e03G/6zZHrNHLu+qncmkSykrfQTb1iyJni7YLli+TvZkk0RA1TH9H0HPFi
xig7hQblKfIIvfksI/U0L9FL9q9DfbTehd4LEXMcJ/Zfyx97MyJMWkczUcdnWjOv6Bzo6AEcTyjO
kk2NPwFCtBxlpHRtU1WfNv9o1IdzXhi0uxCPwC0CgBTEgOu3vVLnhdmVdrrqbWFBFbIVbg68AX4Z
aFR4ppfgPXTyQBNziXXcmQCX7InO76XkJW0QCyq8DlVhvg8XlB6WhN0LtqidjScwN8kySLvmXlZY
ymkPLdBHUlomA4lkeVqj9WSS5wnb6pHRyBTEqiV1E4mVLTmy2EhJTq1KGiPF8dQMKM3d4s9ZMyTK
ogaqlvEKaEe7fct+zXi8L7Ill4C4mu3+iNDR4zdib+faemecw8Bjw9SsH7XeYj1Qc4Kmbo8lCZOS
qPxGqMQeKx/0KFqmIU/u2bSPO0C702/DKU/FEVFx7qIXzGddljWIFgY2A8bnzEt6Q1PKxHhA5fZQ
3zd0cRRQfXWHJ7zHgyOYWg8dDRn1QMGmVHO639Zz0lcIliOdhQdtoRoHXmMhsuATHkn95HO+rgdF
qeg0rD2WE60nEcNPOAQce11h2Yw8eIVvXZpuSJ2NgybnZjnR6ZYSF85a+6sDI+Ygmbrsikh8N4je
3ccxWdQV5FIIgG8epzAy/ohd3wBVM4v8VSPZwHNWsF/pD7TdqZ8Z476ihIUSzs3m81ct2Gpp4/Yk
uJYSqeABpBln9OcHlmD310ukwO0ba0RTweZ2kWJqCAkUoIVcZh55USxNM0sZATJJWn1SjNll9vam
TNlHgOhTxl/qC8q/BpCLiV3ElWk19/dg7pnRLVq3bIx6loWv8Jb2CxWvLnvCuekTSw6Tkv4FQK3z
VzEAokjTWUmoFb+nsCqV9cpTmykzMgzOxvl06B3c1OfIk6XXGyR8MWC+m8SFoXy5BGZ+dgNf4fpF
EIK6ijEklqSWbUjnl5Fa4xXnmqfZaAxs6j8b33WVuWO66a0FwfbY2l0O/GBXt2V+ca25kes6CrB9
z5lOXbgtNeIybIhW4J+rZ6UyRxOjnxS7TXtjr3tBxvP/FMSq+qlxqUmEjLSQh/b+U5BvlFQsMLWj
NYsp/cOZriWvWMq/ZJr5aVqD+Cu4CpwkGz8SW0HN3OgBCyKZa3ZlyfqhyH5wi4XI8ker7iJccpAt
oI6wNQPDlaqwjFpN1U6ISlwSL64yWa2vJEXf4qqlGm0PCFLVBBe4fY0ARH8n2Si3FJtX82CC3zbN
krk06FKYNKICqLDJLubCuYdb32DGtm2mdYnnDOv4WJBfh1bII1/NGIEN8n9dZf60YhoicvYnBQqb
++RnjcHdyvSdkCK/yFxcEbrrTaeufi5OiN39w0F93kNQieVcNF/qy/d+nNVndUGMnF7jHFWYlxUa
quyvkIzDoGHI48mboOPNk3ys+xVHTfcyThdaO8mwoqm5QPej+Qz4yDzBdB+c68/YwCWmsluUeNjs
QHpQiJHTd3yt0q1sXEX4MjZdQWMcyu93eE14F0sSnZKV8Q0RwC+lLNZYEdYqw8dhsp6FqOpRXnqE
QlySVihU9nGYYnWNkraP8hoB2sskZggAsoxjCbU5Kwb9IxAHSsW9OTlq2rI6ys6dYvPCTuk6LM40
EEmDQyuxnTpPdMrBQ0WcfoCpS5oB7KNXvAfBm3s3GM7g2X9dldMEH49NUMHxcQhfrOwECTMNqo4r
05YFX9+qvQzdQKSf17W0NLy1JZj6CEptiIR2y0M9YvU92b0j8LxynAO5vuPec8u+3Ixvi5AdTQwD
3ZEjMxZkaZre2xGr4W9/o/XZJejCJ1uTsON5cxBkjUpZFiXu9mMRpoF0Svy9j77ECX/OG9whBi+t
APWHIi9Vn/agIddM+fBcmxd5eWTkzHZ9MeozFrtfDKcmxECrxbShDClTYYneUQVdxNJwb7laMlyi
0VqyUrwRAJhtODPnGvZgD1EG3fHPtAoE/BhgpS5F47fBjSodRaD0I2eVeB23uf6hbV/aeCVO6RP/
uFPAU5Y8Y2/gkIikYlyXNl9Tf4/hsIIum1GVTyoFwmiyJqHZqqFtco/2f4iH/1C0R54NyTUF5ijm
4hgwT+Omag4kBZXVH4TZeDL5XpmQde6sYDSqpWHwyf2g5ZLUqbIPUBwrkN63P+grGZq12hu5wgKP
o/gza9RxiDzRXDhPYnRgFB/ZAJxzcT95eCVIHOFvgXbsKiHtKwOFRRx5c/1oijUvz5fMITmA4Rcf
6K7ki8FaGij2VLG7qqrFR72Ewh4xFn57iajKuwVSI77fkfpsRUOHVWxyuliizbUeUWsWa53e3PWi
+Z0vcoWyZQZtjzDkrtMaJdZ02NK05a/1dWA1H2SSOiR4YvA1aoX9ljn+WOEE+25ixPhN9rAbG3Gq
S8VpkrwZm391oPRq8TQJfFJztvj6OJL7gKgyH9+zbyxM2o09BzeWhy68KJlkS6WbCJExkqZeNIqx
fKP5Lu/bJlJ2FoeEvH0qmAdnu4NUjLBCTGscM5bzvaJGdFjQD8/oitlOc/5GXk6RTYr06lCQ0cdh
jCpOtas9oYM5eCqWW1+r2Ro4JDTw2HuBdnSsMc3hHtvJ778XQG/HlP7r4mAwyHbVXf4boJcVdwYX
akK4TWSgtIoNK5sClvYoxLHOM07EUYiPof5OEFSEiDlTJCfZcs+4Jwu5hy/gCebNcbDVxNbkJ92w
xiVEm7EJFaOjXVDUlkDnnyFO/6KLX6d8dhLfkHQjOPRaEJEAqDSn7avilpO68OFn23J2stMYWj3r
DJw5GLH7E3t8zDTmUdR4Sk4R6uTMvEPlCCeuW7GMvm7a+1vmlJ/6UjNaOvoULzlXhoJ/mZSnAACY
zsFy7amzDQa07W1y9P5kt7P+XqvxxPuQuz2IzuFNa8piKf7zkzVPMOoOeS5QYng/ythX9vTFGM+F
PrvugnBu5w2N1DFygzmpD5O000lSqhGYuQxt1s1tZ/i0BbLgFMquGwVhFLVKh6DCWWkvkPNM+qNs
Vk1AL22dKZlT70eT5+HTKF/Z9dptjMLVYu4BVJ//EHG7JpW0fgiWd3NLgiGtS72de0k9UEgKAJO0
zz4S4LGjIDjlP1nyPHXgsVII6FIg3bM+ZP2oKD6TfVQVtQGQJloyoNxhysrmcY6J7q1dxJj8nWoR
hw91W780Gg2AtXPXv2OOpyEW74eKpLb3XW6VL7UeniI4z3lNgKD9uCzmZADS0s59D4LHMaowf28n
fCQNOqODrD+MTxXo+rv0ib9MvxP+CKYK+hScKYELYZhnnKPaj7SHptJ55fBR5BnbfghJ8U8DeHBH
PPPbl1Vilb+1xHBTU+ORiKTPIwDY1qEQA5bOlOgL1J1FLxhb4NalspKLYsVpJGX7WAYiLdjDpRno
SkFCwk1Q1VUCMqv63Y7Dc9HsrxjG6rNBBIZIb/21mG1G0y4WAUjlQsIjuGXDTMoyHhOnpPYlkcXZ
uhL6f+s+DJ6VDCjjVgLzBOiRNjNZKVUXF9EeIB8H1h6M2ovC9SI/plG0xlAgQtOwS3SVSVbTkTi9
SMaVvyf/CtxbpiGJR7OXQex7y7tC0p76Oju+ufn9SvE71dVFBaGhCkz4AOn9Lj7vtBIQFNawwxmv
zRH12dRfgGjc//DwWBGNPXTDz6+1HqpkcgkQ2CkonI9kA/AAkMV5/DZgp0msBAYlZv4RlDKzFTrb
IS4hM1f3LXJcGh63CsI8zn/S1sA00Tgsa/LAz17MMfIO4WKRJrq/8GK0BeyHAMIS6icSCColRykU
qTxh/fiwRtYv7Vm8nJ8MAayKxAlp+iGiwM8PGIXxdjkC4E0hh4pZrqnAxgoynfMnhbZTF7KQhtmW
UH0xz6YE3+1/28FuTlZjotJbKaysYxO3LwFTro92Fq1zXLQA2Ufo4029hes1cTbuKYnbsymtF8eI
i2CR27QieV42aNpqzzQcfKeWpmIOwAupcGm3NBucinx/+HFsZheJDRGbShlFxbK0q8fSsELNpWBF
MtXfWaXZnHbqgBT64lsyo2SFhr9ZBJc5fbZIklb0CHbHa5pvCwNLihnxB4jCIJ+I8WCe/QnftDOa
lCmazhJdu20uctgFaUDTzAsg/zzogvdqZExHIvZX/m7CCCmgxID/jywWNImqmCV35lCuWEJ9rlBp
utGrRvB8YV9yvkhGYIjcNefKSdRk3aekXS5kk6KtOppi8zWlsLuqlQt31oTkwH7WHEQao2X2xbkn
iiK8hDRHy51WKHHZU60ZwPjiwuZ1a4W63cgQiEKu1YnlXAW+VwfIblsot3zKv684CsGWcp2QcYAD
mBkoySXfTtGyzuDQ1bezLGq/ymujLsTXhToc0SVREQjWhhbXts9nHSAaJoggthZH+sCMqOkDRPtm
ZbrH4qj0KxTqMG7XlOAcHjmXSfNaATuDgpT6fD+oyTuurAT3pc6VKZ5izgwFpumxGCf92SONgvF+
I5OsZpXulGh5nfkyQANgfTCWp1Y2XxGCisoMWcXFFbgbyBMsdn9x1ISo+Omcco3KDPLL86eK9/Ib
8XcZePRlMMLPb6utE7LxkYL44mKp23FOg5cb3gbBMDWrJXO7iokdgSMD+dfnqjHMJhp7y2WyNoLR
fGYJNPMqz+ASM7LSC5H5CWagV121ON/mdejqgwXU//WyDuc3ZsjWbIQYzDpFprB4hJc5kKryDf+X
gj7vly8LhYnvuzEW9ZO4IuRhlOlOPwATnsNXJ74k2p/Op4JK6notJXvKqC80T5dDl5hTFhSkmM2w
J/5zT4LilFQzLlYKLCAykaTDX8lrIiVDbGYTLnq3s1o3BvfxtP5E+9io5/4hyreIaivQ64a8E0ed
muQizCrB5ntiYBx0Y3ciO4Qfx/V26kbTl9qIVfStLMPCmXUuqUoje42LRruLDntnVG/mY8DWxS2B
sZwWpckSYrwYjGWUjL8dSMdHjWtWOiyUa5zPKMlBof6Cf0IRzJEjawsApv0Lihi/ZjUpllUwMU5g
x6uJqSIYOSyK0CfBO94SpwhrT1enYRh/Ab8eDbWb0f6tAzo2PvHbZgJS0rBNVlETfiJUzeiAshnJ
5n7rbXe1QfnTXIB16adJCVTAmAfpx6xJKAvWLWSP15zTl/eTTO2y+OuF4C28uk6e/HoysNrsLlsJ
7+mYTI/SBEAmtZTjCpeuj1rlP/7KFq/Xzl1+p5Jl0IPcQaN5rErkNcce02aulsny3xr5vrKCcQux
XM127NoUC80RlPcZO+mFi7UEKlO3lLBF0U8ZuE5JPWcKGvQwZwubs0hTgnF9HCUUCwezC/wOer3z
4aKOjd2ryyJazP118XvwDYeJ9PYaXSTnHgTVVc5H8CeBgIx3oiR8/Mf0wvAti8FAB96ziZlKXjg0
L7lWKowia2mzJJDkDLcLXxgmIIqoaWApGN0gUIBTOorOFGsvN+AW+cvCACwgLwahMaLYBfvL17nY
dZJGJ8CwPZPsyIeHQxGmf0n33KNHcdnREUqOOaYzkRTEudMZLCkCFopupBzMkwdpR8izaNHYSY3y
mX3MfFf/jk66vlcZ4L9919t6xIo2iH99gYAwP/7I8SVBDRGeHYGVQ7BkzQPvDLZxNgSe0BAgnxgp
o/GNJHQcmME40+3fnmgjgB+YuJFiqve8AGxTRtQDgqCWj7EnlAxlHQzzioJ5Ahhp7gknsWojEk3P
RDYEvRGn7hfsryvpyPucNv+pFSyNVoK7QiKJtpk+dVFKcKEpOrXBRk39moGnEdv4zmNa3oieWLTK
RnoIqiI9e9p425WOxobsRJhw8BvGK/2tUen236w1B8/+8yxcw7CNCxE42aeQ64IdbAD8KkaEk87B
EnGpp4C7XM62aI8upTmwRPESpj/qwUlYxP95knofPh+Uso3T9rE0RWqHMeNze+3hVFgD4nCNyqBp
XoJZRhmKtm/QY7F+1bNmx1SYu5zIX/6ic6DNq6ZJ9cMV/ytl+6swNd0kpUMJercdZntzMzruiYSA
TaTi2yvRTdJmJmGCDdJhyx7/13cZKVlN+gvxFNuOidaIYEy0Oy8Nriw2rlT5nb0i3C1/f2DtDq5I
iiS87woXsHoKK2EMRpSBE6yoAcxiKpBPH1RnZnE9mAh68BZJF4ylKV0eM7ugIYJ5+nG+rbHtaQaw
eZNVauJrMWRVa7wZROQsAaQtK6acteqAFXh6d8nU1pdpKjaq34ruarRwWbWjkWhZl0y2xI/zgKnO
/dYWckFPdPGrrzo+uZODd6mNA/qbPbZy4Vf5LQBtao1Zw2zq2RkdXgEFJPrWb6a79J76sKJCWH6x
w0JjatSQqlLPcSM/DlnzrYjxx1X8grt5V/yKLjVL9cjTotdR84krf9+LSG3E7Zlg8Ca+EUNkL9u5
frTqLi+K3Rn5STkfR1D2Yk0vHw38JpR0jo/vVmlZDyMVHqxe8F+Cf4DTAwTdlVfmNeXzzGSxVWHP
BDtC3h6/05XYHkdE92jkrhxZvd6wUB3brf+QNZjfV9CD+FGiryd0sS3H/+hq8rtz/SoALpRUVPo9
dJBjpfP6sp2kNP0HlPfNF4DmukhhxFCALZcPCD/IyPQfhkipuv6xEvDwttwcxOvj+fSZ10paHUCD
K1VasdJkFL4oKoSwXEP/hRDAD3n2dWXNdeyT5e9lnDt4I8EMmA5Urp1PnEstMmsNTSTVYOXeEB6k
fRIydzAX3ec1cucloc694PzorZ5E+/6RJGJCJfMOrg4RdLb9axEhjIk77Z7kK31hp4Uf7hljIwrA
kzJzmWaebKxtCbB8rISdZg7FTRT5qgdY6tv6l/x3eDSGxOHEsot3XclpPWMroXHm7cOQzKFVhwHo
L2ilfgmks6hQ/0nLHAxmIa8HnHGKYL2Uh+Z0wI4dXbdEYivg5HBzkx5miD3uSXk1a4bYGNul+a/W
0cJpvpGq7KfXCxEOw20jvwpT8oteco9cmkitF/3xZLvM33tvzyfqSXPePNovN3kYIXZ7d1/AFUSs
VgmRaYsdjnr5tNJ/UiAuU55JOwgVdm4TA337XLMUG5sTfIB4YGB+2ztvYOvGTUtl+fBah9hg8XsL
aQTaQl0bl1r3ZyZkOm04eCxwR+bJYa5jvMbD1Pq8XwCFEOalW6OMA2DzQemgJMIqOLHN4e94PZSf
NUAj251UU4MxsAGIssYsM0yxifsjPs2X24uoSlKl6SGizg3SmEwy1n3UybY0FpaFOP6oo4Z+gfQd
t0GwaSklpkmYz/vFViVD/feVTqor9BN5L6ravXh0n7QYtov7l6MavnQdCUbYs4x6Opp4q0R/+/Rt
m8UEJ97AC29Q4Kd6EXopt6kNc7IcT6dlN4caurxJeaRWOJ20N93zBaDabBOhMyCMPCbKA069ICTk
Dd6QvaL/+rnWDnFXzuj7NP/b8c1NGkUBIkWHiS9/9Ed+5JpaoL3tW3TmLTE3R9Pl0yfA7Wapjv4x
Ft5pFlAVQ+RzQ+2TYVBXPMFvRLpVIXxzmr2fOcZoZoVYxwQBFw7K1kl3Ee6586/nXEQf8ZBRFemp
FWO0n1QwXR2Q6I2bJxJCslrsi+44/JxnVHOmz2n3W/9iQqGG9+cQUIMjIBTHXOdBQrnkCg880IRw
m7xOxGDyEPVe5/AkyqjdWs00IINEi5nobGLfF5FL+wlwtyLIGKyPxCaCtwEB/thiV6ekv+HaydFI
U3kkN+OCTyE8ErQ4H2aAJoq6e+gd07Eqy+H/zt3e9ABfuxoDswE3PmGcObub+KHgAShroMAlK7S+
FNzA8toGmqHX1yBERiNbVRqahNUO4LNcegH86rl5MseO20z4UE2YIhe/cPCfCeahNVcFjJqnZRgq
+pzKVhAytDYNXuOxQOfr+x62K1nirKbmihcRyZEjOYZc0t9gv6XNc4YR3TE9FF0FoPtk40v296dP
z6ylxL6YgJseFRLuNqjzzuTkNJZFPzlE0bLcpuEj7mnxve4KBiZY0oXuSid8PI91ZaCfdJgIoL5Y
2Nyfsww7wmJuUQ7oyEp/cttUryQtbRN/nhIPzgQWEV8u09yH50eDQj7lIx16qYbaFcvgIvbZnnCr
7t3yNLTZ75UdBTlA/i9+aMrF09Uz/EnBytdznoV4w7rC9SUI4Gptf7hKZS8sOKm7I/n87QnB5tEM
/4w9PlyPZFHx2RoqejxextCw8hg8d0Z7IhXrdl5vzuOHvYrF7yPsRjuJSqCFcY/VgIMYCMG+HhV1
yRUpDzvI6bptcSR9QtVRKuOB4/UjDA9Vri00yXX2lOxEMwoNd4pm8bs7WT0whW3UcGmPvCPo1d+u
im1CBIHNMRYOeHwcTFJRPUK/2uqJr6BhgGSkqOyXQJfFlmtugH7t7T9SwsCHqzPrn0UJcOOAzF0y
2aaVokTFu3LV0NLlcxEIYpUgl3ho5/qlygSM5tLsC2CYPF/AiyKUujFV3SgKi7VTf2Bu71pE/fNg
VhqOZXF7FdYgXUA2R7Nr3Y+185Qe5+/LAz/7QsLjxzezbXqa8zJ1mKRfeHfl7hyJaIvQ9Z9pNHMY
nhmX7oI19tTP+rEvs5ciz5WEqam2RgxPZmQnH3U/i6H86IyoWStIbko+Td81b3x9NCRUZPwYt9j/
8U/khtCUoQaVpPiBHjZoiEZLIQFeh2ElMCGhs5G+2lPV4OgWL6i9Lpj32sqdwxJnQYtzDfOmRJnT
rX55IBUBkG/AZ8483I7SP4hHeFPh+BV2t98Gw3GslBLEnpO9ObLTrbVRvQh2tz0OaQfArGgmuv3U
q6QjuFLg5AQjIwxqdWqbOw4qfFndLdrmaWz3db/ITPw3Z9gtpOvkPbueCKn/xdSmP4IEZSXvz3xB
ixXmCwXPJw2GLOE3WwNwr7eb+ENzTWf3GjAmzJCPdhpssDh21CWnXwlHkcGZxuOEdm75rdIXrNjx
KxUwuv+VzRe0Ac0Ja4CVRJuDLylCph/SWzdI0Zw0LiSINAjwnpqTTBs1CrfgOUF45RwHYf29Z+aj
2otFjsFDwvh5ipx+/Kj7rX8LcBxKriBIFiJWvBu05NBuIMBpYxaSzot/5vblSC9FxwvYNQJkCIGx
WkgXAmj6pbY21L37cGCIs48hiNhl70RMOYS4fHAnPPUdu1+E0zrEoeyesk+mcb+69duxnHvs6x8B
zb+IRO5/1ibIowqvGMqxqk5HmP4efLphg4YrLd9oOim0plj0H45USYQLSqPDb55Z2bYpJv7ER0z7
rIybG6hrP9WYvWFdc/XqHMuM4UOl9Aan7f9WbhHh3aQYIFn8quZg6VjSuGnfQBqZ23i4lBAYYPvg
nxjuEDvvnSljfH1Y7Sb/gI4yFTgKEtltfaVasR6O2d0euCVbHqfzHSj78d/y0R74LQeUlO6Pb/5n
RmCSlU9XCzbaWkp/U85roKY/SaPiXaP31RYzf3M04rsGtLw7c46JeEPz2t4rgFtv+FRaWqDrMJQs
nIDyBMMi5QksDolQ/z+IG+JgZQoTF5iPoEGXBP9ErVggCt4eTNZp3+71WHczU/znj7wZ0hV4+V6a
nZFN9Oz8ErzA1AVwfg8T7Ka22iIMXTA3wjKprGM5fQ5HfS1F1jPhs5nLFOS+VHWEtGjxQxwwoCzE
/bHdOO+udTwtK/OBIR5+euZomzqsg8QDp5ICZ6iCLe3iCoXggY9F4RzU/0EX5QjC+Q3nsTwYjkGU
gBq4GrGlJ7Cjee/Bky4ppLOh28fT9C3mp8mQJWj51kVunjkaJKq8IJaCYXl4ItgkoiK5dloPicrJ
5Eq5MgiuNQqCsYc8HEQGkjopKEtT/UJ8O9ZH+QtsRHG+7W5yCu9zT8GR5bEf96Wsn4+fQqCKytFR
hu5ardnGAhpx6QXzoCXx1z1IpiQ3QkyYc25nlG+3Y1yaEo1QfzMdVrl4041sy3PXWLOBuNpDx0kW
so3B6q05AXhRNqFOhiN8/tfEt5LyuGnO+3BXnk4lGSS7MOBNf0uNaqEms6QBNTAow9TWdT7RZUE0
F7tdYLMIzWCl3BkaiEsBCTL7JuZrRU8DKhaoYY1VDUygFehMKnqd3FMPOImoZIOUEmJaKLx6n5No
AMX+FAzp0VPywlTxR+GSwmg5WkDPLjtYnf2BC60z7CEVFcYf8kSh1wI2n3HNTkOTOaKv+onTd/LZ
vcDPvaQP/aHMxSmRhbE4LBJr5qGHZcMiskD5DZ7eYWZcae+CyZ/8+coMRoLad7h+GvHjT3RtU4fn
NpICVsaSRDIZWS7dJ/CKCYHkxeLwh+BlxH/8LEdpgqp7qLgHL9TSYYyb6/9jATz1LcJP8vQCi0px
ZcsUc9ewwC1F8OBUDTQSLlG/j1GdNZapoin9mGZj7Gaj/juYo+V+pO0npgMTo28q+Ml8gEA3qozn
v878dBjx6tdHyrWDTCiFfm212U75322KGqoK9NVOozkhdG8/Fk0NlwIWC5mC3NAdbfFHG2Ypn08G
cQri4mcobTd/gPoqGxe+6K5Y/LqVHlatPpZ6d0M+ijhy6QqBJJYjJnXzjjP5yQtpx+tELCKY545F
37ebdhjmO2HJ+8CvGJwXXQCE/3JuceSpjfqMs2IRAZXhE67ARJTANUjoYJMG/71XUNGG8KEVSaXw
bIBioF4vOadK/CgAaXneVYrofBxW/5dVWmIzNGQ2coi3q9xZm0ruUrc9+sOeYBKd4Mj4P4TVHp+W
Zcz/xQGdq1AGMcwKWS5G3QB1UgF9MLDLnxFSOEP7an/csW+aqJac8zfzGfeIv7EE8rNfC32wtVCa
2KrLezV2rWp7klzdFCvfkWXIYkyrYDl3ExhXZuCnn4iy9ZI2AVIbGqJOJtR/JXp41te5SlbJLVbf
eNIVJdcmbaoDCXVu6S6uRb74h81731CpSsGzdGkviTNC9IZeu43THZliQMD+Bmcrho9GQsz8QGm8
gvPD3iqpy0Ri9BSAynaUmsWwt8XC9lzo+8+nMz3Xn14m/PdC17gZLeWMcV9inF2s+klg31yLbxXf
Si4zQLvGJcz0Dn/+pzQobZ6ynsAfi/yt1B1vD2wfV+e3zxWG7JdGOUOxiPEXKyXUJPqJW2/z4TQp
M/SNIHa8WAv+muAU4AYBDmm1Q9zIdFKnUK7X7aOdzP4JddCJ7AYG2Ffnoze7eg+BA7F4kzirs3Ys
bRvoK+bC8sbWzDVLSvmtexXOfnkQ21vjrC8FhBv8hYfv05HIr/6ZiBm65MlNsiwPQ80P9elEq24f
5dBZVs1gZHtfJ/MyeZUjGw4vKlWItrqzo3HqTWCv2IJP43qU7LUbGOlFiD5E25Cw2IpxwTK7z1CS
dYdH1wB82af7LW2hsnccgs6FNn8VYO8zKYMt7/bTsmsbSWnNtFuYy2Qnpynk8Mn+qXE0ndPpRY7F
Nkqmya+Su/nrLPUMSi9vvNdNI+OwQxZnj8Nil6zDECNtOyxp4WnsJoLpcprHDPZ6kyuCSd80oy7j
UG6O/x7hjvfzTtTbaV6u3irQ/dPX4TaOmImLcfE6LsH2kodtAEm1/fZGzvEiTdojDDZfkj8Ao3Wi
pLd+TeZyT35nt2HG/XcZQrNJ24d+yWIS+huqvreKe+0+souilqRG6736aBDDoop4+eDHhgrDeoCJ
FPWzKdxB0+MF01qRHG2Sec1tjNlzZ6G/eFFlzPs/wc/luZei6X+QGDYHoARB2JZIG17HZGma/h8l
koUNQMlJgb7nw9UNz9gqrxPulHC2orUkdw1BAzas5SOiP9Yie1EXiSlmGMmHtTghHR8hAHu2rXSy
lcRuwoeq8KMVR9FrGozfDfMwxmp4kunbj6cMflIkcZAlDbZtwmb1UvSKfJomqSgVsJivwBhj6JIR
gLmugwhHVpJ02S95pVjawWlr5q9EJqPQFi7ZUON3hOAOIFD1culnl2Gafoh7HTGjkRFwVYA7xifL
gJlAKcnhfrShunuF3JCONL1gg3qg899NgGTFBEETVZ1/B89vJ/V/FjwZMpdyk207EptkVvtzpFdS
f+odUTzM3wuCf3xsvTjiByVwbG1aSToI99PAOfu0C2oOwXxnUWXiKPtn+au1wYKawqIqWRR1UeQM
pjMh5p+kwaAANE5dYmEDyAV6+jDHoGFgJ9Ts76t7X8a+2e54DBJmk8fNExNsPMkagTVUBpGt100Y
BJoyaMI9sI8A57j1VyzYRyynqHGqumFDXNiKT8+vvuPuVvI8q6S0Y0zNotwN77SyJcCAWU4fZifM
qdsmvQA1eqDBBHSFS2DMZ95Ip+H7kmlcjoZlnONx+8OLWZzvKk9hvzRwSbL3ZHhLIKyUZi4p/D5Z
6tq8H7h1FWib0ylSsrnH1YAKRDzyFEtkCRBC2qYw/LzFtduHC4r5a8Xuk9qLrM16xIHz1GriUqrF
RwWgGPFTo/OYz5TQGTMO8rAfZ+TKcsb/ejz/lptMX9DGk752g9lVaNW9sTXAZVhw7QQ2nqGrxLJO
XVSEABQiA+2eyNoqNtcDtp/Zx3lpAsCqTS0UQUvT6RdvD7pACvg1iuOVkbHvdsaW507CXIi/raSL
DErYEqdR5URBp1vGf6jyJPzL5ami38cUI0Oev6avp/O3CqXqo5kMeieiioLY+oHXCuGsvKBJH37o
eQYaz2BlKtNCKT7E1177I9yZWZMc3qpqbBmepUd0ydkvZAVgmH4QAls+VLyy5kc9PR6QGUAilVFE
WedphG5D06DvTNxQeqssKyCJH6e2Hkgsm01ji5uzOBuuL3ePaYiX59eyhIn9c+MPsdIh0RerdAyD
Ov6uhuX++uXRVOpbCTHjUidpmvQsEK9F1iYYVheIApyBLMWVxzUWXH1wd5bjDZOkHrmbzwPQYreo
Q9iQG4swarPqH6UDebyQOE811gQHHWT+Y790pQdyk4z1Ctd8ua2Xo546ibVzG2nFEwWuUfKgc3d/
EBFWCmOctK/Ibrgm9dQHee+mv73nkDX+8TDO+zt85qNWsL8D+FNEHQfjk6nLfU58lOq4Uf2HG9ep
s+vB7QLO26RYAQxrcLtGmQfdiAaUpsPYCWHpDsFyH0CWVXjVEtvRmanwhyFxs6y6mMNso5R+r/vf
bOO5YGI533ca44ENEuBZKiyiN9HSYrIYrqmRms7bMaRTJD/T3ygi1yaTZC+lKUVG+r1QVQ4REY0F
EM711gmx6d09dXcILQE+hn5OhlDF3mmPsdQzlgHSkijHuOrbyGa2oY58i5tvf5oXQkPFcKlpu17W
gL+cfZOOAQA1Z7BUcR6gqsblBx6BL/PeWufjzAJQKBvSfcaA+NaCerWIwCfcKmNjgAqlxFZaWH0b
Szomf/2saARSLF7L+kIUTwnLdy0p5v9CNnGKYEV1avg4i3i73L9FG2yp60BHfyGHa8HuDBGWcB9K
WzEgE0cC39AoZ1JsvEbFZDLj9x+EqdPLb3+xKXn7MpbEWCZoiVwO19opSBGPTN55GwnL2RJM6pv5
Ukvtq/IJDHFdMrAaTRGSnnD2ott4vlvJ3reuIh6FeAdcujNppQp6I1/uSUI3/GHWTjxUIlT8m6pC
axWmKgfZFJ0mtiZJ50M7z5VDlKfL9VCFKZBPADaM4tD8I3pv1VlKmtZoJvx6uSoQX8M8Uwh7Rgyd
XLdkJ+GSo0uBJwYHG9k5aQ6fxVbQUgpj/ibcP+GV/+ldDZo3h7zP4bhgkOXTgUFPdjkEhCsA9FOj
9nGSF7TND7G52sLmzB5NOGG3cHK9JkUrnfenPkwYC/8WdB+xVRMCbvM/I5W9gdrbTEqlT+78GEiJ
Sr7B1PJkDOhK86N2IuO4Whz35WIkyxZdQsPkJbiNcja2AGdUQitrmCvuKNNrgbtmYrWrJEs5PSPK
BWYU77Vbf3k2+MIsLdwQ5ctfi/vCFK4hsatbvic2F5CxuxzijXQll4/lC2ZkFH0RZQDLTcsvesVY
kOh6fAD8EtoN4RKRa9vZmJUb0DfrJLbvals7uuqf3MKZVJAvnw5l12pImH05DC2JMAIdF8GcJ/Pf
pXhP0izokNfbMydYiGgKrdQb9EVeMocWAyMfP14e6ecGEraci7B2ajQunqZDoN6bj6AiWCkNpLd6
VM39FE4LsRwYBIyuBAJygwocRi9fDrAu6uugcu6vwZIFHqSjvR2LlOt7T+hG767CHjzTBl9icDI6
3tDH+UimrWif8Ba1pVhNdbRYRVb3kE8+1F9IwgivQ9eKqXbjAmgMWVMZRfV/eR+Y7lDNsOCQSOg2
YmUZ7VhrT6RHOPyN/BXh+2COZNgyl58zRpUo4CiC08t6o4N8wYyEDSENTHC5C6WIKOZsj4i/ztc+
z2uQ+1Y7XPoK7BaznO5pn/QuxvnRs2OFjto1ws3Cj1J8vsswOn9TZtpGSnLI2+N3q0d34wgkM7/7
hI4+WxLTAiBLQP13vkLvHZS8u7sftK7buEEslqWT861kjSq4PGIs02XnQ0FLoTOq2d7UreKKrW+i
KrDWo+VDgQJ/Q+PhT8WNZt42Q3FyErnYK5wb5ubTbnYQ9eepNEC9l+QSbPIwXc3iJHPuJnimMNFp
lya/wof4DxqjaeqdlybLGWGt6E3dZyFpZtSiTr2NBeJrtBNGdRxNJbvvM18M0GkNl1sjo3Wo1KKB
HiT7OSRmE/tHRKk7W6epf1dYP4SAoJ/W5DRQFt80091Lhr0IQOh4uqOndqGVQsVs0woauuT0F81F
Te1+IkEO2KM4k1pS3+Ufvr0WHFL7LiUNOWMLOYTU6jh1rhUC4Bcc/Vass81A76qze0AfckhnUlkr
6mZUJu/stRpnVew7rhpWT7OdjB9e9mWxAnShO1UGeUnz8zfTNpfQCn7ZhhhmMmPeZBtXB/CTlWne
RkPn/Ul7qyItAK7Ewn8/kJ4mX+D8Xa+5ur46zPdBmcYX0Duxv5FtsEv58vMaMvd8mRAv3xFBd6D0
BTXal/LJ5Uj4o2qbJEhPSWKNS+ecwt0iCgokRGzAuUy+H4Gy+iW3v8gfqC9WReOaEntR7YBknzz9
Ww++ad7mnTHzM7rB8EyVbqQSRQCafQu9srnpT//aZ02MSvIl9fq6TBCN300DHNYwyv38xzjGLMC5
Nfztw3YClzs2d3bFNyUPzyOxy/WJbbTKoo4N+Qk/DUiZmjWlowxC5rc4GPRv1/S7NhNSSU0qkMhe
D/ATgF/Di7RMvqk5FhcZGFGRp2VBjr2/rPJEinnvS2j1pQRHCViiST/dA0qIfFF/mEA/36k2ojoJ
YAMDDwkbo9N4jauaBeLuhmNAo73BIZHZUiuVFlBifyj2Y6gLE2XOdI5qHyUVlfADMIb07H4BHreN
6dMC1L1yiI+hMU+8HjKoA5+cqDM3zLERaS9frBKhSTmLufeyXg89C6M2pSn/cAwPgOerQSmOOvRF
cjFIU9HgWTd1HmlTXtGRjLgBCBTyg57h149dI6PXfvS4qIOer+8hCV3nKlJvewTJDINsKj4uK1cq
a/R0vLw07MRk5Ruvp8WcymaocL07fnEvXUswobWSmIV285mo2vWPDI4zaFTqbakUFzAiAttvvTc4
cPmKM+ebjRfWLwjQgNdUCuZFXmYPtaCPGLre1RPAznyTtKLvD8GP2X5MOWf4x84l9yB1KkItCDx/
yRaKind2VWICjiBfEhPrchs0qaCvjIkQGndx2j1URL4mmlnCViRm7q/OLTNV21ucnRXKBfxjTdti
lgPNwJyREijuaznADyN+OR46dxJxWGi0DuoYie4H/+ZwRI4gB0Rsu1Y56i5efgcnHMtL92TRF/h8
7Gn2qNYxdOQ4YJLy40272BHKNnbreVqWk0nFc7OQSjC66gRG+xzNYnlxVFG9SvAiO9hKCssAoHXL
dUYdLKBN8nKFwQNC/0qFz3xBTJGTvASGPDpVyjeZChbL24YzlI3DVUSFGI63+fnGeyvMDd1w91FP
u80bu0GAa8mMNA8X9OyAM7++GaEXmwUkElnKI6NgB1IzST2YOlG9Hh3e0Hfn+rf0OtkHwMR4lKw4
N+bgFEFzt20UfZ0Rj+Kc4KjgfLQM840jFMTVymErPuyAVRhMGeWjPclSGROzURGa2InfUKYvdupV
B7Nqn/vX4Zz2g1xuv6t/13XrehsqrsW4uksvvulkyTC6SaPZmfq3/TVcyUBILG1dEWo4sp0cxPL1
HzxVYeFlE96YKjYHuHWCXB8njEuChUXEkrr1b+Iqg3+xGcKf2ePmVluv/Tbf4v15BcOXCv1xonB7
vrA9/HS4SKH6DRZAyBqfT5nmjKJt3MmLyolairwD+s9mWTFuP9UHanw6piBnwnKqPZUuqJhXXMoJ
FMg0Qqbwsly5dCItbZXnK2PxCnWP9KJO7Xtu0aRiOd56pyJ+LkVppeyhmPz1haD2o+UJUTdp6HmC
EU9h3uwvLP1k5d+pvxHHyxQKC0/r0TBpj/kN+hWHmGR+olM9PEN4XBrlzfd1ZiJ7hLatEHWwJiNZ
lUCjsYDMDIQLbzwYbIjG+uUSuk0QwTUEtDSoZ/JygTQYozEDOYuj2B4meVevKjGhCkwWAZtjV5m/
75/4kr3sxpc70V/oxM+QmNRmj/f5Clo0PwfLtmkzVkoX1OTHvfq2g1dr6QkMAbfEKn8HbB1Fy4pI
6H/IQ4zr3HaGELLFKYZ8HOBZu2mHROTpN5D3Kv236M0FoVINqF8q8DMTrleAOxlECd+7yhbN08wk
rn6KIyTCSnWeOy+EJ3uAOMmI+ZWlOIJGfWNgfU080VziJKgCGwKqxUUf9zlS29sDVSwpkI8XN8Zy
nNsSkZF6gcOhPeoaSfagpE6/rj5eFY03hxQLKrKv1DVbbHDch8+h3XnRjoUYmKwq3vC4962krCe4
rMY1fZpTlcoPkInb4b/ksNYyptNnDhdob0uG5uncus6F5/ELR36a+pUF3kZWPww0BHWw5o36oSRt
EYvtW9eWgiYmcepzFcr5rQq0mhD2FAMurVMvMfAfZBV8d30lwsH5d1xnc6tCpulxDLQOLs89Edyf
HOOHLnH27pe6r2YqoC0C+SAcFlovYj74Akm1KeWo/gLlehnOSFPBUZ+TS88xx9xx7KIaNLAJQUMe
LWV4k+8CaWUrEYE/Y86UyUuWvKrhH3ZdKXdxC/uWr2Q9p7FV3dhP66sSI0LyBQ2775HQH0LYVVpJ
gztF1R5inc+Opk9DZgZd7M87nhRtvzAZsk4gAyYdTT15avfpB1EYM4R2E61h7C7+WsPHRyABeuNs
sWwMT334kDufBKO20YQsBSWktq0/8WGJZHBTSmkFawtLSs4FKFWhDJY001ZJ90D0pc2fTCDoNp5s
js8AixMtQa+RIvfawqYXp9YxP6Q37VaVOzIPxk+3KSRjpWcexWUBS8MmR1qsBV5XKv0Q0lhSvUVx
M+6pF5FUVdTevjbb1byhm5PA6MuxHANHV5sn490yzjj5mlT1Xg4FCEgAiXQZ8TV2ut2pWoDlxv6f
sgvSewpXh9379lww/7NY5r4OxRLZ7IVNGlqNLl8eUTeTtaMhXcWjYGL1E1DFUWtDL/YSXjZSvGKF
RvWYXzH2m5e28KNWLRSwMzV0GSRrgXLP19o7ZAkIXd9xgEqtetsePAHuv0AwpUCRrrtRBQ4SJhca
kyyBPaTZAYTsy3+ocywbimHI9ZlUtmqlOvfBx2+/s2R8tDDnpPBq/ktLES/T+zXuw59LVkFclijp
SYEFTMu+6lEyUcGydLohbrcjgrs7dXu/d/rH0SWqBKRuq0njUjAw+HcmQ8SXokQhuY9EqLu97t16
OL4AQa0UMd2vfl5CJvXB3WVVjsl/42QCk2M/JUhQSA2IUnL/nc3nTxBexTcuDAIZXSlH5lYvty4s
ga08TRakrX+6wixBgMVDlVsD8amwc4SN1UNS3yLdwhXnRj5mqs/NQjmZO/X56jvVWqdn1+9lTbMU
TslFYmgqZCyZHVN87VhWEoVsxvdTF9+ZhH2At6wY78DUVsdil41ak6TuETBV5w+ssDrmfSjWcfzL
D3zvmJmMvfuoohOEbfkhwRupZ0e7FkvHGjsmalKcteqyVrqh7w25GdbJYFe9Yted/63C/jc3GLQ8
Z8ajNIpfWdGouYnhBPVFpqFR6Yfd0QloZuT6UDqKMH+DfM2it0bg953psI1YKjlI6iDs29xwErvg
/+7iTMZASRV30sRlDs49whm9pzX0pikC4cGgYa7Aw3qMfrbYdpe96ainuTGLRU2fjzopQ+bodEgr
s7OXFZAECyMgcRKNEmreTzTq3Ls4CMeeeSjkPKfPb8icNaxQg+I6wURxN9aUIgKpOIhte+JoZSSz
5XV3qwRBATe6qgW8e5u7JhIKmt7OGnPaN4f8g6DTwSgn1dixpDAfhHTdP9wGzsL3sIwo4FXJyBvD
GUaczqgvs5cMy1ydkWQsHYHMP8yR/onWJJv2YofYzRY+JW08W/5APxAIt7hSg/s/HLBlkHUxQQ5i
rsegqoZRIGBc2q8ph1/mfq0lNoEZDy84lXW7wd0b6D/HXP9vKwgGwnUp+nX2JePz3jeI3keT21Qq
YgOp9PqKKCyRqrAnsXOaTe+F6la2FN2Eknpx7GtIxjit5KXsMNvVsLOgMZh2gDdZsTQ/k+02ZGxc
2ycSdEgZ1ZAwU+B1saGzGGoSKODZlE7HA+cucLvYeEAEPTbZD25fMRkEDRFXPHN5VFywJJkWxsLt
6u9AbMoi/JCxwkfs0UtWiQiAKlD4NQg8gtY7LRrUEuT0xT5KlC2yEOaYUdKfW/hlMOH/UUqSIOEA
+8XrOLVse6vK2UyzrKgJbB5P2+BfSgLNI4qzrmpTSmQiBxJzsYxG9q+NfCx4f2qTGW5LCJKuZLGb
9Wb3ea0yVoioYliolmPXd7iIxrx4giLIzCKb15EA3DHjy+c2mrpfLsPxtilh7sJQHAXV91FI1u6s
E3UZKmykubejg9e+rMIauvw4VWCwXxClwOfHWfJmV7rbiMZeQx0j1VRD+cCn1/op6IN+edml2Vmu
DboeOqVwuqcKRdP8oxmkaFJu2FjfLL3OKupcsBLtj9/383uiznpT2UX5x/2A90OcS1YYwpIshg20
A/xkEsHaaHmswIelMNn2DopZZSGVM6TZ6/StxJ9R2VtEcvhvkSJhRhwI4TfSG1Yx6t7Uz64VICvR
NauDieTGUSX9HejDDxjBboyWA7qBim6l7IPm82mEddcqsGIfmCdV25Au+EVtSbw9N73Z4l+1fbV6
ukg82xzDCZUGyLbOH0prAddidUcEgDs6BW5nLQvgrQ44vP+D5XdWXrC6DAt673E89fLM1RwKVqio
aY3psVWYav7XyZ9P6NjImL0fhuPT1MIg6Vze38zcE6GHNkKj/weFQxRz4a7xnW2wuqaMJHs144TB
LBtp11PoKDa0C3/3Fvlzt9WHV96xQdzu33tmJZl/RKHCeDuzGrbzT3NrD53rzi8ID676u33AxHln
WaiS5CP8lK4AhqUd0E542QSnHawUUCwvuStWaOAng22gmOv7ueFQlfE01nVv6b/XUEkoRg51NUUk
2drFxRlxqJaiuy/yh1UP8FJRe4q9hyKbrb8jifPqQ1F2FjFKB9OfzGffbx6bDYioRfV3ovX12v69
q859QJhZ4f2NhqIugF4gFll0nor6ySVeSPJ9hLI5dP6g+0R/AUG3LI/PowZguUlIBNuKoPCh7dJ+
jEZNvHdY6WJpJpW4piThpyBcxQJxpMIaUhuV/V5z8o6VAB9AtPVgyYOmNn2yLl7nNhU6Gkb5OvA7
BTGjGWUNeUjYJjNTajIr4LtWGltBgmCPpoFZrZm0kiOucw+Xl+doUHlIqnKwl9y5mpKt6+RmBgYq
ZeIfGgTe9WvGS2XN3kCqy9bvRgTR1PbQaMB6rqLXqGPWmUhJOupcwU/hOE5E2GZM8xJLfEp1gt4f
1W7YrgEcFRpkm+eoV2/4yFS6AaLD7i7F8x06X8oBVP6sUCTPUNOvxJTTDg3jmqDoumUSdbB9I5y7
TO2olmGo76AOquO2yM0EQjzdE9jJw6IDCe+l7ttTaVonP3Qkg64vICks3fnEHojGhP6GTvV0m7/B
ndhwbtLcClcKmVzLIN7I4fb5ja2CMqOeQgGGFKHHh4pWQY2gmEfArtCMucDL4tFubkkYz3TkJ10B
X+8kGcBtaHcWwMPLHOSQo5qoBBJJpySsvmDdUihUmH38QadDoB2m/AfaR2tbhlCnxzluX4hn7zhj
5E9TY5BzeGhhxAVZSJUOXRu67Lh54HeHdRQV4bKpf+qCMVNLugYbEK/pdIwE93mTcT4uu9LyhiMS
xF7yLBm/aBnanEKWwJmTgx19nj0WsfQ+atEiYnQC1enScPN1Ttv8MChDzIflx8/miSo5R2aR3kos
xpnYyw3Ej3Q7UI+rt49LESo97klv6JqXxVv8Am9FPQLr38HPq9JqYQXeQdMELmDQdkPY9yiStuCl
K2ukjH48Nlx+XTtivg6aGnr7HfExemzQMglcJPy8UyoZbr4O9yMhFJ0XifsixUXY2YlLOXkCpv+X
lvrHF1vgNGt7SPQA8UGnXHQqnuARFIYaooV5CBRIIekzUBjTS/Wr/TWBT8XZI9ZX7lO9jc0ZrRgo
5ygCzVGaiPNzbzHl6xpwxUQaEEYay/pp2Df01WwWDyJk9fWwNn19xvtDCylUWgKOjBm6d37Pg9If
Oby7pvfGEg==
`protect end_protected

