

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
M0JX+xmEfjDUfdAboIjZJr6evZsG8ncuVsVwOcxp/oJJ4NoTnSksRxqqZHTGYEwto5mzdDp7XLcC
mxe8WEzcqIbsvsLGomd19iVJe/PzBdKvBscHlRelYnUFBwO+fIp7FXEzj4PVtWOpx3dPbhNwrSEp
6fFDKqHyDzwtfzOF333evmJy3ZKCaqHjc7RS/CofQYE8oqRqKcWbqckMAbrfuvgaY8MI9/6Vj/hk
YR5d121ZqnBOg39utmQxzg24/zhB+qw292WUZxUuQO/MKJTV16anz36vQ2cs7CIgidYWLhxMBDED
e60tWPe3yFYRBZ+fxzkLq4qGTsYIdhg7MezRz8Yq1BBiftpyDVfA+XZzKrMXSYq5kBDzEGFn+7bv
dSt4AcTMiSBGhkJGVjf2/5uhBhH8In5+OPV8XSneKSlP7kTAC8eyqxBghEz6sbrLGaGBSRdHNusj
eK03fazEUA8d74dTKbpHlKeQQlhnxZ4/if8+Na++xso8mIqsY0hZRrtZPgkIqguWUzEApot+4qx1
IT2ed0DNp6x3LsoEFk94kTxPVF2DpDxk9945uVZuurzy4hFkDuOKoJTLt2FXkSM4K2kfbMbr8M/C
tSY65TmWNqK9C/qXAMloSHvQzt39Tn764LZ7HZqmXb5w4nrVMjaDDc1hN+wrwIyjm+QUOE6kXmzE
FFwqKeu4yBsvVFh+3SkuMX03y4Evw9nCL1v8P6U6NBMs+Q+4jAcuO0XVM7okAjxRl3ILGfeJJjC3
6bEPQNxAnfO8ggU4h7Rg6u7bBvAmLCZDNnjZSuFZyupDHCOmj2C4eVsfjApSzGPJBQNCCDCM6GR1
32K7s4RUiK+1YjWcq0/rX2GjdlfaXbaiFGxCYVa5qWskaAne0ylLrxUF8IjuQI/rAVGmWQYFg7uE
Hiopj3Q+6O28bFF4VcGv9ovM+TrzPRg5jOSvhYG/ERPiAB1mIqthBs5Z15XymZNOWPhlFEfG1ITl
VNC4uC4E5uSryxNXTNmWoqScy4w5kKf7JMDZoo2z0yLuDX/RC+j47PumKGi+2k1g1nbU54SLAn5Y
+x2qAlFCHzTxbeuRkhYypl3IyHqG3E3sC6CgPhzwuUKXQlzXhkhE47kU5SgFH7BggLamwYz0GvjN
Qh4mlmcEAzJpWaFYWVKbx8Y7+MyptN2d8z2CoqktxCg8o3KZgoqxoCYHDsAkcCo8SGE8TUfLx0fP
6zvHH1ksQ01QqKnDjqKmpHCh5cEeH5rkkHf9XD9HfvdLDhT9EjSUpPsGkw5tDxTFbyE6qCnaDOmS
/3bMQ3gBYik2i8G1+LdcNzwaQO/XrENU1vMZh2GTj1FR+4Vc3pYs3UoBBfFQAVHgDcI3gIW8380c
0ZfftPlL5I3AKoqHe6aLhR5lI087whlj0SbJ1WrER2KCX4+KFxzPrt7M19W9glQz7xzUU460xmw1
GC5AlLPPLwP702AybtM6RSACgKR6hPb5MGVZA/zHrkLkJwp1JBin7I9rLczT5QR7lSJEZAX2SRLz
+69D9rNDdTH7l1KchGEeWg5oRexKHSs58jjLT7CMEs4HHUxAGWeSULIVjL9s0nJ9O62SXtr/9Hf+
T9qrm4K6ag0HybmesZrTOpAxid/pHm46Bcx/ddorURwkz2IAACEgDPUYXbaa0AdEHsK0kNopPIEv
/rlhwwld8r05BzZNrw2uV8/1rD3EJIi3KwFO6zFAWYtVZHfBh+Bq9Si43lgKJfQlMCudKELrHZDX
5YWjU34+rAEzFGB/86PQgSj+IoxrdORHtsDS/2laUDpO57ZCYsKY3RosxB6u+es0omotjyeN4El+
TbtjcgH7KQer4XmTSZh9I2CM20oRMRbiCwK0D65q0HTvWOp0YqM2mN+zpNzqXPYoOwJpfccPS1wz
RswwhIQTrGfr5M22Uhm9yGAaljL3VQYDc9Wn7j2LxR0KmAymhY+DbKUv4qBEXu1eTa9XyWNhNG30
DYkr6bCxEYg9BRmi6Y76NoEDn3CHcgpFJi09ZZ//6+LZfk9IWC3aqvthvdltFiAhM1ZTGMelTvDM
5YWrn0lV3CmKkUPlcOXnSciBhXiT7QomLUdvTHzb7aVD5+HHtsIFv227R1k8od4ITuwTX1kXhSLX
Dkb0Kmu3W3eGyT0FHDS8qG7RGMGyn1ByxBEdrZK659ew2s/UbiOv6PEY9teyS1Zn6IX1U8D9fomB
IruTxZ9LlYu2vwxTYXU92PivisgVYnYYllJIQ1NYOpNsND2wUPXnyuCiGCqnFZ339Psdm5iwU3pO
ReT+NLZiEby5dI2PwWGlD5zrQCjHHMfkh4Ejl7MQyInJ/ndYPjUXs+DryQP5QQjr557ei2jSZk+v
bdjJSNRhFJSXQ34FmnhNsokwpllGk1mdb4nQczLGdM/EO0w+ljHFXMhvuaiaRDPPaYi2Db/lLO2p
C6FLZroD83vEVhG30qE8ZFIEL8wEn+eEnkiXgvG86WOitLDSPJuw9IjgZbZpF1z9O5HMFxLgEyxJ
wn/TIA0BHIFiVgLQOD0sKAjDSrUyHkUl+aOcif1WbZWc3RblUjHKdB5OL0ilShq3pUL/oSNmuydK
fPA5KvlBLDa49giGNsbrNs9Yeg4pbjZf958jtxdGYLPPNMEnnR/3TMjWqpDMpFAZ8lUbh7JfJU9A
5O7vYtbL6+xG3W/G09AQjb7XqHMivgSLTBpZgsooVVkdJaFz2nom87eLDKjhDUIcG9Kri1vjWFAo
uWjhjaPYuwlPxFbLeql7EYVYNlluXO412GJ7mljJsJJA/IkFz3UTtRbImahvVckyMABgoFXfgAbO
lM80I5gCcoh/KpGsHchBxqt0bfXpiZam5UFok8zd16LROO7Q6gT4AydAa1O3UX32WK03lRgyW7Al
DodKoeSxUdTvZ4wSSEu2RZXwUz6zq+u5By9RQj9QcJC6qHg6v+4ewZ2CVPtWRB+iGMpHkAj5DR6g
MWobQOmFzYxioZpaLa0HXMX7l8QslwNJuEodErEaUJ2WtCWOR/p44UvJCQsyEHJF3QvvTzxlrRmE
/qNRyXI1zsQ/Sllm03B3yR+6px4+mTvktBVB++24kUkiPIOmkAz0QWbDeBSJ6j9T6j4jTXNXYFg6
QgZFHab6Hq/gJCcbYUz3vhqa0tNI43Qo4SC9idNmKtzgcf8KwJvWN5wFHPjLCqXVvVr7rNauVmnA
nHh75oKMFpjl0AouKOJCbMouEaXsUEQS4wr1x2LRmvNA213R4QHHzAffbxKb3NmnBXyf9TAZxXXV
Ezkk6QGErHQrv8FtcylhN7qZ0YPBd0rlpylFx5CY5vvbZhzvTYBKtSubdQcZWOqjtRWHzJPYwm5U
zE1Nm3pshPYs415/iNckzerSwFDvDq7ZwScmJ57+M/mM6Cr3foa8Mm6hczBTNYdCdB2mXGRDrPF3
kNG1zBejlZhYkqGLylqXDlq8U2flBon1fmmg1EYzds1znFx9Gu8SXSA7xkSQtH925SOBswvQajL6
7v7VDNjksK4U9ixuwQ6gKyyEbmrCFw4q749u9bZY0Wi5OzaZiuTQVEuoON5zki8g07yXVttI3zWe
wMzuITFurdsr043aiTyLgctoBgbmZyiMVSgVwzG5sCaT3FaYCxU/Rzw2PdbHsWeSJBwl0CbmeUR1
QkpcltKv5Yaf/8koPJHzhGbQ4lwwBlanwEv/PMDrQfUPdmpmzuCHYm5N4xxtiyaeIdSmcxvquuVQ
ldn998QciPxslaL/T7BhzsM7ZayG7FYgUYht7T/QZ67HIlgshzZaforIzfrdCrYHmcwsjnyo+SJk
1E4AwESCDNF4YbtQt235o0xmDPRRAIycWcsd1AOo4GkP9ZaOoIivDh8bX+/7WYNPE/tDBGFczc43
U31PNYXIgzemXR7+cLqC1TNO//NX/4VQ2LkrGrBoI5ohfniiRvESujV7zMU+JzVbYArabBJ64PDC
tTxaNVXaGcYb8usvjMt4+xsZECBk+YWH01cZdmATIxiebh8HY/CBkzIbzoxFShm8GW4GxlzqQlQN
L+rJlAiaACkrWpWLtGr58mUYVt9lWLca0H4WUMpiakx/vKfjKUUv3PH/kxTs8q8gw2VwturN1Xiv
O6R0pCAs86STIIwRzDIkqIfPusS+NsByCEgP4zdMYJgu5amZVPsM69yaJI24EVulOiXG1ncXaXcO
P13jF5BtcJfO3uIS6/MgwLUKpg8D/ehSe8PMA5/80PLhSm8hK+Gr9Ko5ME+CK38ocL5TkFwrWF2x
GW8Ln5GO/4mHkHCxHLp8z93wSr4vnZo15C37QEzSui2rD+d0UsU6U/rKuKts9OQJWd3YIwX3Kfpa
8CcmTdRCWnb1vPFUjC8jA+2DS2mDcFGmHs8bWOnc+Iz8TQ0QTqW7sR6SQCJtqslRtibunDP2GHKK
4at0sg1+Z6vPf2WFpTXusoAvhj50WXWnpsw/LoLoZJzcYe1xaqD3JEBdBL/THIVo/6UY6stdZ7u5
VJQYb14kYhMJ8E0MwQb2Ohb8OglkAtA69QVZL7zycPKHbRIjmLdLc61A2anBoaobGs1OZlThxCW9
OKHLMlDs1TCTbhFj4eSvgcbxhH+zjEe5H1iiTH1kNgt2BH3xl0TSwbKra9OST3ZWG6kguZ9RBcBY
RmbirW9F28wNIDoQ8I+SPism95DAzjBbduhBzxkuWKU6T94vwNqvgMa0v71NS4DRF7TjlKgTVM/7
R6P5bApr5r0KP+pwWN/H1QWWDSc7aJ1KDIszkS7A7LzEqPlVh36+U3ckEBW3R3jeauWGcEEyzN4H
iq2z1JgbrxxfUl5BXGzHyudlDQ6xnxh+XpVxJMPZvejykUgpu93B6Ltc/zMTWqE/hGPOtuMeJroN
c1MIW6ASSMWlC+Wv0vBY5T+aDy3DsOGt+qS6dZQuStFoDjWCRUwLPNxhbvU4ZkQCEKE7W5kPhv5r
cinYSOAvVISs0KcXoAEHHqMlzOgQP2WyHkXroUERFsyw+zHuTcgiLWS75eiBXAQEhOi2jznPHu7w
qpIra2sq0/phd9R6mVU+0gu/lHzVAoeponGE5MtgsGqEtvkggi7NcFYgeHFinLfmvpAvoLTwN6Uk
97ne6+CwtahrzytdwrGlNiVNIncg2Y4egU4CNah8bdTt1PEVSQ2G35KM/RJeOK1ANx4PARj75yXA
ZfDdo8yA64QL3ZqDw7K5tvj+S4mjaE/bY0L/oMWJAMoIxK8iHM4APbZMm3/j6wACiD55unKj+Xyd
BLCvBTuXMvQI8EMZAyQs6JzfD/76r3f14+qdMcbx3jfeNmWC/ixllVwjxQZLY2p++NoP+8xR29WY
ApT+NF441q9TrHJQ1lb31FhkMytV4WYZ8cdEt75ST6L4zb6OIOy6eckf6sJLLHbaD/zijDb2vE+k
Cy1NhubpnLjbr/pwi5z1Q5Z7TORVzm4GxC040mSdTlVN3hRDgxZTGzji7XEaTdQc6/SqWz6fd6Qi
h3Ea7AqUafy2E/BIRT8m2KZQINKzryg+/0Ec0Uu331y/lliO0WEucBskGe3yo6pTwdT2o0va4tI8
Fh3mz/B2beJqdq3X8EyJrL04u37Gm3aOA+frIwvagnuVSnYAoy/XhhZdA6P/rgIIGTyoOIc1l0cZ
h5M9XvPN4tQEjD2zvIUj7r50hG3uMTu1J5rPvxL+A98KDZBg1qNhKtHfY23FBFBWOicTo8hg6dT/
oStfgHzBwBLTPLqG/1rx4K0CY9kIJCaOeeCHBE4JsZ9MqnPg0duz+tchCKwB6B5GPMeJriZWAoqD
V8/neCs0baZC7abgtr8XUNXf9Re/o6btrhJ6Za8L8Aybqkr0KmsDsB/3JYfVjGwI9dDojwkjqjc5
WxdGiy50rhivrGxeFdCglXOg93FkM+EhAc32wCxE/I0oKETd52nSxBRNJeQt1+IbPiR1EbDhrjow
UOazIOxpdBdJgSFso+1nhbjS/ztAja+4i10eLujRMQpcpFX0Egtuw+tUs4fu7VmxRBkCO1bYO00k
evh/fvx5tpnxpLkDECM7WCtPzkVgUBIp9cfuQo98kE9DR7kuApwm6ZRxxlODa4SStkC4HhL9bM/d
79o2PHxVCD3Fc0WOWgFvgDql9hYSGaKn+yGF1dmCQXrltlFaSe8yWrQF9ZFl0vImy4p+olOgbpWv
Vdu+yfR+sd6o1rKvyxeBoDF/501wWwz45N74p2C3/xNUDTZH8C1V5ZP9WAC3SBQ1wwzeSQoFJDpn
ASyw7Uo3KqwceCZUJVPFAUUE8PYkOypEmI5xN9UzuLGggAEoG4idKLtrm8zpzKSV0w4x13++9wIn
H37w6tNc+2R2dACo5vGnxtIOSnS40rsUGVHFbz9ON/uc778ZfNhXzvHNrVAMCTHDfb5qYQPbkjeG
zt1MmIMM5BIjFdFSgHEJmfVVdiHVkffI8qf8IqNl4gbtWTqgIie9i0YWyy+YE0XDKWKPxWy2GKi3
vVk7EW0tUK48B8JmAqbvR7nl1FKBmK5QzbbhIKO5tV39ZbZgnGFPniJemTgwC5CJ3HfKfpoGj8CN
OkwMS41hRv44HcNecDsGPoW0ONHcwaupiXbBcz5DDCQpnknwLiYBrAI2+Z7cnnRP0RdDk+8jnCt7
KJpI/DhcjU22ev/xGeIPF/RmYt275By9cNB8OwURD2cbqxShzl/3yC7nbXdIQBsRwg5ilAWns3Pd
EyRVkcGcmyQOIhb6TZFhjggSiK1H/y0QhJGqL9LGn5tcJZFYeyYp2pQrnB3YposHgB0dOzndqjSD
kxudkgl4e7+cx7C1VEN9wcGMFJ2dxURVgcMhMe1R7bvKDmjeCPyxZcw5elUwqm31yInrb4Kmtq8t
G9RRFj+ePspHssNJA6tJXA4bve+bMa7NSu8me0FMylm9yQQcOwkQ5R/caYA/VO1JZgwLLn/hzNvZ
u2yo+UHV86S1X4Pz6+I/dw7Y/HnZ4DSUFH2alIEJnFKXEoYO2KwBCGZrVqqPAuieD90accyL/Eos
S+8alTbfokh3llGJL/Oxb/JNQVFTeXxOaVlCxKdOwt51FXGfrIecReA1Sd3QS4CxjuXajcnlFZKy
l3QOaaEMOO92iBRHEolPoZaCjHlSMA+uQNva8LUNz+JtUEQ7+UJpZyf8mqAxaECgQexEXvTYs0/v
+b9AFN94zM+NS+pONCv/E8ApY/1CHY3+Hdqkp8mLzpy7NpwQFfhXqDy7K0PKneDJRftuKlARlqKO
7eaUgEljeHTng8QTkpBG3e7YojsdZTZaO7DVOtfpQkNYRtzcqykaRVBLCSp6gAHcARlfifEda1Bv
v1YCBeLrnrkJa7xlydmwcOh4XEIQCm+HVOZW3NtIz+FjYs2Y9/r91XlirbygKMnDt+S6wXbMxrSm
B4k16yN3LwhT6K0Fmdevw1uIRdxZPDuQuSigucAxswPabzifDuU5H7XzKNTMkxQuABPchdU1a0VR
j/+uRft1cFpQuaN3TVG3+UY2FwM73qgmhSbVS5EOxCyFqgunlc323FVy6Sc5NejIc/K6Yz3K2CKA
iZdrnyU2kpjAQBirIgka6L+fIIa7PT1hcdOe+06ebCtN/MB1coW20dJLLUOzU3/o82qFbCJ/YYfX
GYUDphRgfAgBcjNJG9EbQ2Xh18FFiVgHa7Jd64N3GncPkIkQIfE+laWkw6eod1M+RVpdyVbCdvWI
DN4QpDyjL+CoFEl6M0tiF9J7ADQvyW/zfYD8nHZDZ+rg6l4X/kyB37bt6b4n1GFQHuMbP+mas02b
zJaTlB0AYoZWBSpImhVDitsnZYmDvx3pU+hESu2OSm9BgvXppidFtdVJUmtdzpxcphSRrZWaAr3q
/KUIha1mRDj7zfX4a8cs2VuWoxqv00namg7pRlEhUtf+wbODPyGaasxEK1jodvCzMvt7FteZFO18
a98rjoiJRSHiwy4ueRWN5jKa+XT7LZmH75B9CUArCcg2+70skiIxEd5jE6UcuHrOGeZRdiJk+ocS
1aTTd88DQ2rIAEWLmosCFhzi7FQ7wqZqfGRMMGFjTRtfpsjZRMfkzuQ4M6RoObd5arpdLvwMw7d0
rUvEuQn7faacHxkDkUO9oeDVJrvwg9la0OnhLzzPkAlDTvBKxA5U1zvxCxC49sZDUr/X1+VZNDRY
jyvMlzzDKYhQa2bIdMmbSeYtKTdEuLEMgV17Gn7oijDE1/04tbEe8fxdVxublo8bvlSEroUAhj4Z
4lhu7Keju2TyCWTUXr8zedOjABtx04FpmDr6B9aneOZ6xKWwUpEAu3v5ojqefKeV6uBpx+UuiPWb
HA64TV5VL0O1TkX6eYFhbCIZJYNg3PEbf/vXUz8q6dQTB6sIWckkbX/nD+ztiaB4O4qNM+LXSozR
McMwhy61hNKDTINypswpPEviQzrGwCIoRTYzJzxi6CxeRXT7/RvgpEiwPVSfxuMzlOLGsCqtqMux
DJTBeUnAv7J+96IdRidfLvEdpGhQMOA64TTE55obO0rPyKXGcVJaqDrfH/sw5KvsCmcR0oLLR3ce
c6dtgjR4O9PKGn6WDhjXREA8IKDcvUPqpdCXvHN0nOBl4bbgXigFZWC8d6OtDAaQsnsskZ1iNuy3
Qg3kQ1BLIbOQuoDaWo0c92qyeCzYjznq6TldLM1aM/XvstIHHfKZfyBVqcBsU33zUQPyIQlDAi0h
ahekud8ZeZtgmWAjXDdE5oPialZtBmw1bsYhZTDNEPyo2rbbTEnoQqQAusX7SGwU2c4rrdeWLsp1
d7duaPCgLkqEy6Pvjg4eCGRm5hKrp2g/HL5nXx5XcjzshSLBjQUAEM8TnfkZg4REN6mmxF4joAtf
9LR2bMcynmp55iA+CsNy2g1pjf2TOQlYJUPKPXZcvZp35B96aaoXbbJczXSOh1pcvDXx7LNNyBO/
Dnzf4niWIGy6V+uOfrsNBUdYehv4/FWkvWb08ypfRitBGm5G0/OOCg4MJZWuKH7KsDYyhfmTsEIE
GnkbVcoPwvQBkHW10WLknQiimBDbggNdKi+PDnCutUvqhTe5Rg6pSwWNeN4JX5O/vfRC3sXWHrqD
WzUsZj81jYqD8TBWuswpkWvNS9JJBPDBcwwtkLx493NHYiMXLidGZRbbh91m9Simzw2vn2fAx5bw
f4iXikMH6qDub90ZmcQuP5E7Mf1FGoMGiybGRQy/UL63QlN2o1wQN/fPhIM0/RLNKIVhwo2l1WLA
Fa3vrUe0r1W491Tm5D8Tift4skXwM2LJ5bxEQI2mONlSffbKJz+SrbHTK8N8wN44un+3aD6HddGs
Yd4Twh0LfZ3wSoqOVY5KUgOKq/QB/UpaYFfSZOCX+0/QCNULEXhIEtE1yMKvfKNxodRYY5Uv3Ynw
bMuRnyT64OrfPUi+QaFszYXVAqrAu0WjtaOM6Bs6ERWc1dAPbtbGKFaNHvtQ1ES9rAZt60qLz8lB
Kk/jq2u2JEo1naP6kbmabN9X3PZBt3dcIyr1+KaTI0lHPv/quZxQPNZvrkcwOgeFT+Phxsz2On4r
5NZOyMTTDJRV9UqPTH4Veqo2AeOzuwWUJ71QNHkSZcpOIT4MITtdf++fi60jeqgoUVYDfSMC6Fdo
NAF2WJQHFJRrep5tJOfrqEHeZ39/bWXll+PEgi+a1bzWbdK+D7sNb80LwNDcZmS+b44h5XHrYKAY
mpd1zS4LBY4vsiyq6d4SdbgG0+E1o2tDyxgL9SprG7EjsNNoNqAUk1Eg6CN2SXgEh6T7Ho/rEEvA
NO2/JgiSmnODFA+i8NHxL9+kHpn9bxqcuAQEUUMBXYiGxgRFCTFzor6nIROITbE8f3rkxAiPk2eA
mlytkA9jIHUlHhuL6dxvPQIFoyFhqbWkEspdsxr30XcYDlsKA/cwBTGViVNcb6CAtXQfx0tkhi+E
XmEN4GX4QjiSPahQKkGlxfgFZ0AI21vEdlPbPty+04r/LsOSlNW8Wvwm5uBMehb6ERtC17xXaQb+
1SQtCRa4B0KSTfztWobf1qN2EweCwjcRwstYEDo8NRkbvGN1wan3eKREY+Sq8BvyWgpQEA8IQ1QP
psPo4luMAb4q5NXACQ5quSDaVSAi8neHr1xGXKRIH49RB8mUhlkHhpj3wO0n4BtNcwZOeD8QFZCH
hh3NvUDBpf4uEtqw9qZkDTTMBIiCwt5lf36g3iT4HkzDE2lpZbm0AhmHXdQs7/u2y3K1k75082Pn
8brkYnXcc4SbrqXp4wQzivvBxueF6Vd6SvuQAlhIO4ZAhZtmtFKbkxK1wFtgfmbNw1z/zi8Erii9
fG3fSXBSa2XVQkRrdLC8iCE/X91dYHxbBnLWTLFaN8Gm8idZrJ56rSYokVcLQ54DKah1/nzfywj5
oN1gyiRHwWaauKU+LqMpUkJJTjB7lBscBN+bdzxqCnaggO7lnxjlVz2Jwqnu+hkliKokiufMwRm4
xgqYe0gG3lt0fMq8CuDJ5YE6rzrBUvmhKlIuZSXERJwZJPUxeom1ZIqXI9kyPYJlJ7GQQuJUcncu
n0jwtZ15n0dr/l3woCFDsy84VdFU2BZ8L4oz2QS+CNlkapcaz/RiBJz3r2+kBwORfm/m+oenJsxQ
y2VotcqfqbCYsFunY0kcYfSMgjnm06TMnWyR3O8p43DBOVoxcev5MY3XEQy7H6zTjZqF2ompNNvl
7ktdR2NNGdknN3SN3s9lA5ZzHn7PXOMZKLNQdSXlvbToxS5Z9jWzlEUL9jT9hrm8HTYBZg0TmBIS
ZlMFTXJgrlLiA1+TlHjkInQ2yMzU/NJxHLQcVWIIeUIhT1L1qR8V3vNR1AgHJClAjAlCxxfOiTzh
IrYfo1xy9UCLlsDRAmOF5jT9puYeo75Ymd0CzXqFyfUPdZNGMGFQA0UJzaSDdyFKDIl/DDHJDIne
7xIXGNUL3W3nHKnkR4xF0PhVg+7k/LcuxgeSe5iGU8OqfOtdqwvDu1rl4U1ggYNsoP7BnVxwEKgq
YcEmXB8MqKuZn96DQ6sHQN0ypq6Wq2e4OXPecWj8lnyaLyS3s9SiAMUW7g0a0srdBCR3xj3z3+A2
PnXlRTmAylseuwY9dLn4DRuK9N/BKioHioPD6g0hsDoBkbRuLDuJv+I18Ul6i5hcGhC5XLALX8p7
s3LVUWlUL3XkAJI+INnkVSVTdDP5Z6tLpJ490JNYvYHwVjV0sqvBE84DgfbMlAobNS9+g9xVgm65
HqgTwaL96TanSmUf65NnS7bM5NKMcBNPu6zzlN/vA5aCA0w8Uw9AfiLO64S4ONMBDkbfGYgp7Auh
npVcCd/GaD4xLr8o5jqhOOqyvIFA20oayKiGTlOQ2xxMVoo2YfoW93A1I62OgfFVgl3sS+AfNwBM
7fjolfgfjgYgVh/ooOOU/1h2JXOaWL4GOFnVt/TaqslnUi1Skg5C2skuQsgV+0fapk4ir+J/7s8/
JaTDfxE5P0h6KIQsqHTR+2O05ykF3USfB7lK7KlRcJH7p5awz3XcccfOjZBe9qiNQ+AVcu1MOunI
i4Wj/fLie2VK5yPQyEKwBZwZfatrr6Ci1Bm25zrmwsqJ2tTicBjU3tLLKFNHhC/NoayfyJjVGqG8
1fecV9lG2dxqtCVXtVVGatQq86rvbYUEvqz3YCSlb6LWUlHPKhN/7y3cq9KwMc6D+iTnSEDTR2ec
IwT9+QaK8uapPtca2KVPW0Kna1kysHl+0PwQSF43gOS/F8eLjvADvZQRSHQ4hBlvxvanc6XwsEKR
YdPLUis75nNRDtQ5X7oj3WH5aOaFOfPRQA+a5jlZ8xze5iKwci7PsOaFr70EMZ4yDKczGmkHzJSc
gkB7/Z6dtbLvCa5ohO2YZYWCyFUakBBMl8EB7aEm/7DHDOnv8dxo6gs6vhBN8B0BttyzFl4jn+Cl
69UuIdJMXG0AtLt14bSlG7rzQfgz63qbK99m4Q0wF5zzh3Au+X8Lu+yLb1udTuprTudxh8uZbK8E
nc8/DA9AefNSAbm8JKPN18sUoy3sVxm0YwpCEdDRDoOl7r1fKd7m0EVUlOPfopvvI3W/Ex4oqVdo
XW5dUs2CA9BaXS/nY6800COtJDcXBIvu389WlTgydDWtbQ7DUgpbwUHlA1n6GSmmJvYUid8+Wf2b
r0kaL+wGNor+KfewNIsJ+zc0zya3Xv1bdgr8LAKzVL/ZMRB1Tuw8ElXGcY8rkk2qwJusxCR+v9e6
iz2flkjFyRPCuPKBsn9oOcT6BVDO4P7OX4UIyMnL0eQJ9sefxfSrOrhcv9E12UQLxo+b02z9J/fn
N/Ry83ZS0PS9vIjpItJ1ldOKDKuSqSty3EmU+s8ETxt3k1fiABpZTtsk3RuKS+5BrwELjUbX5l7u
jTqMQSeWD5RooGgUMyGIBQyC/vco5udyoorAbiCqWeMnfyTjHTnV1wab6bwe7ordclK+BMMksiyR
WZMFah5EO3Lq3QgztkTLGkE/zXhnmAROYAVr4meMcTzDsGAbOAbPFWQDxuWXKc9ho+2I0GxtV/0p
FSLsc8Zi6EW5QDl/mx5P4KicFB2YBbRw/io4lBkSZCqIFewJNx5avUGHdmwxppZmh85jonSYBb1E
gvj6o3WSltkAA2VAydhPsMo12xIx+ca7WD8oobCrd2zIIddm9mFGj4WqEaC7Y7mqzs6d8wofcFzR
YtD4QrvH+cYsUWt19vkesCfXwCs+NxyfszVLYVbmPYf6IzW7o6fmR7A4h8M+4D4IR0YzcuC+JjtJ
98qRuaoqrCSaC6lNFh+cYDWh/ulsE8YWAR7LVsruib6TL1DMiSPqnxBh+39B46P1rGfFaO0/8tAR
9zE7UJ7TfW1h5yVt1K3C0C3Y0Bm9wykjHNi4yMnpWguXWJ/6m83dqJ0J31lRy51an0fxOqGtXjsp
S5Dy4cMfGwDdb9YG100t6OeSzjQhKNni6BFn/3+pzc181ukKy4NYBmefkYPM+jadDLEkBrOb8hMG
C1/zSgmiVI3SdzCwGPP9df0NMR4iPBv/9s/B5KU7RBGSoio2gXFmEz7wB13C4iaUurMW+9jtbgv/
fFgG0sXdukjC/k+kP3gxvHd1H+1V1nRKwHenIL12uWZaB9ntKY6lXGXN/dT70fUHX/pfPu6dGmXE
CL03rqKOz/VanfE85W3iEthtCxI7SJ+3SaZzQZahYbRi7LUvh76rzWAa4kMEkyp7UOcXhMRUbfqQ
PujQTJRXvADzRxlWqAyKC7JX4Jm+rtZ4apPT08WjmZg0V9Sb/c7oGqv/TRpoSDABuanpWV+3wlTz
W5L8LIvcfqnOqbwnDsFfySXiBsU/j88R++57W1JCa1YWZxb/YUNs3zh9qfvkE025UOOBNF9iyUhH
wX0O/t9zALd/dQ8zpg+cD5PQ5QvTI0tPPPfxIHUamb0lPzkcSOSKiDJVHR6r/tUJbz3r1+bqgiTD
g8KD5V9AOritCvbu4dsQx4PQLFh6evpaurj/Wh2ZuN8mIjOKnEaxmoERvXBGC446Vn3Y7D7nu0TL
UtRoP5OmzIjUGyjFa0lpd2pxyeRcKGfDjEyHtbPcL/yVuN0C3JWK0myORmIQF41Q4sWWXv0UgnPT
RfiCgJ/HZpxaOOwxGSUwmKvPXWlk9tAJ/gtIvJTcyfFhpWNVb8WKMfd8wotKNOncYTq7zIFe3cux
kqZW4clQwjajJ3WLixCvtD0NReVLBAiPk33HpLovGwVpXvS62bLU8Jz9pWPcQRNVv0cNrasUempJ
Bdystn4ZzXWSCZEtSL0vQiLJS/KYUeGn+2rrAqben9oJ5W6ZvvhuKJLcmnuj683ZxTVQxfCxxK3I
5AiQsjd9U40CON/T6tMBdGH815g5wyYa+4iwcaHybDIoyvVXsggQZbQHjWDP7NT1zyuYU7tT6Vew
kOZ3z62F/CWUQ5R9YTYu8eNk4cIff1YVvmP30tIQkqlwHyHrR5/VYlaafrNryinLwHD0LuDKzuIa
mccOQyevNAlHFwnzCnCfqHQDuoJQVZuY+deiaOTxWDRgwddZGb+67/ijQacpvJKdod+gT8bCxGx+
4ZDAFwWpah2PbIBDU0D3VjpFS9ZpzubEnYrX2pWLMvfIcMqqN72+5Rhhqm6a45O2BEw+q5TQ+RBL
h/CcVxI81FZbOPMlWq0tasW03XQE4whop2pLqjhwr/gvnpYEauRhMcY0x2Wg6UDJ7J2N6nr3bYls
DQXeopOZl7ZW7RBA2ei450mXCx0PA6h/1XVQV5IoK/SQ39V8ugagUwUysLzdYBZsKphUotY1XjC5
jgs4kboZRN296De/X6MgmgFlW+5l1Z+pxXlQjWY77QhUIy14AJT0B9UkYmpU/YEUFGrTIEo3IaEJ
//fGKLxwoQtSqbfC6sXBojbhlYZbTwx1yUll/P428JU/5bj3UathXE9GzqW0qAEAbpT9zfJzs4aN
oD8fnKk4JIX4eyr6wZEyCKaMEBJf3ZiIfiJeNkyXZiAPslzahRRvCou+X6h0tz1jEhbZ7GKwblTZ
qm1P6104rRUEjZSaGZWc0vJ3KPUlkNxTMuAken/NBM/bV3bn95cPAkHpcN8lG/P45c78IGJ3SMbT
lcyGoqzxb2F346As9al16G8K7SZoX4Ie2B4Go8HE/d9kHQ7dDPPOhXhkklGZvYIjaz2gu/SGutiC
APttKH5Tgk7eo1dFL15T/adN5n7OJ2kbDqkQdMsROZOFNjOWbW9anyNIfoXwdlVeCmPiAkITDFDH
MKz01XlNwgNK6cOJw6XbwpE06oEe9GH8aeGUGFAEpIsX/AUwuI4LvzFKnEoM/3FBY5uoSasKpq5P
0UG3eRyRVIDini8rGFs69nVsGrkrMZfgTw3GVYMxf0TOLBcVtDADqlOXmwt2GTIBhSMhClyWXi1B
607hcTBVflnCnZCOq7IuIKuYpV6cFIWfBYtz5hcCjjNl98C6G+30er6yfAyYJ44IvWOZeZtBl9Uz
VpkZzk4hGdQkthUWhRxd2ZFlMLG5fWH97y2TRyemcbjhaTrFgRI1H+h3eTHTEqmiU1Jg38zkJc4L
n0uZSqVg3ONNuf7Eg3OypAhqsLngpJcbzLG8XVQLnDqtaMBlsJOs2EFEkS892xeN/dGKZUsVd5zm
xuMNVOaTCUIFfOfaC7IqD3mfDvSwVXJ5vbgUfDa1udZINcrmRboYuMfZDRIfURm1R+TU9KGMPro8
L4W5/5keMEww8Pr0IdqMMlIyQD3gomfUymPTF3zLVy6MBJFr6+UOjKcaIBRQBqw+6tJ2qniS37Yv
j+zDlpOqthYvXLEHeSUn+4CBqL2MLQXPL3N88MzRSp2AZGJL78KZYHg5clKugKBsL5dKI/vJnL/L
0mqCmgf19DywsEA2qWf9jmodV2p67L8BRt8ngcLUXquzBMlfaoJgHsq6OqbsWO9iMfkx5SPFBVOy
a7EMrJg+uQk37Q1lJlF23cMrtF3AzMwzMZKu/QwAcTJewauf8ogFrVHFLV+5Ngt78M6D9vdhl9B0
OOezon4twPCaYZQCq7RJ3SovC+udjCv+2L3fzQUdbUti3O2OVLzkkEiHmxYGKeS2jWCZ/bjptDcK
eB2n7Wp4ZX3ARwgWf+GSB7xs5sF6fXK7F0Nr0idbCozTCCFeI5GiJkD+d9msLq+ydoR9SJOtYFb0
yN4c00XbVqllokMCL47rz8kLvKTlpPoBDxAlYK40zP+eA5H5Eajl0kAFzX7k6EwXkvowCJ5JIEZz
cSOO42KiRfG7pd1DUysShKDaQgRFHlBZpJO7lDKGXCv8a8xsAN/zG6rE0hplcfFWLahfpuQ+TfFh
Gmv1MGZGXKQgBGLtfzjT8D/m8vaCjWeJuzqCNfPwCK6GasWeJiLw96yaj4fig6ARNMYkQd2Gfemu
HqBe7q2yXu/JH+xuS3voE5vxinjC0gcVMhrpt/GbZC3eFitoO28jr6BgCuuiKQ3eDZMkUirdICL1
ttTxVXQ8Iy1Md/RyEsEoXMEb3PmLiRLiPOalNB8gXYFfINVLKFdLc7u7yrW/YkQ7Cb7huW7STA5e
GorSB8zMhnTELJnDZCcihew+4IpBWQgRALNxQM1IjNjiHgNCSGa3i/hAQC8R03BNhUSb0nxj5wgv
ztJG/4XGW3SMnyWNYmATrktPSReFXwZGbkYY1QrHKNVdnP44wZtzToe495R1kB/pIuLO2sf21dYN
hE120OQDkS1I/rXidkS4ZydzeXsu+bEBDQXufQ2pUr41sivr3txzxjyrzpmFXm2V68V9jcfxJ64n
MtAWxegqRdx0voc2KI+SjiBKoxLkbuwmlGS1Mv2Pkqb8VwMt98/7+UtRPv80e3arRwHLBoLFOM4z
3aApbIyZF0uqkGbQk3vySc5EfOT5KKtgeuujP5QAgFHqI9+JHtMOmSX3S6ZXfOPGb1l5PpFDZsFh
SVJh4CkxflfYz659+ipXhSA2ymus/EyV4ZOEx4g3mBsq5ifQpmtyI8jAJ3ryuyLHYuHLvtZq5MXI
JLJUMeMU89xZkhJexZ2QcPUlfZ5ALwSFF+4tmwWLoWRMm3X20KT3Yaz/AtBvn0i9CWbC3XuAzrfP
s0aYC2xguZKONRAEVsa/KAYW34F/kiC5wvWK0so5Pgv11B55mXqeJ0dlDu0ju0JN1t1/mKfotOeG
pO0nry/4y/IDFnQjCZld3LintFFmerBppEF8gG4pN610T39o8IctGwetnl8pelnOBgNQua81LiFI
GlyjO1kkjqjfVFL5fnwo7NPPfdVlL0TdTUTY1gsIkRDlhfMwpHZYRrZ1AdljEchG3LahjuCMZ/vF
sewkFC21bLmC88XP3EOKtgzmhcQmZ9POOoIzDyX2HK7iXsxUMJvdGrABVAEUSXha4NsEas3116BF
LhP/2EFUTam/aXBvHhXogkOt2/W3JRKJQBEy2cR9/82nZn8BMVw22cN/BAFqXOa49Df2+vvHZEMM
NaVe6NsUO4Z52VKRkaby20mHs0vIUt1JewnFfi90qVGvZwtXhOeDBMN/3ike818Q8v7Vl7KfOtjO
82OkbL54O9/wG2iYM4/7sqvDz356bTmGSEKqD282IMtuS0w6d2riawFAyWM3ARSIYi0ocm/O03pQ
6T8ofuwNhRueRWh/TVMssUtzbB/WbnfW/7g3t0yvK5H/k/5U14FenFjGuJ6P+FEn/+7lD+JlNvV9
qYsIPtphPtLBsxqCzOSmbudt6m/SRLg4yiGWCQN5USSUpwE1VtVwFLdxEsCPuJmIar2Gmf3YERgQ
jygFqhFQ/CWUoTrPNNUvNqds7d8lg2z7PRXCF1MFGeVQGqe0P2trrQOza/UOkHitgPD0gqQsqhY4
zGHQY8ZHjdQwonFrRZlJ1Ta2FMkW26PUteguVRlIflNZUI3oAbDDxc5ZDdH6o3CIa9MTW4kcC9XK
5YbFwhvZ68Fr034a88TUavsR8MGz4vFTFMGc4sIlZ/IrDaFcNq+o1m08NkUqO9sywEJruLhdphs2
BYyXF3yitBt3tEP74RnBCJaX1RO3LQD3eDIRQYN/cAeUmJeW80KuA/4mOLca86pOlhzz0yogxCMo
Y7wU2rbjnbSay4+ea72ZpgIoi9eQoKKj9kRZqXhRpypT+A6B3hKcDoYp2YWAxa3Ki5lNi4GN5tHl
vTS/H3Lrc1t3sQ8IPMcUB8U28Gk/IzSwZN42WsxGWklfdVEiS2OFM5UsHu8R7mGaApolKzc/OdU/
lGyHz7TZH5Wj+uDlBfQAUa4nsa9uRzi4tqT9ItGFmuzaxMXqcho9cu1yfFwV8B3CLKK9WtM1A0VT
7HNjBGuA9dkSXtqCh6aZSKZ6WHFfoMiHAXn56QP/jZ445w7oKCMkqfsVsPG6FZHosDLOFrVsKTg2
MLYdolCGo0LxjN57CrUleiOhAs8EROLo41JmRr6MIkzg5qNYvQ6t/Hgb5JiKBAwUtNrNL7oiqFbR
lj+oUyE5yFkg0EHmb42cfwyD1LgVKRirCph0LL+RuU06LT9n5W4y4FR0ERLSt9LRd5EwxNMcSwaa
5l7GHtx04b8bZmKWUPaF0ceQ90NB07j+V0JuGnOk7t0NyKS0ah17vvv50HQEpLG5nXDtF83daNbL
V/IT5qmaXsphm5AiWSXkClxbWfqQqb1DNpT/0kuhTr+ULAtZOUAajWAhKkTnOfGqKx2sG0UnQS/i
y9QMdAploNDa7y8PCCYDubnDu2o9QjYe/vcczZf1cRZR1e1pcw3rQxiYaSjzsLLkrKNS9rT04WVY
6rxjUFwk4FbaR5nuiEIDfXl1LNxk7XmopJ57cgPWYERCCbyyTFKanqf2PV2Vvm3IwSS6/A3XvH4g
rW/h4p5Paea3F5KU4RbZvPs3xH8HV5maXWB+Otv/2USBIlfdqqKfGAia3lLVDEaaek+ddqazO24W
mQcLGxTLgaAqWM1Yk5IwjYBuOJ2DPpt36qBoKP1luB16FQ41rzccSQ2SVKjIDNL8F2SzdRi/FyeT
hWIAd1BnG96IQdWA51tt6j9jLAh9dm/wxKRUt63c8RONvGRR62QztcyXOjPZru8xbBpQLLo/uRya
Wwx3XbkmlJ8zxckh8gOW+/nUKGlrbRWQs52AZHGMimgATOkj6vlV4mdGOnsLjGpTb54heI07hPNb
+H/UzX88nfnnb1/nSSp2TMzsPlB1g6E+bqzWs0shgfCtpSFTTTIWXkyWS/3+5r1nMyVNv7cb2Xgh
RaR6GQtgnrm8AgbkQBJzNIar0Ax/JPNXShRObw/N6bnG20w/Kf5JYfLL6rKdJY75VL1hV/yn8D7y
9W4NIMVz+h+LKaO5HDl3c11s0FqPFa74eD+8llMJ6cjH+8GhMdqilipti6R1p2AmicOv62dTSfeF
zNkglf4O7EhJWDYllkx9v4lUggBvZ+J0/IUgvTuuMnls7GPKXghvQfYjlhau+ufsSfPMZUgPIRNt
evX8ORevmNpE0WS7coBX2RsEMyqqHDwDXZXEBRBs1cBzmsHRIg9drVPDa62p+6KlwHNpVRP6B7iX
Tl4RjAVJV/cZwjYReZqNZ3huUTEoPa03NPP9f0w/1YVNClOgHmYUkZBz7wEjfGzYMve/Q4s9+WlV
5qbypfWJmmX8wan0jkoQgQqnLHGEXlXdY2/Cdo/QP3wlPd7d8Nt6OPXtm44PNJ/phVDdG6DGEP/o
dj0Tia0bVUHzWgfy09BohZ3zqjVb17GcLIHL9/Mau4OIVnkCL0OlsyqaGuVcVhKvDNVnOeebIE2F
IKpbroRdkNVTVKJsVH9ZkVXqWxmigwz6KzMu8CDyygI1/w9Wf+Zcz6aEiiGPZOcJw80zRxqwBTdu
YGsqQzCMMrCpJHNIEoDRl28PcIpKYH5oDaMdjModPeEL/MNZue2l1vYFjZPOLnBfMmgzInXhJr9i
UK7Na8waHbALY7a8as1WGgu1nSkYdUo3NVI/yYa8y8ZqUu5GvK9nWt3SDR7G4TkbeldcAKPTP1Bt
/gZDUqUvkGnLUUde2y0DUssOv0gwEy89pQHKSiX3XWx7VHyIOPP2L51NzImDB1bfTM2j6toO0gIJ
s8zILGcMJkHDwPWWuYnkBGop+D0W+7UaTufhwUF8a7U5F8pVnHTvobM7RBenysshw1XmP9d/w3sb
+EeoNBj4jrazLLxYgzZdVEABkQrnooAkZqD840YPBKH3N3A1J42wnneBGMh11VBw7u3BqhN/SBuv
T7VZugPmu3eBQgHL/cEN0lK3wXSBXWg95lIpbODNpmS8RvIZ7IHQ2c2mRKkhB/u/Mde8Ld/Y13js
NvSPVYxGrm7OEnsKQ5QuhRpXFQ5s3yw4WEiTYfCIbrp5Dw1Nsbb95BQx7+VRSN7EEWICe91/STUn
QHHRs0Yf6kzYhSD9iNf9Fjaq01R9eufHIzCF9n1fPvJlVUFJB8FUDAusMYxQhMj47JE5OBBj4qv6
7lcAGMMYaK/9rKL1Iz3ZO2ROIVrZHVLMbiaHVG3zN/oVxy0BKO6trmrxIOaIOn08g3jI0Wmk+XrR
Wf3BDKuQUIcMxya6CYjhJg4Wm+y1VDv/zW9UPDrLT2hAWSWfUz8TMyaSY+u5Y2y3qMZKTVH2e7sF
AThhoPJeVQA44xnSjaUEMqvGJcz0tcVL3a1uGpAxmCJtTKw6+zjFP2B+2z+vR8cd+xjmSfQtE/YM
jOr6UuUT2Iz0DimL8y9qMvmzr4G8T3V8K//ShwEUvI2Ws4eG3XrAk1rdpYJCR3bvkRGg8sz6IJ1A
ZxOQtX2eedpDWE+NEW4W3DpFH3OklVSuZG++ExxZpzMimJnjyEoO0MzOtqNa6uHd5wFumipl1z8a
J5YJ8HqvlJGhImgdelLtk7/RJCGLZ1zLWu8CyHdv0tvK7HT2sb3U/xGnhSB9DSS8kOx1PNzI/sgB
3WquxWK7KRfe/381u1fB1Vu366a8EYDzY4UiwkxFH+icFARfintjYvznUYrO9XE/15C5BU/bHHww
kJba56sDvAamw2uX9GtVvs18RcLvAeGHpGBrkURm/7aTK7uddAjsb8UHMAaFMiahNX6F5cNQCehe
QD5fK/+AnCdhir3kN7vbqBLx/OL8pWiMeEL5h3ba2F3GWHf61VJ6jXwyHb9n2RaCyJwp0wvkJAoz
IWV5gRu7JMt5Eu1Sxjo2IPIFi7Ke6cN4IZEjtIedUJ+CFOseJ0K/VKLEqOy9o+tXExvrBkmsIIkD
zh665pJpoWIP9oHnBW4lRmXy4WBk5SAI0+DNUkEjRA+I9PvXqj1ND1oDFW+HHNkIxD0jvM0iocJG
v4DlcfOYQrbh+5PR0kUKkEbJrgSwMc4uUpIyMT8vVOw/4G65E+uyvmq9M6VBjhDKxfd0uwsSDoo2
OI6c/T9TiHdhiEkYSpDd4m3YI071pD8pJGsb+Q0PAk6VJcnBFZw3NFZLPMWmobOXxiRrAQdJ0jTS
zch068lbzHaL7sb9AOhizyOREQST7Qti7gjRCcFMLJ64SSE01O3KbPpuscVP6cqqHLX2xzQ5jMSd
bF23dHdWtgtaEdzjvSbJh+JP+lIBT5e9jA1a3GffrEwVSHRqbRZmAU9TJXKv1mC6BGZHAUb2YJlV
D7mconByKQEMrOTC1S1au4h3jsiLDMmCqwovhHkoUh0KUfOqoD6YjuLiyOhIjWjKeYMg9sVQ2JFz
qCyVFBKNuCkC6wpAUo/Zac0A4lstFBYPh1A6TBu7WzmUYI0i5+uitpEcOygJ0aVi5iFK5DYPhFZ8
l9RKtVubpLe13cxznyctugt/vZeTnQlJYvn2SC5bICOgNYXznRyGBpV4lW1LNWl3p7HX2TkStAK3
D+iegUqH7EiU4z9hK5n6EjKvksNnt4nHaJcGCSy7SsvuIdcW6llvDFIMM8+aiOuy6So4b+NzBznV
63e9tk/QgFRQozZdhUWY7y+OWXmIbK+nAGdlp2XlrjIQnd2g5+XLGPKO7SghDQV0DVUheKNACFNd
qeuCgXDH5IbjxPYO/g/CtvP5VpV4f/fdJ+KLNvXBieCRDIKsAm+yCG/V/peIvpIUGihErwNoAkmQ
YHjpsFjl1MlDVv0xHfPht79z97R+w7gzhNCfX/Cfg9wr55gBiBe7Tb8LYFGavGxBLMcnDUfIE0HJ
TzDqOejPkAwiWuVTdm5RughtH1/7mUomOh7n4FvUwZbnnRf9uZodLryYuD64qkTaOWCWw0ZImQCY
izdeX+VP0cM2wYMd/axoUpkvGdpfr9kVbgYgizhxr4R1CVvBgeZieAMQEzAxay9fmhbvq6cKnlau
Ah36qwqkZJJ/wCQPlNYVXoci1xjkr3H5QQCzjYSESMR4oP4VbfpO1kS5z0Hp3RFq82gFto0LRDA/
wbs80XqvsiZgRThwEoxji4hSm42h4q7oBmgp3qy0PXwz9/W4LiUdeciz72rl7t7Jr+1zMIYq/Eph
JfjRwuh8ZwJ3JwtgENXTQxRYhO9Jy+Xxk/g5zW3CWXyBWNx5s1RK1AG79PSE7Smv286nal2JsGPu
aNRIs7qKpjvrJdaIEmPhGzl4CROgNfh0NKyonyBUxr+kgZOL8HWvYsKJQx054O6xerj3yzmyMFgp
uI57pqPIJZcSC9FJ19fR+4sSPsnEpu9vEZtV6WhA26flXosWp2iI/wfWQ2TzWVLyzIGUvK1+4GbI
M+tPvAmBRprIU+Wd7Hvmw/mx4Xym2ByrbuavCAT47XEwvEQ3/QByLKocfW8YSxKwmML4hsjeeLw1
DQRXOUWzgcC2A2BD9E6WIwMIfdXDgc4jx1KX0+HchVd7fNORgse0/xTvOB20ifDIbxHPFG/bF6gG
VUWdqXlUP4vgwiTLld6hpI2YXzZ5hvnL9+jPAsYMw6n4NAxWtCGCXQUY6xMGmvSVabGAQ63scMEr
KqRhY8ePhU7QtEpkaJR6jvUMf0xRm3l2CuWSPG5DgnnF8aXYmtFT1gTqvvDdX0I7E2xIImHoNntR
5M6mAsoboLTg0wSy1lx7w1VotD32osrzSlsC9bnFAeyI8alZQ9aAukx011JXwGXb9VALRTJOG4Hn
FprXSa2Ygk/XNcbnRQzw4qDtEdfmkdqbKUx1/ms7KFyePQWDVwd0cpwfTMhIVfln8LtNR8GOPtyi
n0Fg2ZAQ8F60Vb8Qj4a5IfFjWAVStic/asqooWtOs/bnEueKFm6gLO2dHNic+3nrYErVj2YPoupn
nh//BiUrfPaGL7YITEoqm/B8jXqJleQ3Ldrfon9as1tNSYudJAzr5PAW4mPEx0MCl+MZXAPu3sXE
8993KYJRliir9PPGMJ3+E5/EAKK/OAYJgrbf22swYBg3Dn6kaMt6nge7Zr4TDYyhytv19Dep9nuW
65CRoPiycyIDTJi7nt7x9kj5rvGKk+CH5xLItKsIp5alJFLUN3YTeVpuIrPzqBl2rZJwoLkRPVeq
6irdgCL3SmFby3PfuDWstpp/063OLUhXPlwmYyoMDuvri83i2e4TpoFAnBCvOGieZTT0Ivd+p225
A86dd0NucTxneBLYyPYo0UaSW676YjGUBUtpqsn2ctig983nE3EwrA3y4JkJV139DElirxQDEDP1
sBm5QZVsnDpDDXKxGXb7RolNQNedVoyy8lfC0lKMximcygRzFLUc8j9YgTt6/AffOPVrNqxmox7Z
y4m7svwXib53mEAvO5ILphw8Zl9+GAK8P3hICg0VFetrCbr2029e5mbeQMKhYfmaTkKvYE5TIhER
eUSbZ6vfe6fMWK+O2TtnBVsEcR/fHNMWdlsCL1CIR0BDUdFa/JIBB1ttX8RBP0LkYf43ScrNE0hR
/pJJuCNb2NpYdSVjZsYl+9YzxhVTSh+MBq98SeGav3Ra1foLGadL8qbBof6bxDiuqLHs1sEpIDLF
WgQ9QAKrWKYQvkdgNTMPCoa1vmbFwnz95CTLs9l+85GiScTPszKJuk+Ydu687guDCAX12wEFnrxd
1xkaWD3cFAavcY9GgC+SF0Su3S1jDL/PcjpkkqH+UwNoy5kyGAar6Ae8U46d2kybqN0ynEsW947s
oyDS9a5xio4I5gYLrzZj+5+XsI/HupDWuEritnmRoCVN++1WkANrz5tHgps1sZZE5b9OC98j0hyh
aFUhGQI5bzQimNsfLHpihFZQT4ULUQOxYWsoIC3PWziAUH8meuUWUTuIO3+9N4sS4+t75l5akUxr
n5L1VkyzwO3lvFdEGBwffLxLJimhTw3Iw+9pI03Y8sJpyj3bL1YIL0HnZ7Jq2v3CXz4ksZ4WHjTz
4UfmMJWOaahOKujAUluGKghOdN5ACscgJwfYw1/UWmmhAIfCghRIdxmnaGqAkcnIzZZJS3ijwB7/
xcjRqN50eaD88aR7vwT/nkF7Ce4ktnCRsGbCyffE2331LlbasnXUNgqMNlsOGz1v8hGsLfZdXBTM
4k5QhJnkrg0GVWbakhUbVVPqXp8RW+iQX2epjcKIpANON6vBSeVGb7RdjH16wj9FIv9UWnBWTqEH
F1gUoYtbhwtXkMqEB78rdo5bqChUI5FgSSKhqEMt+NIsN03VqjMH5IFq8w5q+pZ6zpuBgZiUL3ez
TKlZLq48Pjrojlwr3LLnLxm7ijy7/K11O9BGbqnKV2g/MxxKDlTQ75TW6PZHkkK82apHlf4JkaJE
llYRircTgg+crOxU7fS8EFNfZG/L3qTuGAGrVjJvNjLLAJQyHbyXgDqbLoAjznoKeswXOZ5CKAFn
FJEyxezHLAnKH0yFYcIHitXTy3JzsSZVVhajEhTfHU+FXvnA72CgeiIcjuh71HdyJbwGnwX4tfqR
TbaexVY5b8ip6NHPoy4NCcv9WREwgm+S/MZM+4Marqrq2VySqatdGPfu1NMdNdbLMC6w+1db3eBa
WbnicHEIcY4S2Z/SQLdoRLY5sn90pMi///hO4Y5KmqFgNYXr7wJMGkHtKgx0uuN0I+oezrAlAD2c
gk7cLoCRy7MvNrFiMu3LsoBtBeFPR3zr7mXUp+TvTHEhn92/tBNqpYHLGJ0LpmD9DrEwuuBVh4y0
0uYgZUqsHPo8wprOjzUPQ8lk5hrdogGG7psjZvWzFMoLi0nWOLMKE/vEzx4eWGeBvNkYiDKIX6l3
A7A1RvG/PpjBd6X5KI4mx4JHb8VU1sSLdZoALhggQVAG+2asN46SFzuSVdnfb99Rup2lqnuYvEL4
oXycksFkMfJ7Q9F1gAxtsGPxiHiS7hU9ongqsy5j9i6+wl3+uP1P20wuExviyG+eZy48fcjUAlF9
U0uDx4gPshOnIdP7xu/VjbLaKlfArbijBaVYLSZnNaaZEEGP/BgmEqAJ9SfRpJBP3f0vTWQvGJVa
U1KXLL+bMHttd1tA/RnJu+8xBSs0HGxfVxkBRk1uloCymUvYeJiy4D5VXbA8CDti6uZUGnqK+B4K
wJlim510H1oUn2l7vtJEIZSBzY/4nUh/xhCJs27X4bh2HNwfP4K/4GbgLPD/TLJuFmZAtwVqvCRE
5oTOhqP+kpGFekpJRsbujhD+AzaF3nAbXqzsVkQpB8DXDaO2Wn+uzlJdetdbPFIIS2D0nblk7jTq
yuJrRedeIhTaWBGIsD8n3K1srTJE0ZNe9QwCPPXCEiRxKf5O0opUPPj/wVf62d6w/m4S4iiD1bK6
s0lbQwf/Z7EK3aTQcQpTQ3rjfs7X1g4VV2Gp+/rvZPcNGCZpkodG2AZdmK/aM+yuwpptM/pP5sTa
qn6ahmDPCe7iyAedlHDUmJpr03zjS3gBbvASIc/yFmX12mYD9zKP56hYBENGH6SKPqsapyiorfcK
idjUdpWOgFyVnlsRwHY5Xv1KBGn5Ncb+gFTwXqK2sx8Ojj78XJ8IkOsH68ORSmhxFbM8c15QZ6KW
WzURIdj1pRxVhyHChIduoJtmMZTBdTtAhdHGH14NIqPomZrmNFdvI2RCGM/OsVkLBFQr/uXMBgUJ
3jnm21tBCl2cCwqHdaCG6C04ZnXYfuzVgoacecAPfZDSas5fwdufYtaXKMVgGU5aYdPdoeJSEVzZ
HkH/mnSdwwdMzlf/L3lrgxjFZI7N/vdMImuXOXHv+oehx9xiN3TTkeOH2wzFpDPDtO/sFEPDVAGX
rytFhYPTflWJvv2orkDgCSeN5TR/BRQsW76ZEQ5CZX8Qy42rXuV4idjqQAbkhZQN5n3lTsEIVq/h
MoSJ+5MOsYTKIOmHXCe/MuADAspRvyA8LZOUFfSg9ylLjrHMmGFqmZojUxU36tbpneKZyxlhLI1T
Bq8gU0pJbcYUrhwOc/Qb4R+CgBPr5SYkeGM1JFj+EkjoPLWbeKrYvdOo8beuKss0/94k+GRchdsS
I6qyNB94VWFFMon55sEleYuN8mdFY7juwBw1p0MYYfl35Fdqy+jSB5p7/EVYT78Oeawshe+RW1i9
G50DK+C+BHOq1BUgZOZ4fx58g+TLlVyKJZE5+fv5I2Acm0EoBR/FpHgIpdbshdlCRVUxXm8qvBgJ
bu1caLxIorgPBhUfKnG0MgbFoYsLJgpPUQVFaWGij67wHi0Vz2KY1zXh33uakBKr8E98A1Iz7cQ4
32vrOirdS5BWe7jT8FITY8ef8jddFW8eJQZndXrD4vP4MYvJiIIoA3mze22wK90TFj2HY4cGbvT3
cQqa+gJv94x52FxhPZ2t5T7JunguVZuJEGMtVrSSR7Vbjww/Uv5o39Q7wCf3GrKn43nswBNeS/j0
HNuD0yQ06FYWu2SyLKvuXtRTpA9+4mJjIG7x4RfZZ20a4KCgp0HxqWh6qIXTr6PiExL9LbDQrN6Z
6az5Ann1TtrRFP+FUo+w8kSSUdSj4NmXG/hLpxN55hzP8JiStGU/OLlrgrUmchQKPJie2FLtVDPc
4YxuQQ7UHdsk+WisLfV17X2+Pln+9kXAZvU/iNvkdtfmzAj4pa8LWM9FDVp42Tb3IZYGGaeka770
1Ep7UQOqkljV5eRzyn8kIXWE/apBwypRL6Hzhw8n9KGtBa+cek0XYkpk8ipEVp1L25Reo3rNz5e9
oMwwtZlKjTzDencxcR7cHW7udZzUD1CFTQqYHmEABmX1qxxw/PAwBjPSMQVjghKj+8HNDYHR8+i2
5cfB4tXSTh0aLmy5gbI71NY5ibBF+7N8X05ATkK4AQfSaiBVYQp3/bKZvZwCrra75iQYhUBxT3NI
SxnNroynbqXdSN3suooEgfZGH31jAHoT61haqLaufw43Ck6eFcfg65HhcXla9BFqZxCMT4LXRoWU
6tdoq1uMvl/5XZndSwt5BkdU4p7qaYcz/IPggEPsQ8IgkoTzzauuB9LU+5HAdhi+Lg7vBE4RsJ6C
y9YmJqTibyB00sIOytJgicQ6+ms43Y9I9OE/d0STxc3gOWpX9mjdamzLVwB1IU64W+pqV2/2nEp0
LQ3DqhTLvAaohT/pay4gOkFt0IHM4mamKgVXToLYJfxCdJ4qsm/RrbTgw856fbeY0e0sE1keDY3E
8pekQctIf2V2uAu4j+eNDibL3Ok5sVf981SjbRwPIaTPeUWbtsMmviWBPhKtA/LIbOdoediEQ7xB
OImRbr5ax0AUJzDy2EghQzWu5m1/cmKhpNsyHQkFvBLHr7hE3RERIw+SDd4CRoGBybFmGCG6pwXc
0lZoqVgaHvt9vE5UpYsKgvN5llVESqmkZzuJILTl4P98Nk1v1KEjkXn4+zkSIeMfb2BFVdDncM1l
VkNm10DQOFLUEdmA6SCBBrWzh2tx0KSNgvHMutJf2LDpx7+qzhBLUXML4EpjGy8j+9NT6FrMzinB
LEPjEJaoEbBFvjFCuGJgxIlYvA0ecJ37cCdF1DgoDSxwCHmiS134H/0Ba4js9eYac7eJGjVh6WuF
gAjZLW7rWNGyIiNO/etptvoXkrkyhcFtodemEcBUaw8P+wdULf7/I0H8NXFKwH58l1mskVXnPRyE
hSZhWp29o+9D67KLQRkNyZB9OS1kKfjkp4y6zwny9/YouXAIsPRGwzIbcodPicMvbA5wFRKCXvi0
Yl9czyb92f3WGe51xkBPYmOdH40cbe9o3z9tJtGKD6kYyWULvhiViNrmqM3HTIgm5PxVxg/8kNvf
vZ/gZIskmEYmd8UI+G3CIqeaAaKJmPZW0o5nxs5epSoG00/j0PoeV1u1pF6GUT5GB5wW/7nCZ9Mg
Kxpp/znSvUX476/BWPhOlEFB7T4lXWnztyGKr+2aBKQ94q7AJstRemq4wJgQiuWiEvIam3gXb9rI
tnST3eD4gBFpAkuuzd/Zbi+6DFhVLGcFL5OQlONR0FtHcZPYPv2V6mlY9fs4Rxxl+y/DSJzN3s73
DMxOc5jsr745HjzpRwBUhnB0l2N0H8Ku6kmKGRH5EZk0IDgPO+DrYKhtA9/JaT//rj1waHtIybif
vg1z1nPy36fcD3M8qWHNtIIKswiiRNGdX5HyUJX132ds2W8wEnMHJAjZtQ6WzRErXMx1I2ecWQAv
RZNtLIUxC+GlCYPC9xqVccvhEQCJwNKT7HNja9/DTZL7J7I1CyXWm1tgNGmuVAUNYUWQ1fiX8mzF
pHsGOtrZ071anN7vCfESaiT5GCtkkORIXDq7QHsLaw5SGlZK1yK6stfdrBK/+MfltVyoT0TCio5M
FfrXedd7Uw7HymY18jCTFBGCD6FAmJad27QZGcbUa3Yt1fzWb8duadze+sq54gna8EDzEonUCtPh
GZvxVPidLN9C23JBbuP+dhu3kbwhqzUECV6CTCSLcuhMUf1fvUwk0+2NO8/I4bW3Kmivycho05wY
w4k8GAgGer+FE9o18BqD0e8uzV/3S/MRuTMR/b1T/WVdLIjgSg4gwXqbpTQJBUszh/qraJOGV9+f
ex4qKSBGbjS4FXnzCVno0pjQTaWFZT3F2PEEKke7AOzAOYEflSCf3PujhOpuc5sQXK4JKw50gzsc
O0/zWxzV7CuoK3FKKmV5k652e9ta9ZZd6jlAE7Jq0u5IzNDwjI0hVvmJJXpw0CUaGCwRMf1IyxwV
TWBnVrVEflwKJ133fP/m5m4r5BspS5V06q7bGw8UK66jsnSfAdKtVtv1hcnBUsskoY80vsn2U2EC
ZZlXk31ERAbIkpEgpN3pYb42VRqWGrLMIt+CBqPDP+nW7GQ8wVi1qUbp94vyP33LCDKe7uHL4ecC
/XrgJJOFb8/Hh/LUWhusj0GW4cO6ABaji1vRhOXO7Jzamvs6YfIaLIZNUY1u5YnBI5K3Dw7oeoNB
Gl19ZDWVgHfx8GhbHzcKMSMQ62U9wkxaNMYTB7DSBYOyFQh0ofdJPA/wl5BsW3W9IP0OJn/0iErf
AclbkjjcUZ+CQORP4Ia0W4F6mnk4VaiBrMc52PXfocCVI8M2ZQU5nqCYhUhLN5IPOvcgR7rhn90t
xg/Kj9afN7MjLCPIXY5GsBLIuPUUaaSuSvhdHosuRc+27HWa94UyDBnLbzxkijbt8VxPlsT+C5Ir
7sxHhtY8tWjsar2Fc+6qUM9PtbbKLB4jnd8DFV3rGZFsd4qKVA6LHC4Mq3vyNHvNvKLr0GBfFTtP
1NM8A/FJptXa+YLXsAKSaRpmybZOx3mWxpBnWDU7w/m7nzLTuGD6k/QVqLEWSPqll9dVoUcfv6IW
3VROnk6U4vSbGLEplcQa8j0uWy095kJf3tb0no8c5ceF1DUYH/anVJb47e5g60NACLVUlTMjbXG0
jhRxHCrFNRTw0AWEVVBT5cKYdKTRs7Wzw7NSiQ0yYP+FZhU5UaE3plJziwzJCBOpJbbEFstihUQg
6+EZNzCn0sZ1gKKPLxs9ZVtWGSy9KRL2hPxwjoDw0YxF6jcxLcLDpMSRlmFiZWUBTfoNyG1l2N0k
haqGySzA95MR9q7xiZ8hpTLci6H7ZHBu896vj/O1PdNzeIcSehPNk7UjhyiOgxHEbHTsGWBjDc/R
X3MSahhUsu+GjGjX/E3F5JeV33x0SrqnohaLAxNwsSxnywM8OOr27r1U+ffVcT65T9hd15SwW2Fq
L5UtwwlvvWPIptCyNjgnplDIyxk9qZvcp971dLSitVlc4qrGDeKiJP7o6LxZo+GWDg870kLe5mCw
ps6gMoi46Hd0rhyHsXrrGM5W8MPLLZ/1vUbkF/zE5RRfqZYHb61n2svmMks7vd90vZlRe+H2deEw
/s7YIEWLpttE1EB2SsjWpFSt+6xJpcCVWlMKogYP/OrjNPcxKWimlJNezO/SyzNyic5YMbprqZGb
VFLpTouyB6EnFcHtAVEpnKNFiUEnEFeDDopGRK7atrGT/w4slGbW9w1W2vSgQhT8YbpmT65XXI6Q
w5hLkN59nrIP//R/+vsIROJh3HeWFq0DT5qABk+jaEx/+3ifVRdbuSJnmuf1/1d64OfcKEw9jOmM
gl9RnY9rbVdfaPFWKea+Uf8tDoOOkD4WWamCDjr+5Q/JZFOBX2yEY32PZspn91Uzoe1JHg5xnVBE
/7uqTDUYt8jTrRo+VJzfels0Vz11SAyaaJp2qbxr0j8RXu5jFhJyRoJ0/XKHQmCjmw5NTP6KiBLM
SlVCIqgEm1D+QkQjXqvegUp1+147MTYd8pQG/8H1dOa7CWa6y1azKybrjcsgWBZNsQ0YdXC/Ya8G
zF3OQvkhbW2/iHswBYYZ4SVqw1YzU0zSM5Vf6YdKzJ3MfwOniwiq9eAOmodOIDZ8paCOy145Hlpc
u4qqdO1LVuzN8Jh+5dNTzuF4/esJcbesvs5tQSebLO7tchldgdVILW8+TBctsiLlh6N4fC4Q1yey
WI5L756WvNtWhVM5i/a67R9I/pO1AedC+HtMSs7WdKNxvhsxxPbozTW4UI8IkF82fHU35VcoCG9x
/yJdDQzUsK58X6iUQm2YyNuCOWjqbn0KQ9Z6JZi0OcSqe7wZa1FVw+TpGvGnQ/FJJaW8tMZjrFju
8sdGJxvgxiPxJJjDrwQBF3/YdGE7uqwtKJaTSrvOSGcu2m16MQihQNsgGKwsvP9J5xuHGL/MNNVL
mj4eTEtZfMdaD3QsZ778+CtlWjIWjp6IlbaFsU98JkxgdOAhZ2khkJO8mMFtL6uE+xm2tbSwJywx
VU5f4g5E8I0hGprHWBYJK38lHiGlBOhgc7Vb1hqpkgHOqM3GmhN2v17JvFEtHsF0c/nydMmvfabk
QYr2B1IJwWIPXMi+FiTFrsRBKD8kU2BHrDpExXRc56e6NqFOjqps9wACqU4GjFwQRjMgpneE1viy
l2Io1ooY9YIRP1IPlwODJe0f+vOzVjAaPHbuv6wz4z96XCkjUdmpOho0SXYi2y7rfApyF21rdtIR
30DdwtMqB9EggmQJAssMk6BW6chmlhC0lTuNn+ZUYtl95tvAbsIsYUoR1DShBmXYNWRBmw7grMoT
80izidUooKUtw58Z4gdqXxXbG0uY50eaCOja7tBvglb9yKkWDjeGN89HJa7mCxy+qxANmIl2olND
+2Fk04BNi/0LWUdpQNM7nM8fq8J9UGthcXsa9rTXz2L0nlfRURkEuhzBGl3TJ4kbwVNqMKQzVYzk
cc2EdJV5VR2AmvnP1lUp0IY4UV0xDzCNv2iRxg5/Gr36kDh4NNVmkas4NmWIz7msuDOWhXDCdkN8
5ZlRyLLkydhY6FNOBw/DV7dlHLqhKBJc9Q16BjBWSE+w84PL4ZjfxQnMV68g1BIN5J36w/MZXKsx
5iyscGozpTwQwxFdeD6lFxTDFTYa/vZIKSQhEkJ73YW3wmmPYX0+QVNUzM+h7EGoxO0pH2fjZxdV
NAlwzkfwK0gG0+AZ+LqrftHaNtwzKUbJR1b6m9pFqUiPp+6h0Zl9RgdU6/lKNi+xtBa6QqUfXyH5
cWMdrE+40F+72wQif3FO01rKXCp3WXuWaKHTRJZCgslB01AGF41CaGKKWjYnlo+kaL5YgSz+DvAe
u096+uRPMAFMbwop2kXh3NpWsAgZiTQGTyCEEykNjawLzeVd/55/St5PJCrFzKORS+TP0XegC3S/
QU0C5hLMdLX9+V56BUidscgNQHKjSQFwL1daqYNaeREwCEGVPPskNh6823Dn0d/8iCe2f4805yrv
0p6tEh34OKnGwJJSGt1s3hPYRJ5G0vy3lT6O/tggcf92IuRxt4mUE/18TEczWGcR7cIjbIFJB1+Z
bsZsnZRiQ5Fm092cFLv6jjRMgXQ/pF1vsBp9DzarolzztLrbbRki126PujFjiJyRfvZfim+s3tL9
LRjKBhORnYwAheBQz9Aw9Mr6zONSbgh/sv+Tmr8XpZNSZkE8xZLq/ObrJVa7df9BKMJQwzA9NQ5C
ooRtZyS9SdxHiXipnM55Lo0E1EsOr/QzqpEl3Us+PmLB0wJ5njNuie8B0ivSJUwry2uLhF3PDbXN
2fBBDWUV9nJ+CjdhpieNGelLdwawiHtRfzDsWiwc0ijYo8DCDOR64ML75eFT1TQYf7uLj0+GNkuG
L3+MCI9v/rmRw9NypI77dDvGrXpzJcjkVxLw2PFelBSePfBoYa5RJO5I+uS+x+bKgZ1cUqrSr0s1
m6zWpQgpYqYPfQKrvJHhw9o3vOtqBkzmM4MmYVWls9OoFdrgJZ8lMnRZsyO/BYAb/ZCDIo9y1Io3
o20DghS+zNauA7T0GIFUHGLxfh6SpnxDsi/eQ9s74Dvzy6gKA1WlrHqLmbBp/g3p6zJnLd6y9GoF
g/UYwzqzzNhP+wpNkh8R0NbFYf2FezhPlcvkwKw3g76YEJyBPB9G/MyzSueN0DU/J9ayyZ1pY9dP
eACoHYplqQGJKUa33lloMljOeZV6bvpenCV98D8Xm2tMiM8x0i6IyQWs3YeIvzb7gn3KPWVHQnaI
aE0/+/WLm5kbIxprKCZrXt+dM4R8tpPs3nYzroMi7dELyy9TqBdRmHylL5RJ7YVFY8dTNfCwEVQF
RQRqIXOS2RoB0qzSS8IjoCpmgnLSVLEywJSSOsuSaRjYKiXlCS2Iw41BuGypIxsCp2Nwd+wuoRDb
OZDvSfv+y7aclS5S05Dig5udrAubtVIjs3o/EtIc+GUhVoipUlKhfPOpX1jbZ9HBwJAMzLh7WhLu
LlgdXgzjtwI1/tLjBEKP+w5PbpbaB8whJeL2NR/tuq81Qnl1/ca0s/PcyB4/ZqGrgmOPK0J+WCzv
WTk6M+jE3Thb7yCDUrLZ5gyVewrnYVtSnOKQXI/ieOIJfnJf2vYrNki471NRcvLenXKkseF8xFpN
IHUeMgpSnHOOR2CXHMyyIyoD4sr0z/YaxlEW8aIKJiYQufd8MtRZNzcJN9tMvWpAeWZIDI4LVCJc
EqhpUcURPzCglpGDhZYnaNxnCqR/2E9R9vCBichmy2JIHYx06D4JU17aKFXUc+y7yzozaFWK6VVd
avU/J4WBPGNnxQlNpVoWq9Fv/OOMDdT+f5evnoaKEp3RE2OpwmHrWJ5Zp/bO99i6jow2qzEOgZVw
NzOWMpx17a9vL1kMOidr7Q7IJ7f/qtRybKxzE47Kx1zXiID0dCnL8F9W5XQ9dw1/mnTWPpfx0lvp
NxTJ96URDMtwidg+ZJGhnFLviAlMQIQB8D8V4IqUaycsM/s4ubY4h17X4k/piNkzSw+Io6gHwF29
ZmtwAF9Nl/9N/djgF+yUEckThWkE75UZf64ok6aYkZs25VhASKslnI6K12t4pzeAAQFhXidof7ak
YRKqIzetkVD770JixkHVbym+7CO10IG2MMJCNB34wXHB6UceYhB4DHhEGpnh+X3tWacNbgeLmKKN
XCB3MZt8qL3a5Xw3etKD6h66o5PHdMFy7VE+kSadgAqoP8E/odOAygP0iq7ZUEra6JRzi1r1H1pB
hHhSuIdZOC8NY+vODDbUl/uxafhABaYflqIox8cqJtsjg/+tvbktp7KAiqr2TyM9xJKme/xpDpIr
hOhVtm6KSaFKhpM1Ltci20bWd5g9FsrzFIoRYRbVdOYQ44TEWTgbEv1hCEqkTCFdFibZzlB+CzNj
/s4G9iwnvfkq2ZvhKaz6HzTYy8cD2Y3/qzBnq5Ehu/os/Gsrg7WcN9g85/XfrARpggscynWsAszn
3dkt64Rf+e8EJ4+06mnSo8xzcjgdOiS0a9ApDRh94112KHz9OuHryfuntAfMvkGbMvt+5iMxXBzx
bVY46EVdatae0GTw4ZFW1Mrcw+QxpRo3wVzun55bDpVES4ol+qUb1XleYyj0Tn240VcFp4sc1lBN
/i5CdZ14JjzN3BcpXFJkFdnzp4gqRKpeCJN0CcDgyxWlX7vFmzKye2RfBDS3/e4UNUnxmzMo+oYo
3TWAQ6+0XXKXsStlXTycf7d5Z6o/N6J+OKMw4rptlpVMbyvqAUN/WQZriQp41eKlz3+AzOkVvE2Q
g0181q2MvROkkAAWo/nQK7pGivFrQCjFVwjtZ7vPP56b+BBonrSdDMY6GmZFeSo3k8BASRavEyDv
cM8jEWTwE7ZSRXfTCD0pme+4RD7AAgLBsRLMPzMwjxzQRYYDr9mWoPiMre1msxAIOUlJR8+8mC1a
IESAhma6b/01SFVyOEsvZgvfIsjs6QY4k9+fdkO6HueW21SLQBsCYhF/t2IcZkE4DwZgVrSLf0zn
OCKeD3AhyyY+9v09MH2vMfikhNnSJI/N/69FEVnrbFy6+QAMuMatnqgEjvuQOwqwhbKC7Oti9Oqa
LMuMzNj4LVwr+bPwiGdQcUr/AvzDDOoQeUZ7zaY6e8zOtTTEB3ysAXKdC6Ts8bICrJsNV2VujyQs
qoLFvFtjQEL4ruED77LhjjVx/cRiNyvWAFd5Mo1keVmJdoHTsHH6ai1IcbVQm5OdGJgJIXeDfeaM
1YQlVKndXJuJIzT4+fF30JfkSD9kTIYEd4tUKXPaov3QFiW4z6FXUSU5IVrLZQpKUH2vsvG9+Eai
I23dLJl6PgpYT1dc+BU/YOCqA4LS9TKtSX8BAb9lyT+KKIDApUYcBsoaUn/wfWHp3P14r+URCQgQ
3+upfa/tGiog8JH56wOYMUjZBMB5wpNVz4ZknxNJfh33DOJzl0zhkGhW7eYL9/MKJUWjpmKKoC7m
csVsV9eXaV6Zv3BR67UbBHTQS/zuvjZUfJcBwYHXzcLuGoKT4jLzZ9NTo8JxV0bSFbI27mhIM26u
QKZ+SyzehunjcJyJLwdIunAuFBM8ry7Y5xm3uJMwEpETHcauLvo2ItGscWnKugf2wLc6caTFpZE7
bQHCwqpGrKEXnsn5wguKct3D6MHtUqyopbE4MutO7eCzWUydTPQWb36h9MCiNib+MtWTAzN9Z4SG
vtOR5SRlrNTPXvKHoV96Gxp5l8Fum0JB0fWg2nO+yK34+ehNqs49AaMYIIPSNpAUeJiZzmE8cAlh
m/Ge9qPc8tGLFfrswiGnLWQwRmfppmBQjJTXk6sBaf1DFyFXvqpL8x14bbnJUolUV1LjC8SLSWJf
Ig+Xd7hr+TEC6oXgI/Vmk2YRZZydZQStBAhlC/Mj2wVZ65WejBk9/aB/mUxXdejQw74VvHpJY5Se
qVvnDghv49tb+tWZMcRzlHXoN+ChEQxDaMLWhqVNJFw7tz8bVgwGZbL97RLmxeNzbPB9fQH4uOIE
lv4rVvR1qD+oLxQJNItgwASikYcD+zZ+JoObzjSMlul1fCUVUPwYpz/mPOCe5WjQmjISf1ty4hKR
XjW6p/dgjlLnHjfvvYbtq7oKEBR8WAt7O5MNZFbA6saG0zvOCGVBbG2kdfEzqhr9C+aR2LTi30gp
s2mLTpBkJHTZFAUv0nXPbvMkGRSuXrJLopgz0jSJONwLZ0SSu+6ZYumvp98UhPZHlZ8HP+xrSsx4
iHtOAOtzyQfsYCoWZWfY8bk0ZZfvqQ1knRr5Z0DGlOIHfUJwqP1V1YsEvLsF34Djw+RdUD04nZam
ZjF+bAzHHpHZ3qwIi8xYEDCUd51NI500R6mXUkCaC/rJAVdgTThV2Kn9QLjPrjJ+kzcdgg/dKo1/
sg9EYGa6nUeX+y6OpvkfsMk7+CAeP02L4krUyqnCnljTsmilEwMp03oWVrFQCfmGfZ2onwQHDvuU
68VY/bm2fl4umCxfAJIKWXdKMpBKSb9m8zr8QnjdJ5eY6Zm0cUfX7Y746i38RkNK19XExY5ZJFcv
PHD2HgfXnSHqm8AOfWp2qyQ2W5BX2ThedeDCU2EoPwVED8MHT0tr7b+1Wn266tb8p+HrcG3VL9uc
Hsor/SuXGqtJ6DVvcbe85TpAjexCYtU23B3uI2ARXyvi1AawK0VmlRp09rRmW4Gg9ER4Citksqds
o4dH/Geyq4aN5zmmLGyRflcBlcqVfP0hw5QQ6+5yJY3lnpsJD2a5N9EvP+cd10RL4jLqJcnfxKAA
lXdNo1Xnwx7yjaoDyuOgSGoeYcysTCNvoVoeaRQgWZpFh6XjIsq51oEQ2QgqyIv+bhl0KvzV+gyN
hdxcNhMTniGO5nJd394Lcz0nGE2HbEK2L5Nm4v+pEZTV4PZJtyu7Ia8p9dXnZxdlas/RJ0g4Ub4W
zljzLpXshBHunfhETwErk1rniPIedOF3mmxgsEiuW3BRGpD+1PUj0bObuS0bO+h61Jqd0RbUEYqT
CxpPKMeGYdPU4k6Cxto1pa9IpgeJqUw4WTx99JEE7+QpGZRcaVDqq9LXoBy5wyNP+LiNIc380xhK
EfqWhy8TS+XOYrZw7mR3WN/XnXh/bXIG/1YcaaoL9ae/OSYczlaaZXiAVz9NOA1X55Hdcfj7/1M3
Ynz7eMZhOcMcTKwB9QYC1xrKyH9VqL5RTo2d2GnAPYgXotdlQAGplNcOo2M2jabi7aUEjsAGpUZp
x+5VaJ3/ha0s/o+74zFrlWHtAHEGLoryrsnxxK6UuGi/NJZ/5CgpDtQG7VpsP8Mt991FUtVf5F+c
dR/Srtx6oBx2w9pCXbrZnEp3ua1Bcvt8CeQxcA67sbcSAvH03ksu16iqI5NJ3gSQcRvOFa/B7QQn
zWXsB8f6yP0EtqVJZXdDi0ZcRam0fnHfIYazDQoGcXycoDTHyYF/PpUj+80yWUpsFb8msSqEkCsr
6S8dbRdkEIlaJVtFM6oroYwO0AwtVgnsBbzfVmdyXbDz4lXqkJmO30UG528JY8m25rKq4JrPrHcK
IeiHfSY77tE+B/dpDiBraLH+JWGJtCrYgLnBkyt4zADFYvMsvf5nYXl6ftaMhmY7BEPGvrYv23uA
8cQy7F1ZrwiXFuPVpLSP8bWJegSPBmMZ56sD9MMmWVd3M7pvHV6CuiG4If79IZb9jKojC5dFc+lK
7zHam8/VsEK0JF2knEpgS4wpZn1UiySSPosrQFPzPV5esLU/+vmnAOK34+SA+/na2XYce8Tk7gKz
r4fHakvt05zY65CtWOlFhXsobB70WyJOopBDI/2gUkDjGYqm0d1LSK+1ax1vmWJg/xbexkht7n98
JIFM53kG31htNRN+8ep46sKUTlGyI+gHEWe1tJs2rg/QrgRfbHF+V9DaZusWcyIi9lzDsTJw5nxM
ub8G52l4+Tkwlykh11SxaoUbLSsOENeiIc+E19xc0G1XraWAKX/lo4vy2n5U9D7IizJ/jgENTpna
U6IyDKuyk74zHWkhQoGf+zs2Is47qiu5LOnW8Gl61qREBkRnmdsn6jMRaPbDu4Sfc5WdV2qT8uVE
6Y6usZdOvNmlPd1MvMiJ1W8R0TGchGLAvoyue66TOF2wqtKLZKGiGZ33yUMfvCdaAROveddPy5eT
2vjpy89m5zEDBQX/IlDPXXjfPXCHw2h/vZ++3e5JLe35zJKykEoXmAI+cAEPeKvOcMQxlyUg5DM1
n3fKcJN9lwMPWWk3rbJoZTEw8WqVGX4ZdXB1y/FkSuG60phIUQl38LfFZXq9hOC7pOdLYklP+oZG
MLj5W1Wr3brnWpGOqh/6ySpQizD0sYNw6UNqCs9EqnIgfw4/tyP1ZdUbbPhZ21NrwiH7Qc1Z136r
0RuE+J4YFL1cp/OHWpXBuyndRQRDY4cNQhLhzaOEZCGYBAIuxYWY66WswC3sKqjROOTG2qHEJrMm
Kg+eYzQoZAzcMi8Bc+5DdBYm8hWwGtflN9Orr1WX9/mA9BGKWMIKW1RRaRTu8m1lJd4NtWIpO8hy
lOm38YT3kdCk5DL6Msd3sF3sQoyK/ndeoM3OX8miNZrFByAikOFAetUKJZGkPEULl3iui0iiuS+k
guE6sgQdv9fIb+RhVBRHSE2BFOmQPdhLVyvhpawAuEHV5Ej6ZYOxIAH1BR8G2ssp+Ou7fmLnpe5c
8XqriNfd4tSBcmR4KGmY4oVNObmex9NVlocjvsn0SbGdDRubSalsdufugonMydBkEwlGaiECSyVI
9J0U5n8d0jxDMgr/BJMANwNZ1v6AIkXsq1QjGnHsu88WlRkHlM3D8hKHPT8GZxzcOnpDdYqSVn6b
urM4Ke1eAgufthdFzTnYRGidBlr2P3ycG8lX4k596hvaw3Q/xejg2aDUQaUciFYwOB8HbHn2z94N
RLGtTwVeJEDPclDsyXv8aa24OUkhCJApRz019U+83cbcPnTSEmjajI3KZOc/Bvfjvtj7ZP+d4uzk
ecp4fHx7C9xAjx3+1jtB/aT3tecgv39ClF/6+k3ZJUgctdMX8RjrYLxk7xm/KfIeMRgaCDfPGdpT
jG0NeHNCB0LvnkMoQeIkpfGFXAxAEamAdxJPpDQSDREpM1Yb4hzBoWetaZJ3aTAiFn7XFBSK9cRy
8Iurp7m8CG2+tOUSxh3dLdSOmlOwLzJzIPcLQ/0wNQufePmSke1zWnh0rH7arYsuEqPAlrGqJZDR
7QVz4FXDEZyyJ6epWJVFM6TIkQyExHIXY/WhG91N+g1mG9z69aX8u1nmEU3C6GlSrgh+P0xXYROA
tTSXqlRUiYQHABD3UIKiYUDlH+nzOMpEDSm9zOeLmx7VcZAzZPZT8EU8vxaziMJ5gF8B2Ktb8hwl
6q0KV2kugxmZgl1LtpqfwAE/yu1kYNXKWgoXFC5tsmvsBzJdZ0qUNKxK4mjcPVN2Obl70zMtTnYe
q7qiullOnpP3SQC0PxsueR5zC4s5Ce3dmjlJo/EUlP2Cdy5C/E3BEMFGJMaPHrdOIEbyok3jYqcH
Zz6QeZT8AZeNeGjZCvEllzEzm7pl/Mfy+AcTZKs0wQAHE8F+5PO5qUTZvcSiw5Mfo17oOIkRXJtk
G2xs2oipaSu46MaKezZn6YqhnDVT96ucnRRZcgiPLF5oxTChLuRirg7cv8fZYILjm+PJ3QUeqXI1
ikd8WfW7O3xNBz1r+/M3nVAeqfuxHkYoIoNBwxoA/HAkSBLslpwf8MnmhfLtkapKuSMWCCBe1aRd
+3dqzLxoJxUOVrcXQ36LwJ/lz+afw8McD5by60bzPdtK+LWnEmcfXsrsfA43q7jsVTlVLdf9wU2s
mbmGtoZyBtKIw4NNNXrmwPMeoG+Ge9omaba02UGc6myy2R3tHoxg6J7g0om6ETDt6ZJ/e9qrefMe
PIjQA2c+4pJPoXFPTYdlV4WrAn0JXF7SlDFDYaCopcA4SLV8CFeiu8xpI7VEJVK3tcFLBru6B5yn
q7l4/UrqCbP5VDObXDoTYdCXidbkCpYmlS0kqdAjkNXhfx563FAH+/8pS5fQ+MJOARS5HQdvGop0
0BmrxSTh/NnSu/OjEnZ2oc24VsrIR4qs1RhibvGp5imXzb+qD6YWwzhQzWEMu7OgDN+BCjaKKtnx
HOm5aMxWauQuDHihV7n9avX9JDF5iiMkgJWtLcvoWfxfdZmS+mKmWOcoghAFHocDP3pU3OGIIDoa
iGtZ0qlUOXl29iUtE6zLKfKLDRRSA1JjuDaMJYygtLmDADcCj1dZXpyAHOSPr0sPSqnqoPgbRrVd
aCFOcGo2Qg6TZ5SQRexQMPsU69NArN4XhaAb+gCJINp7gjA3Bke72MoVh/BO8TRzAcmm8Y4JRadb
uXDtzg0I9pZeAYfUTih3zkU0YR0r2CpaHGkEZUdQppOyUpJCKDXs1+2Id/FOwtjURwNTZC7nbeKr
MPp2LI9N0yF5Z/jCS56sPqzwRHd/4GmDnysIE/0NDtjj3a4wLyfgmSRgG+qVjuEYlb5GF0B0A8sL
Q7WVb5dd1L/J24n5Fe5XBWUsjlNiKA9aFmdBv3mn9sftRNes4uXWfm1dzOSaNZz0LDe4BzBCjWV0
j0wfsmSsps4Bid/McnSmqv2FRoPuDg1dvODu9eKzZMcim4/jtu08NDTiQ1zCUvuhqfciTRJMxzX2
WanVZX2dPdc30ZQja1wDK3zT9giS5zVNYfaJhFvlKnnmapNgKCk/g9scOUZ078mmRCpkw54+nQMY
G4tIhhQV142XkcJnin8E11Zi4qnu3dXdensKDhejxbL2NOzjjaITqNtTQFlWoHN/QwYUXNQg72zF
2JLr5iqk0Vda9m9IueHWvjawwW/cSuGtls0XfiQOAs6QYHTDQExNLCSnDyERiz5BRyPZ3cRySTgK
ecW7VjxbjCbs5Y9RIBkGT/P5LnIaW6tqto/jqz16sGvGbXU3CMggBswHWsh6u01Sx0RZKi0x1dx9
Xm13vWY1ESbTIIYNTPh0nXMi7pOTJ3xddq0DKi72zPu7Gp6QZ/dv+cbMYaQiXyk5eDRjjmaXBOxY
IWIUG6iDamP6BRhnDhseDvyfGJKrk5rpCjA6tGyEYZ4OsPb9dTNl4NKfay+UtmMQx8ViCzIZXkTC
7B67YzKNMGBp+iss71W2Eh28zOl9ohTtNi/PNZO5+If0NRsVYCV1/vy3RGmRg/ZkQwOkjXDaLX9I
ynrrowaxL0sYuBC0GQOrizwvRgIKW72yh+BbIR5zJCcFfbbD9mevLym07QRy46mwE+J7lY/PNv/1
CZr27hiAoLDGb6lKbqmWSaDpHOId+mDxO9j+7WB3eS1NactDaHtTS0iSJ1n7KcQW2ob22e+1Tc1I
NnPX/vvXMsfjO5rpiIANNPH+m9ww3MKeD0IvQzNNh3nX4Vwv5eGClef/XEKjwE1kfNTmHsViooRq
2M8f7yUyv9eFeJjvLDK/6C6TJyJNqBV9ppJzzZ8Yde1tOroLSKeVLjFF29hhMUzgsugPZ1J8ttKk
VqLwGnnwKlkjXKOt2TBsIfkkcrofHhB3K4e0vaMI+DMt3M/bGJS2b+Xd95L6i6ttoH3oXLIRES4o
zrKVS9KGwgzl38HKkRs+1f5/O35dlHnNlnTh5p/dOrlyO36UX6aBY4oDAlbkYIU5imRcLe1uGijr
XpBb9k+kW0SZ1ZFEaiZb/0ba9dVFUTEwo9gvO7V4ETqAAK7QJNzgfcb2imZB6/naDAkcGfuapyRZ
ymMFM3U+ijiZxdVF7lGIXtawEGzTgz3t6KYrAu2CPAtT6mAs1RXX8vTmHfLQwq2y6G5zY6dDa+1Q
l+jaAhqfMiAQ/+g3yepolzYV9na4cdrDxKj8yYXND7R6jG6Xg+gRGvKtq/fOepvQKGeCZvXf8ba4
sigOGX1ug/og8BjoWP9htsL6S17qXsDf99cgTQ69LAlGFhnpyxPnH7Z5P6YL2IHRQDJMN0Xvegqm
hjTiKXxiu0qlt6a2P1TR170GCfvtSX9qr0EIYk7YxzZyfRWApXpsENZULFI86it8moihGSyz7N08
MVNV/qWt6/l8mMnzN0jl2gzMAfYWcjMzJmOQo3DTkWRxEruOhIrWdNPSEwr1QipgG1m3Vt0QcYIp
YOo0UtGfHHrebG4EW7zDYs3sVRAadq9deu07M+9zX2pKrJGr52SP9K9mfRG2qsRNjaJdggvNkg+0
XLxbUkHwSmepnj/c5IhoGHBYVTn7dDhnP9MF125pRV1JcPYrytI6FPNLzVIydzvEhv5td4O9nV6c
1fuVYFBAw9u5nolrn/YvrcAn7GPon79xtp9zs9H9BkS/co3Cq+BeQ4wnF3Eq7d2X4S8xaCTzMgpA
qTaeNOOlbmNfYj3bUgEtYjIO9LOrq5RSrh6k1wljbIWUKEuKiX1wV5DNdAk6deCkuSbxMmfMhZG+
9Oc0oXVtrqAbH+so9hmb3NM2RmrqAmf7ha80xOSbM7jO8QN7OqOn+82roCDfHXqL2XlG8LUiSUsl
taTbqgcihZjYBnplpeUMD+MhgJiB444rbrWYvqHJIygyqlvim0G6oKOgkyIYT2ouAFWfo6zVw3Wh
R0SDVas2ACyoNbudXnIdMOCHF4IJRN4vbPxWI6PVIRGcM80NhbH5iGdYWJOiydmryXBys4RRYaI1
zCQO0FdN5o8thI2wUTQAyUgARx1xCxhTjWhzWGOimeaLAqsynsuQxX6rK/Sdshteuou9mw5z0026
FlWTKXR0J7Vwia1CuItpxdZf7cwYObiJRuCtm6/Vad33tvX19e2W0wRrymdFxUaLROn945m/wMML
zIejxUDxDdT9bL766uFLk8//JYM78te+EQg0tGMEVniJvhJzEI8icI9aFHdPhsE4nEy24nQb0hr6
GkPaf4T+pO5dtpMutIgYYVq5IJw8A6zQeTyLetSQM1D2ahP1VaMB7qVq1dgbAtsueCM29vba/1VZ
3tcFmT6qMIw2r8WhvY6g6TzOIcrCM6aNQUeNnhdG7fyfdPHC+Lc5E+ugk7twQpRyd1Fc97H7QxQI
4kVKnlhnpPXkYCiskXpME5Bv9pAMgBG6TxGBySYeYjqzk/HG/nfHHHoxFHsvDy70Ov+LFmDljEYD
lq7ijLUzWWjR4+aQwI3kH2sCHCMmB4n2GkHetSwsJvQwichZ+wUdQesWMWH5rcCwFU+MVyY8ouRR
bcyrA/1UqUy+TvV/z5bi7F81+K1fZm6QlS48ZgdYvv1DI5QPkxwyMPo5QRTBXqOri+ZgX8BeHpsT
PCRrBO/yy+UrULsDuD7xoO9lYjjfsojPyNRxXMbW2q+GufC9e6TC+0A1P4mfk67vnwE0qLPjtJe9
g+v6Q8HoedWC2/3o790TNG6Noq8Jq51vaLNGt5nl2KTKQ36+zMYehUN0v7wZs9nKeZ4WAnPi0hXs
nfW72mgCT2o4mE5+eAnnWHp0IzfJpmaYs3p0tJ2/fwGw335s+Ihhjbyq6iXY/QStXGm89AyJjsS8
MS6TBrt6Ow3O4VI3Y66eiCpemGq8zPP4Frk7hDumWdA6+IiYvMer42VpW6xFELpiG00Cqnd3xPwD
CztCjkei7OQXttWjzOp7Pc3Hub0aPxCmPyuDz5KuBXmavWqOgx3CaKXt7kkwhNI4vMxFQGLDkuTF
1qiQd+eAxrjUB4dQGIM3L6jYbs+Z+w2PvBu8J316lZRKhmcpCWH6UvCU0PDAy8arwKhhsPcLI3xW
9/QMY6uD4dwxOFDZ2L53Gb6drmIYOMP3OI2ZwW4aWxmFXZxeDGaLc9rfIkegMdSyMh1bKR3RDBfg
t1EBdYNXMrOn8Do7kbIEpZkIBxpO7x2+GEAVW4E8j629K0YHnLSZ69diJRHhj5bB13y7Jn/pZYAv
jT+/fbaZpt079m2A03yTNSgDYJmXe+V8MsrljtX0D3lTzaMo9nfGO0hqShc3JemyX9bbo/kcESZo
ygjeNEsf7XnysVrMqYj7X7OfD+dKr/1SkaDPezlM3wCfhhaJ2aY+hEL4mi9Lb8zBRrPqgzXtbYx6
nQVslGqxNyYT1mV55vB3O3wVjIQgxH3wIaO+qalTlbUB4HLGKv6ZdKiHdnZizDbksZkflIZX8iQj
hA5xat2+YBnrfBLzwtYQ8/1k18ro/GKELad3K3ylJC13qkTGk4gadNXw3sjske+hKVP3fZ854Fmr
w0SRGuVw6D3J9EfhSXPhfofVYiHNvO06KaALTR8nlsx+tcTL8BleFWBZOj60rMo/2CyRoWkFH39U
NBK/X+NhYM/ak0xvBgqrd0YLUaafzb0EGrhqHM1mQETe8F9xAE9vprSEe3ky+/C4tKsevB1W63Vk
tRxoZETIJVBUEbGCW/VC6UuaLC9T8I9fhU3ggPn8ugYTTyKAblkWSBeuY3pVgg+v9X7LK1gi20BT
PyW8n7W4YPZwt9nP9RNS6uTvQnBzNbb7PlUE0Fd+T4FmhDFTNZprsiWCIYUGTzuIuukg4r4mit0m
aTt7jNPMSN3xm2n8vzdktOJZsL/r5jIcy47Takbpa2Q3BdkFJc2YoN+eBciMt41bvDtQk36QOTK8
UlfXfRqvvE41WuT5nnsc1UI8G2l/GalaqJV7bt+mkytMc7Lpg33m+U9YpcytI56xz2SVqihXAO4t
yJmp+yLVFSeLwVoTPYE90fGw0cSO6MlidTYzJjs+qtdFlE5jQJ51GRvqNlo34FPXzIkfAVD0/T+u
Ki+ZzlJ4aS6DgQS28oHeu1F0+DjZ1sqLtxPp6S43oCdyvsssMh4XFmlgEaJVxonAJuWZSLhTgwNe
nV15BGeHVYu80w3G1F9WdyBlRpHix5UOIUlDhEy9iYrg2SFIuh8RpCNDtivqHatsXNmSb+b6XUXR
33kxmrMPxaCc6kcHbEsJg3hlGCRvqctFRppNbgEHYE+7IfbCWzenPyajFJE+GMwEQ+s8vnYNCfjd
dLSDUjoQ7eW6szGZGBUu42XF0uSaNjELTtbH68XLBUGogAx/HOxljW+Mrp+2g2Ti2WMwusEDDyKn
GIZkLaoaeVQ4VLQdaR1Cbe2N8KfHfqvxUmeo4jt4tupYYYnt6qZrkYoswTEEhuPBoC+f/zFQ3XsO
QWiEPKPZ8cjI/FoMlbaMBhf5RMpg26yrKzuaql7waR83ex0h2WSx3O+gmnqfatHVxq61nUUiiCLF
uT7P6ekQjq8y9ELKUDiFR0gk0sDApNyOwLZE3AcXoC5JWey1WCXmskj6Ea6OzPtbHbz434U2iTGa
ziC2tegJDx91nVv5A9OFbIaKOX7VXFnPvp/jvDdCl/VaD88ODlP/a+ey0cjrCCcMfKWyI3EFm5Cb
pwZJF0n6ITHUSY41khQYmdetXB1hh3fLbDdoIJc8nQ1CCrL0ucuFrsrqbFMjpE43ey0nhKFqpytD
RbOi0FDq69yuzDhn9b8j9N3r3g+OmRVdcv7DXPZMFWB0Gss2Xw1oJGE9DJTqBzCfwCd4W4fW2/zF
uoHWKqYrTIfnbQda+xvWsxtcsLMoeAuu5uORpTP74zgc3NgiiEoNlh39oabWeua9pRa5uhlnjBt0
OtJ/Ue+Td9tbAp3fJlc8/WKONnSmHlzCdFhPRr2ADK5AkaBfbvw3U1LY8y0xbiJ2srqxl9N+5USO
WD7krE6lnVgllH6rPPiP3H+bt+EupDUwWSKQ5RSGOqR7QTCo49oTttkna6aDbpG3Xx2wSn6EgZZM
BIOaLCFUycrp9GoYQJCzaOd5grrI0H3Ddos/poxoMtC5EOLV9837Wzh3IPrBNerFAVehlmywesNN
i8isrhbeqQGC8pY8g5wbbpp8Z4dVxeM+6kPf9qpgugMu/TPqD7vebPo+7Mwlr+xBMAK+AYcbwyBr
ScLswAdc99yNpYbTUUxyhsr+mGUmLuABanNazVc2UaETG6jgOGOjJp6tzVzcyrTjNdw5Wm4LsJCk
YqBisQKvd/ARxjfpWCFVNqKgkFYtdNZubqmYemiW9uzACwT7LhLsaCMtghfEE8pL0A9JQiQgk/PU
Q8DFLNX4DGa1aP7Tmb2HPlS021svmZ8FPMwL7KCwoGnYKxgjDe/gqNZwDQqqKSltEtS/IVLcOzl3
0o11QG2PVK2tZQaFibHSN7P3bxpzI97PEdDEn0EQ9A0S8ToUMCmcc56BGM0yanUWuZS3v0JkB6mR
T3M8cEU++cJwHwjySBRlWEvRC/3/w39x0md+s7vcos5oR+2BYySRi6OCsaY98vzxqz4ym62d7SQg
vJ7b6l4i22ny8bRU3aJOh6VwhWjQ5rqXXvBZtyq7+K2L9AF0ZR+zHSMgU3zM7MK64E3IHNvynbKR
wsr+e2VJchWFXAWL3wUQD7Uc1RU7wxCbV/Vfd3qTLcziJvKHiGQH/f1iOv8ux61RSb+Y52aZUeop
EXBddqakf5waGRukidSBjjThHruTT71A5v7hmqh3hMSHk85ec18CbZSFr2w1M+LhyZafdZnFmgul
D3NZe4fXeizICNIzgSvht9F5ySfJqwwwrXXthzugUrnQDx1k+w7AVFA8duyDwrOvXv/4NKTa8A2W
vaGctAtwxwHASQz6cXNICg0gW2jATJ85Xnm9iXXMRONPaJkLYXmcv18pdPoRbovw9olrJme8WydI
zgrcH58M/SLh0RKv+AATRGATgmZ6gCFhCDbxkDOBTmBuz9zkOSBvp9CkpD4vH5/jmdj3qihmAIq0
uAJ1ew51gt6nR6/xEaFTqeUf2hwIFpcVZ1bS17yIo8bzqgwrhorjZtJu7BKRizYbcktSgoVETiJa
lJ6o2HvKL7bjcoFOQvZPgA/Pr4/FnEE7YPF7Y8EXvj8J+w1J+VH5HMWl06xTSbkrTazbMXcj9Eqw
bN4OuPvo9wocWVxgE0IxHTQ7NfXXvnQNQkRtnIi4GUk9u3lo++pjbyvFjVpg5r4LQZYlt4fpocSv
mkAfQ5MTAcCI4+RlMsd4KOtoUWuszJ/PY0++4NODaU0pVo8nk4nu0D+FRTL1MHkonRzTZtH/IKzj
SVpys7ulHSVybIuWwASW8oYy2h08CsYmZxkNze/r9J3gADA2kRfJ9tlBuRTzeuJam4+WsegzezFZ
IhEx9VtAxSL0vUOUqIn1SimcnvGfdQkn+ocqX2jdSHz55ZKquCiDU44s7Eo1YfJUzl5vs6QdA1R1
dopCc1pCPB6xn43C6xHTL3mwwXFtAr//hVYnLiUgQFaY37ZhMPRcU485BisytBcbBBsOTfP/pwRB
b+QO1kvFIvgflvAk8UXebQbILqVvIT0ZfitsZHIZ+k2xcE0Sg/SF22gCGevBnWWvkGs6TqSZBlg1
pKe6qqLAcIP2XqmnEVNaFQnf4dXYFvv6HrOM6/D6AmbPojx99I271ssnSv7QbPZnqSjDyHpC3A2F
KqQTqDtN+c8h0Ap24zqF3gc+FOpWZVBeTpImSg5W5u427oHzFP0oNPUUh3LN8Au/2nFHp/jVZdlS
1s9s2A9FMCMZ3fZYkel8UW39GJa+AmzUxZZjWh2h+F2OqpIprtQ8Zv3BiYUDD+BLIvfGUcGCj0vN
yBmJZ7l9SPmzE1cChMDyja9tEjHchc4ei8b2xUldVry7wP6Jgw9pa2UcASjxWGMOBq/gHQCuEAAp
mQToowfR17SYBm3F+rsw8j77c69mwPgkzgM8RA79AABJpTFRsBZVBYUAr42doK0Pna8UJxqdpm0Y
vMIsPY09i22MRNY74bLOM7TO1TA3gBnrf8Nrf/BzzJ5xhjpZISAKBQcVLd617h3YvqgCvzNlQJ8w
RfqApURAnkR2N5qbbBGifj4m23lt/dLCd8z72JFDRIdQsXQ76oLfXjrFJydgFrvn94fbD9AHrRAU
yo5ne7qXQe2XX3jtX0274DAZUqx5et8ihjOx7RtCjCuU7yGAGVM2VaCnHE6keg/22SuvTBzBYPp6
7TGlyR0pFFBvmGgxzL0mWpE0JfHQQfGJUZ758JHQx9Q3WoC9wf36YZMvwT8g0RhlV7hvMzpw8z94
sSTNsyO3wuosIGbwgRJfbTZgo2bFc6zoH4ksB7GYqlbfBZpDzIBAyka8MUF8ohCHtSrLcbA7vuUZ
b4LC5UptTsf/ccFHwL4L3cKxw4IWYmUeillR//aUHfZj0Avt5M04tLBnF5fjRBR8kU1QLUVlZLAw
eg/UGvXULBsqeE7NtXlHIjjBZ81eIxNCOi9LCRt2GZ1x4PwX4q8TqIwuZ74MazFB1y0Bgeg2EWNQ
IQaZRGFBXpFlWRzkW8duEj63vAHXZJcyvKfgBwW0fdwltfq4j3nDUAXnlL4F78IrFOAykUjgVIRL
v0swBF/wy92dYluBwALX8LDFlBudt/DW/kbmJxtdS9keR0AcmBHv9ffyLzF9ck9SixPZMGEcUHj5
6UCB5GWOp/xvBEZ6WrwrFntOCN7t/8MhUcIqquvP6Lt37iXkqYTS2RsZqXVO38ZZH76F1ycuXKcy
IXjwhuaCHbVq9dh9S/ze/f3oLxruYYwNBN8JPhUWBSrYyxU8CdzjtKSlNiLBglkTBOqgxqzU6omd
rsX4kub8zMoTBL66ER8/eTktq/5zRJfQ3nIJUDnMsSxXp5VXQg5qjH6aPs6HDDYTTfjT3ba53nZC
E/ld0rR3OGc2k5MDSfxd1rpQXKlT1S+WqPyRYvcNuppxtbMEvvxlVQZQewUGJxS/nwJpkVYE0Kh8
thiOLKCAT63lFWXyXIs1jnb1nUKv8YJtzRQg6YKcnZMospf8+Pi3C4JnmrQJm8TDgl8PMj6a2ZLz
zVHpQ/okVU7X/j6xgJjNiaplBe7UzAQ9t+9Fwvb9rsLO1/dn+N7I4t9yl4KiUDsHe9XLRyOQyVK6
zMNVHU3FYcSnF+Bt8kdxE+iipmrxAbuy4JJVjBRP1Hn74WAxFebh/vGQ8mp29p0FEPUAS2BfqNQl
HgJXQiJyZW8NTci2LXO3eZjAO+S23tsZjq0XDnxqNg+M3F9AYviTnZniPVe/hLBMwaqQmA8PAKoy
zjD4lg1PizL0g022h3iqB9IvHgLgX7Ptfhy4XHd2co81VQWgaJqasCGjEKkRASsk5XH9Kr6ofLuc
MVixDyDDTz+NGCnOlFWVko7/O30wwz0hUDBeR6N43zqVhO1ghwPPNexKxmXOIZArS31hG4JMV4UW
Qd+N3ucEplovzzYX9iqXEYrfnPqYplf51ugTJ0KVyB2RD6EXh0tQfxCVeYhPS4iOD8TWccuuPtEJ
SJN0r3u8oeCk1blDnJIePyFDyPua9kycFSbbPpl1DP52FDKfo+FbME5AskZN6iqBkH9kLVp7sqg8
Vhph90wHk3ds5nNClsLc0M/flHoWQ7bZM6Rh16AhZ6kxYoZfP5+9AlecoWlmkYLXRq3EfZTS8MLQ
ZSh9mc/MxvUK8lzhKdc4fpySoHi1/d5g6dTU1R7LfXLTIvg+mhhdxurK8pHk0CFcoePEfUNOn7wG
FuiTKIU2s/wh3zKwvnh6TX69ChRlOJpnoIWgtOrtgZ6JmDcrpKpUMHCUGycynE3QuWD0ZVTgb4WH
VwbVfIQIK52zG8IQmoS9akAYNQ+D8bJ9j7EJP50IS+QqHo17S1yqBcUJnVhJajVqJ3r5qUoqsQ+m
HAzPbWtyA84Jp84i1uafEOxZgz0M5cg44QiNIXNZxp9fpdwABB2V/XsJdHDF87x1/HBrPrz3+CEW
I1N/LnLX5WtB9GY0j05EXfIGReuh7ID72/wWWIUBgPegtSJWDNBn5aSggL5dtc3+WrhgRBqBkigw
pswSoRHWg/kAoQMrvDIJdFux05SnbFJ3xGQm5eK0L5pVuuJgk7CD44OZCPLL5FaSlxEWNydH8QJu
VkQqEZT/C4rq18k1pX3t/IYHMv9Oi+Ogn81VZF/2fyoz6QSEsuKhz0DdeqBmCycY0Io882xHvHix
Ko2bSLIg75u/D1hACGvcp4ua9B6F7y9jvAbv2/Q5ZAKKJQXYEvmzlPWP8s0QANQicPet99CCOQB1
5hvclgTouIgWra6vUFoX+LxhtNnSvkbYTy4KUkVTBIUfy0eWhuyEvIAVniOFQt8qnaHiq6kASwGh
fPiZ/g1vxVHz8sGTuVD4tbcD62BAUzFYWeov8ImvpBWOp3n6pIsUPjsSS060gygfymSwSuCsBRJK
C3XpzWst2NIHwbgzAG4dOhcjZTW3HC5LDjtHt1wLfx5Gvw7Ok1yUI3qhfGOKEKWxcfm1nGuzt5Cj
rmp/ml7lEB5DG8lJJI28wC8NiT0ed6pqDV0zML9R63N9jRMeqxhuk5yjxBDN+s6shPAmRH7q6Dv+
4O081206I6W34kjGiaNuytzpKBieSr5wchFQpNe2/jBskeqceejZ7jJTy1+1NJ2rU/I4ynIxRohH
BIzxcZfeIvpAs8X8h8yCdD7FJAKolZaczvJg7+2kUsA24sYjxIBDaBGuUruHNdwYCWD2IFGmZtcF
uNpcYdbgfHbIiRlazIDkAY/Uk8QyKkkK8d2w3UngugvruR1aWEIPHLWNUdICjiiDxGnKu5kHWczj
QGrRRN9xoq3Hl53o+1PpFbgUkB78jLthGQJWmoS3RvTMvG7G8QH0by0I87podKyGYsFIGy/OBVt7
uebNXnDD8g+gzFDbZHzO+ncQB8/ERKle6sSNhkSbiXEWdS2thTV0p8fc40RU7h+7K88oMWv1BKLx
i1ETBnmWpTlE5hwp/QfZIHz4kOAqQ+CJOezkoGpPu+mfF/ZwDn+H7y9wS40xzyMxt7eUiMaf2cae
0t5dTjcwvYs7E3Mw1fZR6c3jfZQ0hZOujqWQmi+JnMHfTXpIVl2Hc+FYIz/mphp2EVJv0jRKnfda
W6lkcOT6lPn3r8cwJiUhkXdVZgvCfKR3sV2Hc4AtbjU4IoC3V/M6tyIjn8Uu6akm8ryT5lzFRYu0
lAjLkgCJDzhyxcUQbMEECufMi0PsCSdfYkMSBZpnm0Gz/kCuYkHPqPh9DOkozLPdkDCbdEFT7p1J
EPKn1rylXNPqcwx6FHijx5RFe4QBgj5E/6scD42nGjaw6XMebjvebga6bDjBIUawBfMamLq3Q53R
jw3H3VzRb89RhfaUoxzSHDxTTUgr6jcB5i4ilYLddK7Lthk3G9hjkSWAzfHF4JVJEgh6RwRdfxZm
IMmcnlkWRejt1gI89pRq59XUntYyhh6vhv7iP1Hl9ZaoSpGTMtUlLYWcoGuEvNtYaLNcZmz9RlRc
BUywvA6u84gMOUFpd0Yum+sxsBjrZCpJg3bonuCnjOk8z08pTpRsTwPemGxdpZoLDgsyI6+vZlJg
/KApydI/OsU83C75xSTCH7UcdLg3sm3qPIB7hqDHS9VGzeyG5kzLQWmr+R24obCFNdIY/r2t/q4a
5KXJu1JuwoJOHcAhq5lIL3U0eqwPyRB08wDxx63ssuJyDlSOfaapQI3SElQiei4oga3OF5KkUWGd
WVAttDCSZ/q48r0z2Y7sR94oiH8SpS1/oKL6lob8ux52a0FW1BFUshd5Yi4yjwF2FDNGHby9Xdes
ztVCNgbrxikTw+nrXpFyWLgBnV/e2+Gio9uzNG7woCiY/F+v63McojQXsZRIfaXXEAnHxEivF9g4
+IjGxh7Ti3AP1AcXzvKlDeXxaw0lE3DIK9RQ7nnJImO8jSTiY3l1HJmC54tVPtSIGLUeSH9hqvo0
GaUnO/H8/f//0gcuaAFM/ty3HJ9id6iyAyE8rerkSnG6gVCqC7WZ3uD/7PX2FTz4e6p/u6Uc8Amk
9pL9sD9kXv+SFs4jHxqWP6V5/FPLQJ0XpFqGXoT/H1tED6Ctt7IFflFO2yOD7taQVi3QBA+oTOF5
sD5tP1dfK2xGFqdwhG3+J3A2xn0sjtR4PGaI3InC2RZh8AXfqau6s+I0renO9IM8m+MIEDI2pU0J
xASroIZqFV3IXk7MH8CctenRKgG+hQ6r/7rsdSqKXeTkvGSyBG4Tb9Ti7XJsTK4r27SmiGxIKmMo
wIr617blYlLNFG3SAbN+oN/nCyjpkFpoXPvaK4yDHHUKW1woUDW/3qLDqvPgQrrkhaF2ajKjdoZT
IKrsBYZIG+oWW43b3SQm5HKM0I6S86dZEZcaQdLMYDkgjg67oMY4ar/a80xuP73wJ7pHRWXeTgdH
fastTrJayM2RQ8bLA67l1mSFb4KyOzn5KtQt5cBNOwPlfb/LLfcMOcTc8kLf16jV3AgIk/4Imz9d
tT/o/qSmUvpmjCEBvzKbJ2WhVElKcT+OEkGF3fvRY3/NpCmh/Zm40nVSW0F6JqfJJuDj6SnLrmYS
i1sekxCRe3mRS0xnMtVc9PePhXXL562u/g+a8hbWxoPS9Y3c0EL3tUTrn+iDdjdbtQw27oztoB0Q
X6vxE+z1FZAV1DGW+dPrixbCmvOARqwcK9yUSPN8Q+oVhlCSNDonKehHuPpcwppak6lJZ44myQg5
hPuez7QSUHJgOspDFOfPS8QY6//pjqwgOJgqVcBk6dEyzvFVYKmYi4O0X/wRC7N8xDosD+PZI1B/
zA3Y+Gz0FauOWZNGiOrACektnBxIMl6WkR4sTAIShJOdCW2zn2WvftQ5m2adPyin9iJGqRpg+s8W
smXJUYTSO9TN1MVzipeWDFlHb3whMIEvqU5XUeZju8tZZo3f5ai4W/+I0vy+901DEOU4tFr7velY
NNKyP31DlrJ1IY/hxVwZT3QkXtRuzP4gfkO5wgt74HoDf2lGdejg9FQ0B93dEYySjjVrpKKZB03d
xQ0uYiIuaEbO6rUsLfYPJ1iGaC7FmQJEOAgTygjFk+NXkOqsJCFUjmYnAJIIxkcUp3yTpuPG2q2q
h+oAQ2IUMiB2aGUek3ZKzSWVJwDrAgC2+QRV7lPqZMy8S/Z4zU7aP6PdEnBVt0GmliFI8ZD4VM1S
/0MnXdp6gY9qkIxSg7ZFD5jk3HHO+XuBnfcLA3bgRo/Y7Pkl2tLGlIVp6wISCscUsODuVMTlHalT
LiurGAhgwHNfmpcKqzmflxy2mTQ5U6Kiw21gIeVM9V+xHVEpi7abPJrainLGuJW7FxIDDsFjdVPj
VwJAe/KqV5ETOK9Piv5bLx0L2QYoe3RojznqVwK5pRN2GzPr6ZaCVpJLL57pbExJhMrpMeA3bVd8
QO4JworuH7Qk3XFhlaHX1XVyPyWPhJypIEhJwuORG2KBMeFkINXe8MQ45LFayKWINfxB693uNckn
17eAPDKas8Rk0L7OGqvKz6eYaHHJFeY7uaUGzqxpyDZYZjoYbD7pRIVnBMMyWkz4RjHI0srRQSa5
UmN84WGJ6g02uu7HgrLksf8Y3axsOTWVFBs9jlradvtZhtWUqmLQ6I+X7YjVZtEnCedCHSKrlf9D
Byu2Sye4oGZEajb2BgRcr8bIM89VDJtlPkBNfu3fwvZuLG8llq/LcUYnSUTTcGjRE5fslrZtT6fE
F5hLWfVZuflfEkuyXzhf2HGj184mvRreZyOY+Nk3ijzGkFokyOKzOlAB4ZUa4sm4UdIoIq6C8dMO
/5qt0uxjpW5CuFNhe0HsxF9dtiZqcjk32df2d1slB0+W2ZS3MDFVMaYctXLj2UaPqr8gwks7Uipb
3y928QaXAUVmsJV37/6YWJvkO55u4KXP5idcVzKMLCMhFSCdgIDQLmBSnyIsNLl1zk+JYsu9zNsT
EANUgY+LINhIeHtiToUHstkmmurMUqwFmt5U2LHGeUJtS7Yj8ZGlj13cSd8AfWY69s88Ou53WoaI
k8w5xeuEib7ZjnuLqWqfRcW8B6DRHz+IsaK8BGxDT5KTZZdh/zTcqAlMDgFya+ViYXRXqQxUc2xe
pNlr/kcY7UU4Y5xkkP3TzExtXdedDhQ1DvAJdNOLJKhdmtqJyZit/KMVBt3xTNk50CFvZWOIGZt8
kqZiqR86tB8M4ISiuxknyHbfcNbH9p2Wa0GkK671kh87wtwFnkhUonaR5FmivvUxBW9l/iryJOmQ
Jd8w+eIXzbaOs5MFoEw1tlkZTjZMciqp06I6/M0IZxUpiCeqcQ+3pwtIsIsUrgLjqqLiz7Vj24J7
SKQQUoXfFk/kHQCPfOgqMP7czhxSe3BSp5OcNdVX299RgudgXHDodPijnadNAw2k0qNtM4HqulbH
HC18oSE/3b6qJVZsBHNDhn7eM0/1ffqXk5WeAe/c8NVcQwlYY723jGQKXnWego+xPUrQglhwVzLg
FqpSnvOIeOO+fhxi0p1+8vs0ppobBWDU7KIPZd9PKHLg5KtWDngKcwdR7QUeG4Cr3GhN5sIL8uoB
4Zh0vb8sWG3XDLQKgMoXLn9ZZdbbAYl/5X0932Kop1mxUBeFALCp9JMWaOakjLef6lVzjnLSWcfl
dN5wuBL/TzZabztlDL+AjpKHDMYr8p7sa0ypR8tef27/+eOoZ9WJ+ImcdWreb/i7ICO1QotSKXXz
gs3n3OSwTuS8q2bYi8DRUM34gpFMZ9eD4nZ1b96yrvUsb+NvOZoc/zdtksM3Ea793OCoBQnQ7d7j
I2RP4bKOKZPdUZ5lk9pzc5IYki+GIyn3AMEE6LLXEyvHgsa4rqsLjvRLgfxxUlD1sG22YIvIcn7u
JgtsffCkcXoeEoTPMPQTnwoCaKhaoGIIllee3hcfLG6B5sLckngU/YhfF9t26x5doCyLjCmJmglz
FP76vjDg9epXH7TREJx11Samgz28lcZLVaPvciQO3UY8rfjQkudMVEZk/tUg8tF+/DuEvX75srFR
TzQT9slTtXa6dZvnHtfDzg1SqMgIdTXfJ9MoWML8PQxR6hOqSAargUUuXWHhGjvUkOdRExJ8wxp8
loxerasYSNAigxxMY8kfRY2r4W+rPNI/woKWBKeVbrnlg9zpURG3qtwGrnz2yuKHGGd+167cgdSr
x7PN0cBqFnqJrKR0BhtThW7DGivZ1377cVQ0XYckdxIQkaeNaVclHTTP5+OYhOgwkNm0J3ybL2G9
TMltCJrsQm23545jGnig+gq1Zc5aEM+z3SaZXLiaHvhOny9PaMzhR+Lsf7qOjFvt6QD3Av9hLURV
aCdISOvUPc0hpgyCbohfbM7vNVNuxXn1Nwh55sRcT3RCLgj3ztKNb3aPiSFYXbssAQqSUrNWFtUC
c8Zsx+Yulmg8C38oi/TTOi7689PzfloI2yIyMoUEFuHk1U8WbUWcKaT7J/d/edgEXUTioQq5a7Av
k+M96F3wx8Sn2TVsSG7DaU8+Fa5oENvPfwhIMc4kd6DHO1j/7xXglmINUYBb02HcM7+XFuW8r2Gy
ZJDbqwLkv421+GVkA48VpqE3pQspuRzkYeLnIHiS5EOSMjjwif8XOj9SBl7uK456yg3hb1/udCja
ovVxdHVWZXeC1/YlqgjTe8KhXk3VwF7SqPsCixje/T2DgLHI5Hb/Yi1jLr1ocY1sDoxQh3nR7hhX
6e1vBRhu/AVdPUC49s9LNyYkabMLmZc6TW7UcU2aMnBkfFaUBqICTGayB+dggRkoFOkqCr0VE9mb
eLpSCiTWzj858dueLAAZvJYjYwoVVXwBPErnyg5uYjKQ1q/VDUdfw5BJxFfPviOCmYrjropUHd0q
Xdnv8AfDZ5mMbFgCCcJQxtalOs/P6bvxxoxxiO7sReUExSB3ndod8trKLay9qhFNbpp7RIZT6rqD
zflEMRjlGkRw2tjkB+TL8+96STrBL3NdT9eeImnRHZ70d3nqSwuvwjzqn7fDGk1Vd5R0M4XedyQP
nkcOsZej9ifaxSi9fDd9FoGdxPyARzT/Xm90NC2CVoEj6Uvr6YKyDd7xMN9NrFeJlr0RQUgh5m63
h139QvV2T6EHNBSX5t4LbiqlqOFDfd9FKe9m4gI2/m0ZPGpZUHAcHYe1vs530gZq1JepYDVI4RtY
OqM1MeOQowOFykIN3yDeeJf9vq3kCAKe61rhW+MovXs1Os0pynpTzlVbkeq7JydUdf1ild10RWas
LvNGBmJAl/YupCRNjfQ1f+xgDg6Rcmq2niJhFBbR717/5VEP5K5De6ioti+oDmgoPHc774F4uwZu
qc+5Wa+PyatV99D+iuedvnGTNl8S30zxa7wJCKrLzJAq6zLMTxPOSTOU0cYLlpw9Njrg91/xYJtu
rAqoPcMUQcZ2Kw6D9SCeU6PJIHIXhvpYgpujQp4uuWY1tnyx7vCgKVWB/DqOujyn62/tIY8ug5kY
HFv2fQyGfv9ytXmHIvyJDWXwnTq1i0s33NfpINI5P2vSuP+y20F172JEg0ipODPRkzdTzntkByUR
7QHvzHu72wkKo+nGULlhvQusp8YRlLiLLmxBykQShv8Ip9zc95iEB7mfchiGw7EvDFKhGeXCDFv8
Mei4CEANO7VEk+pHNWpJXXaWYj8TJli/nY6kznDdSgPdCNsy/GusntnCnAp9YvyNh15q/2J6SsEP
Movs1rdCVr7EwlCGIXzzYTOTwSUm7oKrdlvTkKZH6Eki+Ty/wg6z4xzHcEnfHhFKtH+n7Scmhv6Y
5XzPj0f1TjnUVx/baEqUxGRubtD7ZfoU22kFYryYRcTXTGNcQbebzLP1s8ZEZj2/ltuRxx7iLlKy
8BjP3+VuGkNc/PJttz0CGELs6BGnCsMEqLfcW+ZhyDs/QaVzuOe3J8VLNZn4avmIOof3yFnohY7G
ba+tKFpvPz/2Mc50lY8zrORMJxbkkn9uSq2g7PvZPIHPxTCftZxFuq9kdSQh98p4cMiyy7QmW6y5
vD5S3Ys6VtdeAu+8zGnEdIe/si7XrmeRblUsLYevmXPqRp/NCvQDzsb1jkF2JUsOINRTWnG0QW0M
Mj28aeTchirPPbzT7WhmbH+6opEztBq7KqWxJBEsCJWSi6B+PY+wyhe1G2ZNZCFHcpJyKhCdJFpp
IT07vrcdWpwb+60LxmWdQ/iEb7bDp92q4qkdGTQPPOjoCViXk0tLB/njhLFRqInBVFdpq9v0UdVx
C/XRvMQZLlx1YAMSuW7hQNz8aP+7kgWHRIBaCQ3qGnM60f6QJA+VuaI5jtcKGH79MvJhgx5FkIQs
ytawtfjjbJn8M/wMEq395FNaGs98YMmaJp2p92fsVvzepsk8j5YxZS7oUzQ/ckSZpFQic368/An9
JZnZXdvJfZg6tZRbDT/azVmk08ItNc9PoEHagL4m2rAIR+op6SU+rHmwiA66vavuTbG+xsSojva1
6ghr/aSfiICkNsjEvU+BqSJsRn1uD8LA7mCr1ufrNbspZytTn3T0LSgj1q5HxH6GBkKij4U7q7Dk
y7bYWGPNAd8H3RH/LJWQ/uGHZWIT1ExZgORVigFnO+mxrL6bNGpnR16Bkcrs77vPtIP/ymRMWY18
OcNU+DZ4wfiqE5SR6rU7S1o8wiVPuCKDjxj6xOVL40AmRMHWPYeFiVgEAFEK/MzoiNG1z0jQ3+Xm
twh05EWQ8FyM2Ek92HL1URtjPJdL+LwJQu/sDEk9YzkGQLk3E6/oitCHBm8PJM1ze1hD5u4IA2Oa
QaehAZ3kC/7Tb0OTumzTCH0K8V6jo5n3kgWqJGV5MyN8Vz2vMkC9bm6pCehTJBG76e5jx4eaYDcz
933V1bZrnV91naGiQRnTTpkLlnukiX1KBtnxoRByNMoEKReqjmHZDe9o3CeH+r5UzIDZBW1Qa5aJ
Pw42PibHDCORDhy6XIw76xAAMkCaUdd6uwavA1OsnahRXqrVaRFBz1VExB7ff9FEEmclSb42Ub/j
e2U0AjulTsN+n2cjSFJ9frWy/w6wQfeFlFGFCSUG9i1drIXPleYSBXVLYwObx4GxA8ZqmqFTmuQ7
2vQnIB6clLKBItHbzy6S7xqjsq4r7MAZIna0IttQ4jQMwFtoheyY+SU3DE/3hlnl7t1lzKiDs3cF
bpTeaFh4vLEuXygbztfiNpou8OLF5nZS08ws58zwvid8ue7AFTWE4Acw/YrjClUBQ1s8FxIix8E2
Ue3C/nVjCLAxWaC/ZFjjruoE6z4x8NDEt05LzRRrcu83PRzo0doaPeTrdrWvKpajO8DyzgBEZTyj
47JrRfzY6OpuFcn0wAxIaIDfiQnfAQP1R2WRTmfztPEnrKv7KGazcANIl0RHf3fOyOgYWtzyUVpe
IdZZwM6o4VaLpyKDro5zHzoy3ipAo0yk/3bxiSZa/QPPPvvmdqc8Yo2hMai3+0Hg2u5ipDC/LZAy
svKLF5HxMnjlpPiUaJueaWPKV6O5LY7Giv4JLSS2Azr6pkmMGFmHI8c48g6dJajNBIcS7eYKQQL8
2rrzgpNRMFQc+j7wL4YMxpBm0IamZsYolQ5rU2tScfmlDcKic486Ku01a3m9k+CAYXRpP/wgwLJ4
27L7RJ2jOsYXbAh31Ghjnnf2H7ybs4w2C6aHtll6xcZ0BUJges+0BFjkKfVEKvNSwAx0OJOSuO9h
gb+Lb1FPfV122EbGc52Ds5/0sqLNNtu0i0LssneOqP8ZrMe60zs7iKBNLS3u+EoJ7P+ujS1lpl0Q
rc3GhM2Et9J14Uv/iONJDEMVXHhtM5+zofwpathHTALi/BhI15Py5NrDwwTyMKKhshR3kzyP+dUa
Nc3vXm1EAO1VKSs0Df1Kl3lV59hrcLDoqi2DSXEzvAL3WL9acxvNcOu9ofcT2TZ+gY9mQBHFn8/P
/T46yD8WD2hYBqgXOUjee6lX0uwEw31SGqZZ7VLlcvpP1aVRB4faf+Lr7T5X/Bercc+QHo3aOJeU
PgipsXd3E4M4E6/ErK71mZ9IXo44VjoakN0KXXlmvVu0Nlr7otdpUQEH1rPuBDglVGHIL2AV1d96
QfqRXl5/X6VuQDPAbyCV5WvJy5SZcaE6bqNKr1/BbJPlBlUsl1LAl5nZJPZAfWtyBJCOwrk9If2t
BezpP2EetANKfdYBaJqe22gnNRDF61uHaSHAHDihivRa6k5Sa5raZcpq9AcMmDHaFiDEyGbnbROo
b/ahEGQ3ZUjq4Aa6Gjrhood0ABGn4e93WuLS9vb11a4G148rkS7MnAdnZ/c7Hs1CsBjTVGpQwbBp
PBzBCqJntGH/uKr916yuJVMyGG99QMeQe9VnVV4Sv8xhyxA6jnf3mKK/GgNrLbpYLTHjvP2OOwRk
9SI3kJHlzN9yzwEe8Xscn1fxUv9FZeCVO89L7/rKiN/GkBeOdMEPr5pPY+4SE+OIun2Wx5hhwi2s
3XhhdHxgEqlDrQhJq95nm3KIG+70hDew3fPH6PA3Tdl1ihUB/fUu5cEEo95yTz/z8eY4zIdBLxXt
jPp7e+jHxXEvKn1Bc/Yt2DdTC+XuRMYKiTMMq7HuPcPGW8IiH95bJUoRIasph3m7TsuTvhp6YO6L
JTMYv+GEJ18Oi68SAO2hYNwnmLQiCASNquLtGh9tmqsrFQyW6bPB0KKvGYg0LqrRaUUaqMFNiWzO
dUeQf0pGfxrK5XLOObSIwGCmzk9Q0qCqpoWEyzm8FOFXFBO6SETxLL2g1QwTE1kc1SuWKCJLaarP
UnypK9f4nDiFSkyB6tboiWjzJaH2SM1vAEeVuKHsnL2M+FXZMnz8Crrb0DcIAMeVteuFqfpCNhQy
ErOj6/d2HJZVbhUFbqi0FdwAXQ5+V8OZ69uiioJBoiKo3tOz3S2swiyMP7KGd2geXEGxD7Z9ia5r
3yV8+NrXobjUx9GbsIh0hqGvFXEs6NnbSpXLW+qgzuxL+jM32xuxh3v3kUvmWHmKOQLSOb8IyWbD
kx95cFt0hCwrMdfxn5oNsNUsekd/Uhh229owUeSHxcmUAWgZD+voyfP7uBAyQRcOtQ3RWM8L8aeO
3r7nOtZ2Xh07BV4kP8+tB6HL4xKKb8A2M+d/drOOptYIGk4YEdst3ldz1gXVk5YDVAFz23T5LJIC
3N7dKpwks889VhL0mR/oMU2fXChredFXQiB2aKU7mJyNZnWXXmE1dYNBXSiyUbpuvk3Z3Jg6SC7S
nCyUlgjFRfh2NwPy/hM/vcwa+4BLpW21d7FVCPV0orooJl6fAyk4KvN2Rs5md/srgFRzb3n3n+gm
7r2lJibPqod9rblckwDCbN2QKYwsLno3ulCedCdfFCUeH3zYKBXeBXYGl+/w118oRlXI5Y/kwrwp
JROUJnjJSBaoECFPAy7OscpfLmL1HbvaVTqdBIJCNQbxPGdHdfFvnLHaL6posgCmke8D3HinCgzR
Osv50wBvXQ4gi7qHtMsSw8M2mM8V8EjyqR9TrtBd1RchH4ZyKs1rfMwjRHzLT6LNBd8oiWgbLBFh
u69XuVTRADV2yC6Nscru9EeQ8NYNnhzM3rAp/bMDx953Iy0wFdSlGkukg2Sim+lk9C2ALrhgY9wo
xMg7nZnhN3pifxGEiigB3ypKhOH1MCAuVkg84gCqYoF1zLIErRXRNbA+WUy/EVyUNp8wA7ghped2
EwbO8oRYRblkeigRXag33qYyM/5jyc9bmEHVj4IYQspGZATvMO8jrykznambFElt+BOwm2e/t9GI
QUdOVbaFd4Lf9Ahg5bpEvBYwqN7rC9om+xsvOIa+/xA8AP8eHMFQdnwxzxCIV9zyV5H/n7SYaM1i
+VvQDqU6kIfDqs/XDU0+6fuaKWDvUyXtGBzFMWQkjCehDEC4SOYDdibVDnSFX/Z9yw7RWxuhYlpR
4M9uPPpAfotwLiugWLgAnHa4rxVINCTRlVA4ejunsyOImWQ4Q7iPLN+FbEmPhRKJC2vnbj0myCFd
mUw/pUhAZgSqyNCrXmYlZENGlgEBRZR73GQUYO3rKEz2Hur8PW994LLaQytlaSg+Gh+xcZR62PnR
KuS+prcjeSKVOWTWK/mGqzRacIeboQ2eVoiZdaF5MMOs7IYTEkomnftNn3sqhFKJZQY/gx+X7t/W
6IJ2EYyCk3vll6y928btL+WFeeXKqEtb8en8jU8gfWja2yXxAcCy6n7rrr5ieyoK7HDs7pyfjq8/
9O8MTSPY7AtIQ6wHkM0r6oLBA2a2Jyye6m1cXMeciKRp3smMKx1Cu5En4DA/pm1oLvz91BWPPf3L
5rbpDMR6RkdFJXJlVi6ZTAOTbwLvYW5JOk+Luf0lyF/VjxW4pR/jOliE/pOjpPUMmzyNpQqlvBLa
Zj5lTc4Fv9I/UvTBych2/46tlQHJlFXXIzVt3V8LdoektS+/pKcBSjSVmq+IfqO8x0Wf3LiAxjHA
dtvxEc15mcSRG0m/TpdyvJjKy0y2bvVWY/7CHKAOsOwFhj8sLH3MJhcqTvwvPmkIPVNLQFmTiVvW
QxNx3qCjndBvEbrC0mjBnNRwr/RIclyX6mulIfQkAl/k9AOTPjkLPEDuxZmb5IrrFOqRKlCkngNP
CzgB577A+NxJ11fByNFNleu3VcKh5xl03yEKNkHL7FW8vIywnxm0S2wO4hyxy+qz+0w2v6nEcGMe
nFOgemSXMOV+pI56OAglb0z/xC9S3SnqksR1Bpp8ZDQeMEX10LdSAjRSK9U/HInm9nObBu/AtvVQ
aM2u6NDZwY/OiAoksbP43iDexlLETrS+N6pfd/lkTPi4FE+jVzdV2V2mK5G6yNM58SLYi9KkrdoG
R5mOTJrD152f+0vUgvZnadIKFiPfMYNA89YjBECPvFQ2gheey1dMQ/IK2dD5kvSZJ6Ufs/TY0Xjw
SdZulMihAxX6KeMNxKpGxWmlfPmr2umA1qe0qPkbcLlKv/SrnBdMYUsHU3d9oUnqJriFI2fyuiaJ
YtHYuthvHlaWxImsGS73ksAXDpJhZ2hODy9VcK72TJljdPOkGMynFzv6qi3jC+3wZQ1bEgnIaUvv
GYUQxfe09K+LBXuY0f2C5aN4jQrVdT2eRaxFblLrbojLqbfZpkOBBKdgRqJD6jOxJMN+Gd+VSNen
Zk9GotlL3aZIv4crPA+yOnkQ8rClO3bIF5ZYgEO0Koa+hDnsKSyIlOrK/55DQxNCPjGJUjakEJna
eSlKvBVPqP2d9UlA+3jE4fqImVn3reaGFf149T3lwGUjWrar9KRBuAIxHotERmzKOv4A+Fn8agaM
FB4dwzUTKUh6Pw4CpwcbQaDZtekmZyDFXobGkJ8Lft/MgtA/TIlIdvbnxk9AaCfoUUQ8OSls6NO4
f3TG0bNwbWBcXSkLTcRu7FW/6bMNLGpRuhYHctCVQVFwxCxJMuQJxL6pMhbXze5+jvMr8wjB87pH
E8g7Aksw00ygCW/4TZ3DubU8wZ4DvAseH5YaQ5sdO50jIGqz6y2lx5wDKrUKrhtruCutU3to3mul
9Ig1EC9J3O2dEEowTgpecCGRbBrQA6HVh/J8galq8rsweWQ9w528glWTLDamXz2r6BC16G6DOj6I
PoJ9AngBznOc1tOOeh1OLfMK/mj5u0Pi9VB4ASRrPH1Ga5HWZ1r3ail2x/BKz78+B2L051alIL0v
O6UiZQ3aUiwn2TTBJuxPxalDywEVZAashze6sqrWDYbWl+ls63gf8Hlg5yQ3Nuen+dzqB7HrlvZ2
rn6oX1BdWMXeMx/+d4F/uWK6yrmgl2J4FkwdkYEetr/GvKU/S9yNFvPzMplOzTU/cFxVtJbVmvj9
hvBeXMfjwiWD5jriX0a4v1LGDXEO6mStKrhefnPTz1xWHEM+kL0nklsM6Y7DuiFBolStoSzg9DE4
voCpl4ot94bdc9tDiSMdTjk+JGWjZzI+mIPUT13FBaHUuRhgqG5VeZ8rAcl61AQJFAFGPVWbWOWT
KDjSxnuNxLjtRwiBg5PozStzfLUnVHOU3lmWOhyjM2xcvdVgnAdHlz59+EGpdW7f2IfVHTipzoaY
NFMdwGhNJTY+75pw78p75YsOg3S6GFMIhAXrZC+Q9+zQMamtfYidwAVY2eHpC8brajz7OxLtyGdz
bmjVNfOhIV3ackHQX4o+G39QJz1Ie0rwu4qtI2X456xbYQXEC+Co4mgt8m8JcYjVxjtOiAFIQr0x
ciaivgWXcwjn3yGqu11GS/SLHTEY+7xQbFwiP8QKm1nkd7I2fzlH1MLyDh1RdxHU4wu9Yj9ntuYX
u5LhrXU0KFC66VlRc45GbSjFnboGqpipkd7BtK7aR7pjj0eWSmzQLyYTDjn8EcSSe4KWWHOjoisd
73XgGlf8ib/3gaNRhElzj5V5LPD3PlnbwmCAiJuzZ3HLnB/OUfRipHOv9v2+FDfnMb++dtYlOEis
d1RO0AGV0qzsF1Sn4bQq1S7kcEt3h6alNBLPHAX40qTzhGilNCwo5LUdaao8qzNdLGTzt4FCMlTh
uXA8E2McabFUWdz6kiXUpmbcaQGr8CUYRVW3X98EL9WbhpMZMW030jQYvm7Gk3n6053S2hohfebh
Ym/P5cfuuWaboD9gmCuqPdIKqPUwwASQUpjmWrsJXxMvePdecDq4E0qhXA53JTZK6Iz08cXTpr5W
oPhFUra8LclRUmDETPsQ5M3OFv315pomkx1mgTlRNNUPlg/i09qymLngphRJguHaBPvXZLidMTX7
6LhaUbyr2/YEIjfHdRDO+9Uzytf88Ydw9fmz7zIf8zTw1bfUiDciV+Zc4wdduHTQGx4PekRLuxAX
hpLA3aFMG50bGFNOUuD/3xi5p3rUu+/9eb6k5pEFs7LLkVHLIoSjZhxirPExFzagJu91r6viYKW8
gy99FfsNVxOaVWo7AGLVCIGPnjH1cEUq2WZacOAsV9Ax0vwf8Oj7QrMKuol5nYsXdSOkL1qgF6Be
8dTUYU9885DkV6s/Vpje1j8p0FFip/713KG/N22pkqa6S8+2lB+XngE7tUDrtMONIBGnyvL6/A1a
YAxrNm5/smHKIJ49162zZJAPdUrU0eGB/HC8AteD+iw/Ig1Xyv9AroS3QfNVB5eozZVMTJgzEkVd
B+9qlFmYy5f/iut2ieiC75gDQS8mQKFnrYQsNBi30iwan9OtqdytZV7mzEqU1ajtBsxQkeq6OlfQ
MdRsBZX4O6pppjLy6/h2G+XYxEIAGDWQ/MS5R5p3HVe2fKqvdCiZ0PzyZANznI5gXmR20Qh7D3NX
qP4G2n8srJZaJZMqoEbomAl5sQ0nfjbVJOh5RrsCrOXDKaFNZBAlKAz32VvVYGVhC5L2XVpXsOzB
xi0m13fJwEefjAuvzN44Epyfq3MrZqU9U3GWvLGaa4brdcwrCxvNorGypxoHJmFBFqTF7kMlbk3P
ghifUz1U5lLV2qTn/2PIB+qAnkMSCqvM2CRC0S7DHiXNq/9EtG4H8V1Z4t0QAiT4hpt6poHN4Yhi
ff6+LwhDeLItq0H2wUW2JIgDHlVM+61IwlJVy47URtPPdjqwN1FuOBzGWpo7cIxkxq7Y/1q5TEP3
XYl+AiBTMgNJiercFKMKyyVlNiQ5CNZoZ1Q347g7/ZhPBni1YQ+p7ctxqYo2WZKSF16Y0Yrk9vnI
TLt079JbC+88YlTpIB9ERT7LK+sxcRXpX/RE8PL11uFr5tMGieCjaz6UIeTze4uzanHlk24oR+55
hf8cONtmGzb9tSQ4a0y3sYjQwK5QuojtRYW9vCz2nEY8lmw4mg9dVF8Cgwhu8las9kmpUcUwOiyf
Mm5QgJEUIXwAbE5YVrOa0J+mdRDWIY4q81y6bUNxeScUbOVqORDv+qe7jw6rJrYnQ9HutLCiwk0A
hbKmvOQgQ1EaFEKjC4mPAUJ7DK17MSAX1ygjLccZV0YYMA4Y18qmOzMfT5j6rOZUX114NMHP9+Ar
PhiszfC4datRwGsmdJvV7dZScpUHay43GsqUa+jEMmpeJlSFNf1gI/CVZHbyOFdbB7u9dl4Ugmmj
Pqkh3wC8Zoi+SEnHmv3u/Mw81Zm2vJWsd4R10sbRXdrwz/WgCJ9if16dirixwIhGSA9a/o78TJjz
kkrTnGCqsi3ahZkYpzoqm9gzhS2fL1RT1+KL6lRG+C5CyATtCyIv54oXLc7s1dQsLNLe0r84TAQb
pda+1baEeP0qYcAztRVoUXOlzShr0J/KSVA7mZo1REo8vRJN0WlhZzf3PCPJX4A0dawNe1wTKxVm
LGMc0Tw/kWua28GICm3YBl4WElkBp0+hKA2kXNcJN1/iu573r9IwrtxW+n6vDz4nKwOoHYhuLb9s
2qA0Zwzflv0WLys24pJX6ZM+m+/TbItHw3ffM86FyhfykSUce5/m1KsjCm7uMdAnlULVJR6Twz12
61QzhdOmpJz3FlECoSsdQOSwQpxMcKjyvxr+oiMOImcqnpNtMseepNk/kiQ0ytAnrHZLWVZTbKc7
i1GA93G2lDSPoVu9qdT/0VqP3GcQVKU++3nZzgK4qhYrssf/SCVrn/VwWD8HRlbCEiqDdr7M6Y9W
6u5x39yCcWmyFW+kevoL207IH/RzHShYv3dzTJ70fWlszLlZc3Uy9XyzlEqUiRkWkU03H2anFNP4
SqocjbmzVz7KYSM5IuDCPIqb7tFeNpHXCwn0iieVQmWhQWqCC4av6BqTkkheU/bfiZTFJax7hjCk
epQAQR6m4cB2nnZGqbVL4TEoJ6Zm94kHej0Cogt3D+ETd4rs2jjXKd0w+/CswS4futLQuvKNZd3c
vXIgqQXyH6MsHNb/i957sxLgFXWMvC0bZoSS1wc7bT5nM8QTs+cvJkj4RqBpqMCSa4l/P8WrkezQ
+m9hvrswjHY62wAX5ORUpPq9CwfQIUpwDefaUBSPHf+crjExLEY4xhwe1gxgfoLtqXIG7ZO0aAuy
GuVm0+EPIOJZlmMgK+/3b2VYJxKfUbTAgmz14FKWxZUjVT6Aa8OnkRKEY7DZFPQeBy6cwlQQ8fPw
AOj23KjKn0iT7KbcEM/MTdbcIowGYrJ8VQ8KVn9hSNh/xaaPuMGFiMJc6D4sGoysbsOsJLzmF6ti
Nr2Zt/W4cVQNcSCYxw8LGKgwZGFPiPMie+F2IkdvXhmN8ZrpQClu6vgIl5VrM00vKuJzWbZe2WFQ
cmt1ke2IcqpD+ITcJmOzGUmJsbwCRJjOkMe1m8pub8ei1OKrUsoOM+CMKHBXsD5MSY6xneN/yr/y
WcdccmlsV8GFNrNUKitLyXJCojjT6daASWGmNi703vWn+hUk5g3htH11SOeY0KtXE0Eg0pXu0b9v
gB4LU1F5LS2HxqMCMYzBOQbExfvH/btYbqN/emcGsy0yLdrfhXtrMjA9OxayIcPczvTwbjUWxAfu
bacUHnSw/XY7ZsSExEmYTJLZYguueqwc4qAGT+DuzvOLxjjnkntj9XvWTPqwKCsRquNlU3j+UlHf
rzDyCidpe4hsMqGMAwZ2PoXIx7oi0XQyPBxTPN1svSRNJyjrt8kZiIsTe37cGTpSs/pIm3Xjfbqv
ypJwaLjJPdvFoOjcrfCoxYojO9u4KQ6FifrKEL4BeggjSzEhWAu1AIserCtEXjFEu7PERNsANgN5
/sD3eOeTbdFogJluzpDwlXMCN57KV21FrEIFYU8V9qjI9Vy5Ik5dHPo7JvyIEyCVQOIU7aEnlNJb
cOodq5BOqHBarPNEDkzxdL7zUNaNMPbdmN+jFm91/azQ0SbajQ8xe4cZOoOhpJKobxjksEHCmITT
Dqi2/2IR7EFrHkvZC86ECeuji0BWwhHqcZ5K3ZEnDETx1pOKGw7GJwcnkfcm4MnD/7FMjkOFW7Pv
LGnuGIsfyCnFlxBRcDc6YDwcgtS1kq0L5KIvoHRCx0yarND68PK+ev4Uuh09KZAyRjLVkLXFEEfp
Q/nUJwtHdCvcvYE2dy20cpc9/rSi0NNbsJVdqIDRyooupMi+wrwRoImrIklciKIr2KGVk0gwOt08
6BGQMpN9PRNWZzudXCe6MUD0q/62yyZhSXvpH+PO/DjUUMezPmcHhzp4yG3dfyq3ggBgwMZjvuOy
cqJzs8aBUU1hWzX3Wg6wKmFWn1l+8K8SRKuYQ9pGVmpCNTExZ39i6oHa7NlQl/D0j1hNvHxWRq7c
Far2lx/uZRYapVY5iALBMq130Hk7ewx7I0FEii5Y3eVAqnXcHSv0qu7nBaG9vzg0RyJkUPX9Foet
ZjVuNeq01iflTrCBVOAepZJfwnau2Uhwq1bvjj9bk2OsIezQd3GKNkWJkgd7jiwhebOapvFz++n8
9Mt4OOCaVKSe1vzVhztiOxw8pSHHomMrXcqb1cvXU9p2uDtKf2Uu2bah7u6nRl+Xf3q7DpW5GEiy
0p4C1FhF97zTf/WT/Y+coIb8IdZuWZV3aqVvp4HKwDq4C6r41KPJ+yAID4/iRo6pb0ul1DVMiym6
UK+uYshwztjWL5GrBWXLIARVpeLI/SzA8ArfUUpqgK2nQ9gffzE/Wa3JPmj9BcqhWzJaK8/F05dk
VgCPJ1D79oTOQ1izYzSHZOXlSqPJKC3cvR3li9zOOKeUP+ZsFktoUQxPCgIky4twTxXL58R1YJxa
Z93Hwlt5h5dcVv9+M+WNEBjVxx8aO1Jt4nVty2bUgAA6tb/RKgoAMr+thf9a9xOUlYY1xnhGxgic
BhIgp6cj1jWsed3oA6SRaJYqstndee63k7fjP/v+khn6K7v18zH5yCthc85CW2J1sw9qTCNMybpT
tRWben1byXqX/LB2FyvAbE4yKPCGib5LS+ekN/tjQK9Y+BrQNbowYxjCn/4quTBcyZJzSR52vP/c
1d5SDH3Y+SRClR2Yw4tVx1T8kRDU60mp7Y7gQPigY/+vGp+lXC5peTACVJxLxF7Z9fpL82NIPQjG
qQd22cwgak2Ahj712h2ExtyZZwf4FA15rD6syhRTwu3zTEDjT6Bxcr64UxT5TLPXTRFOQo0oO0Mw
YQru0HMPwPnRkIudMOeynj32O5iEFO2eXpz6be8JQ0rxbWYVHhvhMryh26Man0cp6vu8BQxF6Omc
l6vtd0Kkis/nUOkpm1EoXVrFaQOytyhHGNQFI63PcP5xZa/w64Ec1u97jJ4nCdsNGbh5kQycsIKQ
W+0Bcq267XcZf0hRgWf3daGd2+0G9gW6129/NKiqhS1FDpWNcqcclbIuV7U9DnBSem8DLdbTB9dz
2Ao1N2xqnR3zt8RKITp7z5Tcz7nAr0HRKEXCcEN66dy76BeLpkFN6wzHn1ItKj96jSun12QqjygI
bIqQrJEigjmtgPx8ceGgvuWsVbdd6PIc/Y2R8prDR8NhMyCEmpcWawtFeYjJ0GpPOQP4mQ+4kbuz
A1WUf7NOyp97VszB59e+DseW/DubEg5SelMb+p/VSlGy7ApIJYoIw83Nj8pAxwLRYO8/jwvxAnK/
SA/YMdBvUUY9/QbgWqKqxkKW6PZvDZ9ClZG9ZqEhhfYEmVu8uAr1wAVkj9qOnbgxiY3mJOgmQ5ZR
Gp8WIgl4zlvaJzSb7+mK9dTx9qENlKZPpH8cuFqdWfuEo6bSC9Zz9Opp9vRQUC5gghpmRmgJXYCs
dYoiW6dnnRh8ITbUiA/BvWi4PMvDZAWU2cK55mj2ym/UOUvUOV9Tq+4uHjZnJin4piSoZh2qUK9p
jq3pHbXlcpE6gheOURYnVWY+C0J3itEc2DjpfUhoItl3Cpwg6lKL6VLbBSpbUu8EMT1FUCGD+kzR
UZOvTx4z8dlGS0fOUa/ZGkfmO1C/R6QXsm4gJ2jUWP5GkqWJmNCFOdNIeoGs+bLR2Bxh1bUOGwla
j3a1OWTRM+bxhXyeAGzEOkBqJEIMGzHnkWUkWm55spM7Ll7Nmxo5YYmoTxqN/Xp/pAUAsCn+fwKh
c2rYBqtWR3ToCJFoKObfTBwE3O7D2ybx+KAjOER7TbzwvPCRvB3RgK7I1QoP1jDZdYgxnrlGj0p0
tPXs0I+j6SfMan1wA3FXb/zinsXqGugTJW35SFMetoJlwp8lsJeOmzoMab97x4yslx0k/FtWiVyv
+/gYRhUrfJp6y4CwE+VAr3YMt79LiuKVT7wucSVIPBYRSa+KMmyFKWR9gbqpUof+bccOIe8vH5nw
gHbzG/1klRzWr8I4i7aGIK4FG5apdmairtC+ynF0eGO23PQvEKph2rsDEpYCJjPonSdlDXG/Ip/I
+TsCCAU4aLGDAR1hAV4HG15ssOTe1Q1h25CmZ2tfLz5sN2c8jNeGIEum7erpBLfbn1Rf4emFWKqg
+CDRmf3sdrWqRGh44W4bKV6XHb0d5PPCGx0Sr0/KJftsP70TUWVc5xni424G+wFkw0M5Ti8X5LL5
XTMXaShEHV4WJ8DD70mJRarXG7cLGt/7fgXQbc4/4622zGfBNkbgghVr4y0hbPzwY7IIdju88+NF
Jjuh5mdXmUTZEQBP4pn5ld5vI21nZA5cpr2E5GjU5Yg6nTxKwNqqOgKvWtvuKoIvyW1fG0sFP9VH
sc2j+Nq7IuH/wVnbkLfsK6JMKWVtZHuxDc16Dp5SyoHolKy8fIFXy+N2+oj7Y0Q7pALx8RJw1eQF
4u1iTAs7YQ+pNzx1MMJExUjKqLuvhDzWQUfJbdno9rFMdikKovMO7Wtc2kic+xJEixc2zR4K8q3U
U1ckR0xBFLXnBSC7ZGalxr8DuNzQX7WRXueNftOnma5B+ttb8qUMybCpmAvx6dvn7u9Sqbhh3QoD
UDeKVEG/vM8ScuukG/8EV836sG1eC0+HQyIzUxh1rNxnwessDjSWjJlyOp2BfIU3A7N8zHp6aIH/
htjcM8kQPkUhfLai65vpU3l9Wwv2UOebIK20EpyWiwt4rg9xYgCqzVw1HmnbkaB6tftYYntP6n5c
3Bxt3ZbLineJQEfXFJY0+W5p6yuuc+gANDs+aOJZIBL2Xbe9KKbLqbI+xhzWTUjv5odidorMlvmf
2/zDdQ6DwQFNGqcwVvU0sSKQNj12IRY4oKCt+GLNJz4fdB22ZbyYfbTnpHEBtERPZSLfthbU5j4b
EXxqRHCfN8haabdYfFCWSpz1ceazXf+Ol3+4LEc4ccDhuW4+4ukg4rnbcn8Ai0zfC1nilzrpmvS8
0G5Ce26tssMpffLPa6LMtwveOhIZI9gRUNmkxSrxUoqVbdIK8k192lHo+Q3lpcwCaMGsFSuvm7Gg
z8OvwiEvoreb4Q7+32X9oL7sRgQ3TjvNaiwqAjZHwC5O0JZzS57OQxvV66uQVEaPV+4FqjmRSwss
m3lhG7PUT2nTh8d05xhaivsV5PINjlS0WDK5UX96L2grN3iN/KNjdepQHbpWIJm3dj31fa5a6RkT
M45hrThIaN/7Ql+S7C5Kdq06bYT6RNPRnEd1o44u4eXVYXpg3M9jCvG0qhRTa5IQpwFnmVrouxBp
iScp+m1lRLD4lzWI0NNachRhnmbBZM7dHvUWS/B+HSA3q+4NbkFSdMEweyPz1lidE4Q8kqjZxB5b
/c6XnItzfcdu4+CnYobpi9BHtOY8zgEpzx3gIGWShEC/N6ByG9Gk+9JdGL2RowWrfD5STbLrA8rj
TvQxA5oiQiHCyVeOaWAtG6CN7JQOt9kBBVz+zv7o+GbV4iQPqDXYpVOkUst/6S1CepoWO6DSRpbr
U8q3wzjhMSvwTzlRl8RmBd0xkzHUJq8j386kAzrbSt6ZSvCnCX2kB+yttdil0S1pjzZpUYC2wcO/
cEMIzHfvt815+z42bqxO1lp/km9Z9MrB6SK6WIS0+SIb4NScsgdl4+BtwuFvUBAYaXeLRAowJQ5m
17BntVIXLv9ZbEXtSXcJtQzo9g07lp2ryi/Tj9m5fQe/2nWod9nVfErAnXFAxBbw0IUYxFi1c8cf
kBnfhIwLH/vqpbx+exG1cChiIy/CVLCSlW5Mw8xlIy0xL2Ox+im8lYbyiYh9hZkmmuu6Rn0GZXto
+TajIZr/Y1TLpiY3csDd1DukFpw2H58U9/BlOXmBaxuO7cvg90dkt/s5+8ZaW0NA6vFcf3Nq1QDy
YArMykZKddsQKAXeGdyjSDBC0mc3vWgFAM93OZuUvHhnSTAmEZXVDT8Krq6ot8sdBXkOYBu35Laz
Z8neJtHHQ0ZLhF22GGKWQuzavTUJIjg7IatxTIjb2sYy3Eik4zrCid0YMWBp+limr6hLvwoM9zhD
juqKyDxmBdk1piA6r82SrxMuGA8I3/RAmhFd/dn2BR8spG2ZHUT6knUeZKuNvhGNSvBw1ae8sbxK
5N9XrLzaKRsWwtHLaPpZncl1DxR9QJVTUnyjuFycf9TnnY85u7qL9Rf9O9+XhexIraRq+IQLBAJw
+U3VXqZin43Tdg6GTSDIqu73J5l9ruyZeQ1qLUQAuuY3mAmYTEBdXnKlomYwsI43gSkkxUHcdYAR
bTW4ACoRoydYbDTNn7R/eHAS8HuqSYACILQ2LQkHyt6pJW1bHk8aVchLuOX0OC9IN2J3m7qA1Qas
XZzHsI+Hl49kNYAkqrmG/MWuZh4JMl1MQAjta5+TrNm5tFFwPv8VufDPRbfPCaS2GLnmPhAv0bu+
GOovywyAljKL0RTeCwRN08/kBgm8GilRNsi27VWRSdab6OlC8QNATItz4+N/lWdhPfzZT2IzKbTK
o99NK5w0c2eQMnzItyBiJBr0T4Cdns7iuq0Cf+R9OAfRV9x7f4n4HPKDilF+ay0/wbk7TU4Va2Tn
CcIEqQB/QRD3ZOJ6te3yIv+yQ9/69TafM60ssqkGydGlZ+mCqlzD5/eek32CiOM1W72ObmYsYOhe
NtPzxKczEf8XqRyOc6oKs7Am7nM0IWHRVfrAnYP8G3xyQvW+WXf8vmNYej4ZhaIQlD5w8XOgiWfg
6sX1A+fVwBb5vplqyFDr+74EQ4jshOaaMAG81qg9rgPqQ7RNY04pkSQjbAQXjt3rlJogwwUMuWXZ
O4eqY/oSmQLV1FAjtTmYti7V8htbnSk+o3h5xS7fHtkaWrAtD161OUNfGzWevJEKNi37NmA/xXUs
NeQBHf0G0UpCgT2E+VwXsU4P1YYrCL4wjyhHZQHNSIgO6384bv6om5lgmaUyCEdTCLgl2fXiX8Eh
1xNkAt8wWwbsFFzB24kHZ/wJBKCs51LXGaLFZ0H+QC0WYp2jsnKc+U6lL0pR8gBHowE5DxIo5I1f
6YOZmUponzkpnwBMpnTLLs49El7uFibNVoCWFIVZ0wza24Nxvu3K8zK65SJt1wRzTH2bYcQIbgjR
MVXoxC6RbDejNqJZJODImdGhrxVZstyAPuzPu9EIw+yD430nSJCyCAI7wAZl6I4yuNXqcB5Eum+H
OGEFicwrQHn6RddCdSjMC/542sQhXvQ+jOaJilNwwybk9eh0+VxCJ/YHLdGWT9HSDGazFthXWDNK
5xTwMHR5nU+tEqM9+1S3Um7LV8kCXZr9MNHlynpp3gAlM7kYUvwSMjNwu9jva37qdD9UoVZS48Gq
H90GmtbO2JEBcayiJZUHr4X0qOvMU/CeWytgDw6UuWDGQp5RshbUY70K/YczrfZr4gG4r+JJemXJ
aTUNS/77eMbATf725/tD/ZLx2tmQ1N0lYwdKBMaZouhUFT5XYBg1wU2cp5ltIm9iGUQeqW7MNtoZ
LpKl1VXuEDUKHAMYT/mXccYabWRfv9WCFo/Cv3v7P631yzhY6p/JwhcDbknrGMt3zdcw+vIMthpA
s5HpmpNoBjrWdW2bYM0VL8mJ05pD43DIpnNxZkR4S7kxnpmSlXQGZgRkGuKSd/QgUiitfye51MRz
gjJY8iOKhK/b3cSEGt29l2lrjA4XK8biLRX/COrA0Fl2Ze8Iww3sN+UMFF1ER+aOpGwYEMgV3IHE
ypQZduTU46w+7CNN5NxWz77pZxK3T0nasRepe0C6KMxUQQoUpMha373Rfc4ovt6Ys2V6WGrGvLj4
RExyb/Zu0YTlM2tnBNxs6GaCmB2xcjpqhiznl1Ol1OldKbuL/Y4/4NSOUn2Btesczj3qFq0jJVPV
6RxIUcFLz3uESyIEBDp9ztkihWj7xwqzKSM4YQmtzwMzlD28S4CFdI1nTGxLEFvem7K8FmDz/ng0
N3Z3vLYgRAEL+FCkTMc1b+zSO164X56MG3qrlPUSprpuu/myOvd7QYlWyhNfhuPqjrcGhk6DrOvZ
nMvnlL8+oCSO4E8H93ThCcYb+8ngE9/tmC/tXi2ftc5cJt10C8kay7Be5ikdk2EnBLnnxgUekwmA
atpfx9m/R1V3cUvo9h/ANyWwZjXBfA9vb/yGoCwWKi+qjRnwKwiivRcnbueHZj0TdADsg+wEzJXb
1I1aLo0yBDacS2bb9hXS2x/sbfYyuxLZq+yXEslFGatICDhkHD1kqdZAD9xE968gvsb60x9KQv3i
eT7HttkNt3Bkq7dt3K4VphIlISsSIMgoeFs7gw70CTfqECKGq3LIIbWo9vaDzTzimIsFVQdNZOu8
tFVmTk2TqTXmsS1G8YO6sWTKQxX1UiD+pmc2vKbREa6pvP8scrHmd07ao35oJQ37VLgifC1oTEcY
/okrrhxYqoHg4vka0JFVlVtWGvarR//Ok45QRDmPxau8cDfDcJD7ZqcRMvKm4N30jJ6JWcrzg2VT
XBhOec3K+4ee55KpUlRZDmqdHsHqLlXPI8grRMe/XOWA4jPy4A9YQspf+HylkG0OU3pVSBaeUN4T
/8Ysmr2+PsD3MB0lihukdkz2sN5p8P21yLGR4KbEmeEi42cfQov+Z92XXEW4t1z7ygNWaqaf0TR8
muPoG00mZZ+dmaK3Ha1Ai3LL7Ma1yPegozxBhv2UIIny30Q45UTjh4OwY5J+I68Q1zrvwMCq5sPC
AtmLLACws/A6+Y+v7OkgJ38Cs5RBqMiroRyo+rxImZ9zgOTtivPV1VAa4GorXU/SHO0EMkqU7evc
3wD5c/Jf9V2Q4tgDv3y2t1mGo7x8BnLkFqF2qshWy12w/0sjc3C9kdzyOA1FoE3VC0SnSAf0OsR+
kwQh+EeKisTdEyeGZV4YW5AS/6GWocYfnxj31BChZiJ5uHgKy/VMxfjAwjWSNrsIJi2O+Zyl4ghb
wGuW0JaB0D5Gb4TbedRUEHw0wdK2w/2HhpBmjPkOBlrjsgF184yd443NTRFEW1bDNHKCjlpC60fK
IaRctkkX8vOc2TUhpRE2W3KplA8RXu9WDME6izEzxLfNylA5vPtueW/wXqv5oJLPNGF4dN3SEHkk
2l1SEGMySYtVvB47WSkcK0x8QvJ5DaH41V69o7Zr87CplykPU9X4h0b3BOIs87+kbMljarIYMG3a
jdko+P+AkYlbGSbhkzVea2dD8I0LjclveKqkygOJl+fvo1/qg05RCbhcZp+HCjixVFb4tj5/k5R4
7NpbK7gxmQ07lvsFoDSle0Ld2vGpd2WLT+cylAqFN1TwpGoU51v+JkNXPzfd4XyfnyWBn8r2nCxL
lkZlDyoYQkG/VUMpNAouneKg0Zu70fv3dr3s+RDN9YXXtJ9QPsFiNTY6eujS2vCchlLy8WBEzPcp
NmU7oIv92r8qcQIAbPRUc4KiEQl3urAmYIOrDlXe+EdDbfu+UW6EFHbvjoABz27zeadvWhT+iap1
zoJHiWHuuYw4GwfQIY+vni7iu90n0oIWYapItJjLdRIVVqJj9TGTY/87BT29CfIjbtDqBxx1K+R0
a9m5Nnnlo6CuO/BInCwBvUQP/LCpO6hx8vnQtLh/20+1iTgq3WjX0608HyWGlZlzh/4LAwgJEcPO
2Q5ynN+xsXytuWBQmiekzSM6L62m1aNRv1NGZb7TPQnq6ps4SsZJ/2PFktw453MU21RvNVoSMp3A
rlyynPLhf9Z8Oa3ka+IRED8edhdemUSwQGw/NJNMSwDSJVbv4Vd3wGStZOHDiAqVEcEgMDcCor2G
YG+Yv1FpWM2VDK3b2MCE30AgR0DK9C472SYCLDWIOPsKk5zgFhv7rYIGHdeIHPiE7/G9zB20DwJw
mCH3G3fESTA7QhLfkFjWAgS/c/dL8AnTeWpE57k7bo8Ie3O+Vcee8wU013B+WNTZh46Twe5Z3RBS
u8LKEz/sCuX87jmRoPfCobtjP6AGaYc1jhbTG0WeZj2xQ8Hv8QBHfcwSTYFNsT6+tCaulmjGuQPB
+3GiQ389O1NdgGpNEjEhvW+mYKxofI3jRPQUbz6JBplWpf8u7zRUau2kHmiy3xcvTeWW9T0ayb0Q
EOEY02XWp44PxoJSAMqoj5LNTfxbgzt+fs1x0oszKYB/FDAnNngnACfkKcHeaBq4e9brv8xy/hLu
ARZppw2MdawQa3TOor8Ufetu4OIxEg6+W8WaC1YLIUQCzWB3E+tfMoeoXMmo3YoIrmM+noqjGTYT
URL4/SZtDKSzzQaeflFWcxa1ZQH9BFfMtO117PNqkhf+ofmXDZwpJpyb41LNxOuv1jGdJUuRtQhE
DD6aw5Rjxms/6TFtb82u6ytOn2zBeKmFs7q+2Thimn7iM6hS1yy1+Ba2CNrrV0nCNSubfn+67372
dBCRUDmHVg5YL8nxekNNgh9PuZVJw8DslURrejI3MdVSCRK8w2YgatQ82KvgAoCKM2SdrLCRt7Dz
9v7wFCBEu/rnvzwEsAyt5e9pL0Ras7nmIfWhYHpLuUW1zT1Srtff1LT/22ckbZbUpLZEpRkXBqte
4CFRIfeCk/UJu8X8XDY7ApvcKe00C4tbG8uJkc10o2bnRE/ZFykoUToENrbini9sNy8Oh50pBvEs
2gEL3tuFUXRwF8jxZ3OsywPuaZ3gG8R5wjm8NzKYXrMu4KTZuYRZqRD07jnvoY1ThX7akPthqd7p
SFw3lPEpqhM77OK0W7jB7T1YXGDvOBXf87xHCs1b6j/ZN8ccp0bNwSRXQg8NU+Akrlcj5uOaJgcc
Uhk8cf+vHTDbeiMfAPzSPx/cQ7EW1Dtl4NkMHLcBF4EqjOTmJD8qG3YJWQcgHeEEc6SHdcJXLKdp
aHHwkF0/0hsraJhOLZ/TflVRRaI3hFQPxbqnMXAfl3zbymaRJuajOIkcWep9qXYC1JZjx/SSLSTx
L+BRlcUeQ5YX7Id7JVqxMW0BPD0D5mybLOndR7MbwjcJdH8Y9L0WcojeJ/unvmMbfbD9jFnM2TnC
8Ljf1ibeO93Qc8qsPHHydbkuLmHKLtiPMFuMP2JnlBBv/MSDa/nehWLP5KSNsg91+ok9/JBoie54
t2YjYZXR/4SK9+C3VuNKbYPbbuejFfOSBK1AeDFQ6TYiy+aTG2sxKJWaaAOMMb+J4CMz0PKa+M+r
KNfTPL9dL/ZoD79DJl2aDGKRy8EQoEmiMb+OYIUhyvMRu8wL0w+J146wF5ZJzNvWKTFcYn5uvep/
mYexriLaCo9L9j1zN9xdg6QYKdRTjHDHO8J9l+HFyRxoQi6kNCGjLNRlwYOZPKA28HdrlauNzXmZ
8F6pSDaxQH8HkGe/WI2JFjlCTi9+PdvaHvO+HJkDRJUpAnBaRCz/QIC3Xr5qUZi3C169kbaUttQy
DknOvGEqGbmWOU2hk7MWlznEd7dH1A4DDiy4mziN0axgbiuq11HS0TTHAwbxqwUS9SDitL5W+pUJ
1pCu/okIFf2jKfF0Wyo07u2OqfnDfT7G3qd/ZUBLQHhYbskKkgtaRmlAgLjEaJCa2E17b4VnRNjE
r0Gy6rWChojSyoNU1v/Pd35f7T+rO+75oDMBl3rrgHKNFyWbxMe3uuM9r2X45xrUn6izmTQIzGbt
IUSyy7FJg9Z57v+8OiYs5j6fJnuH1Lw5S4KRFw9tzgBk/b2W9jGj5cgj/jCXskQUi52V/Dn+aiFu
wcMRDjDIJHqS2+fJ2xJphwkHhI65mMx9HJd4XInZ908O+1Jfi0yzglpYvq0egeRX3yA2BJNbu7nK
fpVg4YTb9BfSp7cybnWCPkKOA1TxaQM9Jy8mRpoPAT0a9/f8JmsXB5X60+wJISlWqflippmv9E1V
gJ0wzbitPnjnM2VDol7L2oRzeKqoFM1OHEuZgWSLeIL1piEX1T+hO0TRH2rkj0TUDy7qGiQI9xuJ
V42OtWC7cpghXmy/bmmxTvJ+0BD8eQWqjRrujvuyWJrDm1ZXFeA7B0iSs9n7p1iTSalVc2LUlv8N
Yj6ZuXf58GsUgHroSQbq8Y+LpNE/Cn63T8WmBoRSUWXgRPoLjIhXHqwrJJpJbG0O8kuFA6SPX59G
WQ1ktelHvKeMrLBIsWJZwbiB94kP9W4+vTgiSeeYVuzwOV2M5VP6vNdXBvSS0s5J1EaPR+CUcBSw
QiokU58BCIom8OIuhNIeuhe0V9JbgTMw0cCH8wf0LJE5o1d/li3+iDNhVj/CC63QKdNwcPk0JWQK
ENKcdLhJZDI1kDyMar03gLCGe567TM6sLgkpwNMOdqE7K40ze7OooLtnB9yBtEEmNp+iT1zkvGKu
nZMg6bYCYc67nqMe14eeW8jqf1/646cJ52Myt3buU/Ph1GM+uLMCqAmgY2Cjqk2/Ieo828mpNWb6
uY6M6OxjL5Ukt5RiMIbJBpCde0TxpL6NG1Z+jQc6ViqO001BRbywvkPTzP0zJeCXq9Q6V7BPiVdf
GBRZjoNPz3SuOiNyvzGbi+8y/R2ONehF/OjVjvRjKI/+BahYddz4DDXaQUCjl6Q3ikX7TF1lwU8f
e/H8VpCNIV0MSnmz/d4MU/Oa+iuA8FXfYv1hPZ8K4ULmonXS6U/uT2FQphft5oBDqt4lJ+/ftLNU
+navh/fx5uqCKP312MnrHSQ2TjEm9ktG7IPlOLf0iLjHzshlFbcyfZw/aSS4bzQNlEwOaJaveG0e
99eoOSKHy8THSEZN3NOjgx7gvFtcDC2+ZbjATZItNX1I9keKdSxNjHWfC1pEfWF3aDzo+aGE+MTe
OPtrbAj/Bqi5hzZ3sTMxgi2rMjXtaqnmLPqwBkhhR1AZXh11mVHtMkjxhPJPXh9zPXBSvYNsHUha
8R+IMTA3p0HElp02LWfTNIr03+fi9xdOmIzqT3LIiDVpqbV4rTtXhf/D19ut2I3yXNp3/G8k+uvC
ys6+K5wwCC2+BkKM8niei2dtbMQwPX/pzyv3gMzR+olcGxgEEhhiEIh/GcaDo9sMN2Cy4cL7QvrF
IoPbQSRQscOdPbQ4DBo8oE/7rk4XvW01FrQTtScyvFJntt9sfnJgbmRt9c1Fv8k0OPZDsakRsPvi
jOIkZjkIu5HSwGZg9ie7C6MAOGceikhnCW1j9+uEzX2f2y7p8HypPt7ZejIb3JiP01Hrhq0Dtig8
2fyIhoCaetxELkpmeetMpUjtXHvQA9QY6pnOGOJxm3cN3g3MupK0a+aMktmMWtb8mHAv2VMGYJmc
PCFLAgzxg/RTA0pl7ucbZTEkqjm0ibGrzrvbpTIutyl+UgN77lkfw4iWoXL5Qf1PG88ZUWEzuixJ
gaeofQb53VPUAC8U5S5S0O1Totx7a+TwFJ10WCE7huUcPn8/YOEgILTmiHh/Oz0qVO+06suTBBe6
Z63YBgdt5mLg5SPPeUfXDVfh+Aiyl72x79hyMjpN2IsHmxIKxvzZbRXzAoE8atEWaH90sNUdR4Q7
Dzpf8xMKJVRYJIuJ1GxJ76EHPrLNVCb5eZKWlSHvCL1NybID9GVKrPBYxkEokOGQN42WosZCNMB4
hblGMgtGmaer3ffTlsJmoBfGlHaPidEYQ0nx88RAwkzx+NUS4FA//JWFD3tV798AapBwrEXfMXtK
1vhKWUdH7T6kaBz6mWPvSTzxMxLIeYZ38zSnx6KQXH5EeERieg39gaySDPypsTqGlZ7OUhfx1ah7
QuFMCcCi6ApPUup9DaqFfnZjZEE2o2lBy5FdXsTUEXBKIy2zMafN8GZrNEHGlrZWuxUUs6EqJrHG
2Zx6xDBNlSgts3aeGEAuD+Q1j6KaEfWUuwlq6ikp1hVAcKhtS/Aqui3jNbVKJ950cb9mAt5C3bgJ
vHwWKRmGx4Da/xCy3UXqvtKXdZwA43OSI2XE1knSwwI0p+YCkc2p7xYCtDndi3HkDIUaY5Fp4lew
ZFSqHsWtM/Q72IWGmUvt5XK/a2VHM0UVgYoZjmuSgNmlMBfc3L9CpEPClTuL9x9ZhkJvo0e8pYZ1
UeNcMdjh460KEmRkXB02Kfp0wmUK85xoNXBu7/9Du5UqA6DR8wovuwTen2GQRNymfwHnZyzLLgzB
VINwOBdvxJYXyAgQu3w3FB80bznjAeODrkDJuyLBMfAmCdfkMjfAzs4YfEfhPaCUk/qIlooddWY5
ul6ZMqO7bYL+tu2kmt/jKAQTqt8hT/k3vwF4qrX5Yae1qd5D6/pCoC2WaMaXi5wnOl4fax/fwWj/
08s+eqRyp+Rgbn7nXkrvyQfMql0T7ZYOkhpKl7dW9JmTmAQM7L6K4UEhYmKPTgTKIo7EQAobC7mL
nFmWgRDe/ez29sLlP+VTIWxyrcr768mJZAuEtenPs9e+G5uYcfLx/sD/dIdKBEqYNMUTBx+8tauL
feyzvT25n56qakPaMmA7TmvB3LVrN+nSxxZJSwinbphwr3hrevJm1DOpBtGAIv41WC1ldoo7fijR
IkQFAv/TyCAyhJ/FgPUuovWa2UxBt4BAVwRBQ+GXLZA7HGk9n1xQD7n9uKH7IBy2/IgVN02pPyie
b1/wyt1onBHGWC+WYHma0fZ+DpxfroiUenwIqq7G3PublNcYlUG7zDB+RXT01TZA2rzBaLJFQ7Fk
MNGULAxK5CeTzrkly1PPYc56MVcYUsBr1rFXuPJdnafdDNRlFOt0Yns4kNjCkp1yVCBLkraHgZKk
qGGdCF5ylB9QNwjClQYygVSFI6uNzQ60JXUHTGYimKTPIVSnu4KcNS7+UsGvfpqGgaPtdT99nxmJ
AHFb3SOkVdP9wpr6bogwdPDo/dQ+dNwkIgAX+xRDpxFvZbNtAzSSyOGGoXksboJjgCvhXZhaenf5
0uOcyniBD6W5CfRyvoeEjlsq84xO/KEQ2LuoIcvnfCwMlWQk3Xb96EFdK1akN3grOejJq+aS2Otg
wtCxDmtrvo5+vyMGrJnLNe4tgqGpuvqvSj5YfxO8oBVvkKKcnvUafpyExwQCO+ZYDEcYpCalW/7o
V7nr1QAQJnTQpKLvgrpd7hoGKbZgwg9WGq2sos5qBgkymeRpb9jGsYH6pU+3jMplr+zV1t/9OHXS
UKOqOdSoutnC4lG1uD9lM20VK4oqgbMhKWEEBR7458Ct0Ifc1lQ2LtbVE5nksHkto5LBbkScGqs+
EFX2KDBU2OXwLg7enW9Sp6fsmIZj8bmPz3GbGWvNFn84rKlzbcL2zGwj7umG3CxdjKasVRmot6lo
FvXxdlWhnFUFzdoNU5j3LQ6Ph+0KJSwHrHgN2Kn4Sx5XITFZrcWCLj/HsKqEvgv3XCl+Cyu7fQKQ
Q+8CVkN9adQbeIU0wc62uFL9G/dH0uQm5t598XFZpDKAmN+p5fY6ooqNHNe9T6WAMNO+nPd5VJDi
+ZVHOfnMI8tBU89aWjsTTIyjtCvN0AMMjxnsvVNE9suhWZIlfyBSv5I4MN12ecdvE5zsei3+wL1s
22jkVjh+sIHwlouK1+rcbQpMfEy+Lwdnkq12mEINFcefIXW1ASl0NvBcdNDS2sMm8QRxETlIHto5
MPrIfpn4q52whm/No54cWoj2IUTFrGcu0lib/k6HZdKzp0bMIStUSp7aaH1hmQ2yvSGOWKrvWBZz
2PWulgCWIbneF7VXxw2Cm6lQqtWAGpzelw+hD1H6ZQ5PXSjGSBYRdtvb3wEewbMMgebLQCJtXIiP
4cfoiaL8eToFh9rDlLPsTQBjx8U2KtTbyIjYvTxXqRhlxL0NtCiQUkdZEtQIPZ/NEFzTcxnZ8CAI
E+T94/6JsmKXT7T7tReuKeoZTJC1ZyUcQfJbUTGG7UVyUHXkyQlRpyrvLNE5RJp7kfXrcb+t27Vk
a7OTb5SxSD5Qcunde69WTu6LZp6I+LeqiijF+58UmyFZIcZF9bIje/7KsdD8H8tFwH22AquB3xXp
GCNGuLejZClEEzzT4+A/AX8/sIPZAiN38YQ5CQmGCY0S+G6YxnUoVanXqKg8lnDbKLjokUaf7qxT
VUo20Yy3lV/1Ki4bbUZEzEJKCyR9y38JfEJJyx5+BYwFTVNc1hLxuU6XtBjh3+qAHglL/i1zYhrX
JIEX+5zPNplwbFQMw7Q1ZEHYlRvtLGe/0jfTITVGXHosz34nzxEZyK92HLbOiptkrcEbs8//Z9nt
K/1MrqfqjaTedI6ssHUwix1Tug9GAmRMqljdxe8gA9Px++RvUWARHZU5u6Hp/v2GLdjMl+bjWUZl
zTVrrcfH+bimby7m3+80GxzeMeJCAYJLVGgPs0syLYWhGZpTrCZpxtLunT5kms0tGw2a61qFXzeW
85GwMAX1NYfDFvDYStfIR0FLF4mgr54XbZLPb9sFTtodnR/xAI8CUswGN++AG7u7l+d21c0EptPN
uWxQH77KtXnBJYnn9S+grJMYJzTt2rX0y3hJVWrb0J519AxcbmLOy9A6KwVolOxjav8vFf23khl2
65AvtQEJgq+UEkTzK88z7PESE2aUmx0VMydQlLftsK7t/5envn0h6cr6hQI0mG6v5agXlmxR4Jfk
ILi7utzGJfNjK3P1PijDSxVC1yKOcjHP5SZz3eEaI62IMBjICyvcLKUEVw5AC9yxVntv8bfCKxN7
YM+QWEKcDb0yG4KSdtQ/CoqyqlU6+eKszt2AMnMnaLjNfVAGogB3ygRrlgQOw1OpTBuumiACcvow
qop0RtB69UDyNsj4d9FMDLdkr/l5MYCRd8eceRqtcle99hfxOdWfwa6naO77kEl8BVifWD0RJMje
4XYTEqLJVE4hrx0yGoaPGeBCWbyrAnWdgBztK/FnU9XvtMNDRdaNapko4Qb0AWwKlZCdTjL+60w7
xQJzflqAlaAStbEMnCQOcwhOm2VIpPM4FMSVGkTpcq9EavZJEbJRqzPYy3wRFMbX1pjcDmWMrNq3
Jom7BjVm0BRxXaqwfz1IFi6iVjz1miAGmkiUJxhO5Ql4vB47OFMidoSPg8XJ2mkB0nhKQMpacLkx
fO8dLpH02gVAwbKKnWvtLuSXch855nSSP9s/YUhT5wFm0GlpDWf0qOsxRRdHYx2lHr1npYBb+pWT
HP4OykU9Mq/YXzAwAT/+1LSU3ZNm32mt+J+k9+US2GOYx5IS1lTVhzWA52oopoSaereAxCoqprpn
rZKXjRJVv1zQIWGqkiTItF/SDiFlgY/IG/gRuPvf4Xlb8DBAVE5MdESZBx0Q0CgI/nDKNL/usYk+
hypeoEa5Eo8DM7eo52sZ864NlFYuLc642y1xN5JY35uE7xxfEdNNUZl3U7ZNsZquXu61eHzokWmQ
IBdC92G18sLFB1UxQrOkTi2UHHD1iF3xKcXKgeV+UY22suz5MNDvyuDQhcdNb9+WCttellUNdy9U
S9kztpcVuDokTpW7FiK563fCKFHfeRj16uxh54rQxNW0lwDNiEICs/ZkqaOQEEZMOxU3GecoS8oe
QvLbbes0wYGRuk730BC+9iKL4aJkZ9IHeTaohI0TNgRPiX2wzNKKFTBcA3XlOs35jBn12gu1d9Zu
mNEl7BXfc3MrpQjGXu6Odps2LXmh69R7EukO9uJ8kVPx7zhw49uM6KLKiR1bUuhm1iQhhqPyYYHP
mC9pTZwJ09ni9Y1jU4f3NRM5bg/8hs5N94hL+z9iaOaIAlsQ/hfvJ0Nn7timxRYa4Za8DcSJZOlf
7tDukAZVJS2wZoLzXz1UxCMXiIUP1Bnu7YDixv9f0mSS6WBqShXhMPipBqLlJB8QKmgQzQX1F0rQ
TS2R8Nlug7xtG1Yji93w6IdzzqUCrt11F7Kjdb23Gf3DYj39qSwmIrUJWLXeWQo6WhF+WlFWucMd
T5oyIP8c3wU2oTaadClMVpj0LdyKyBJgsknuT+C2Fw3aKEvztxJXkpFEnhlMy9tlmBkQ+LqG5k1v
ieGEXe2SjWT5zM6HWLw+fckVb5HDMCQpZ09rcML3J8tYMujmsGgPvYdL+HvO80fgqkDS+iLc/92W
MjhVFQQsyQa9Sh9seChAwSaScRdyFFxMmXGAkhbLl81UdR14w7CNRGwVcH9kcw141uegInLokxBy
2QScOgQf5Z7af/Iq8PUzDNb6u82gKr8IonHipX4zrkNP35uYfD6WavTthb4BGk8x7k64PJ11Bf8Q
Bs+lYlR5GRSW+yKE1YyDPXvBzPvBBYH7GnsC871SBbLWjsjFb1ZuZT2Q510dcHDYGQvG6s8mViZW
MNqQ3ouDjvA621zNpvFg++UZUijAUKjm/jr7oFyWT2cygZt5bboSEzlg9cSDeVuRP+FzJ/XZVxkK
eOLIOAL64LrrvoKsN5rPHHRoZBoM1fd25F1RVUfp+m79W6HWhivjxmX6OR4L4YdeoR/isNhbTrXD
YXcqV3VQShUU0Ztb1tiOxBq6Jsofo+GymdERlQMQErGkKSRDGAcjEMhOR45fufOTmHxnYG4DUIJh
uBOrEu98exdbyz+S0kGOnT2q8Nlz+29PrcGq+yCKG1oToF/zR+f4phzmtJ1R1yx9UTuq5ddrn3/U
almrLN2l7jFiSp9qX/CEzVVETMEauqKZDb39IcE68zZEtPsxezBQs+zRsD+lYF3gFLcD8HgM715N
loJNkvE17fWfebQ1H5eo2peUVZloqCPDy4vAfUPnqgOUEEu5VR4rpGjPrGjnzoOmeQJufQAmO/TL
Jwv9ExbkH3DJ14kaayMci6EZsunejKfHJyx16h0D/ZhAqNSceK2ne4rCNyul8ViA+W7IZFdTAQCT
W9gYE0T2RVpX7o4LU82iCJLrpcnBTJpZUr9ojYtSArBRxaiqJ6vNMoa7Ytl5Mvx8MxM5D/dIWDaE
cpl9clx8nzyxT6jbgJkmBZSQV2Ip9ld89cj4cbXNJJ773ouh0KCbKXwgdL5/DttZGCX3To8wBBaQ
2xYaqfs+mj5Ach5ZNuG+fTDSvrMzCIggFs4fHysRPydB7qE/DU3fwZln3LgAa4oJL+stn8jVlWef
g0coIvV7rqCHJk03BSqhJoehjnQLs6wXaeR4oERFYYdTRPIoWAkJKP9Ay8mZqIk90d+9/tukytWJ
QeR44pd1uT3UyyBgdhVq+FUTtDSl1oiEHTEzQxcIZ2SddUXGUXr+JnUX3WU0MUlwsWQklYTKyVE1
FmHTDGD9EbNG9kW3jkAreJ5BaUrdDOGAf9VtiN6xPBly+dm6shVqYYeRgmheH9F+AOT2ln7bhPbK
twoNMe0Ty5W/GyCmmqvnb3zSqS+OGBYfVHdDiQfLUW+P7+0/lOKUNsu2ycBr95SWL04hADkSzL2Q
xwH3yH2nUSk2IW87+c/B60bfjDBeP+RJw2Q7BLn60SEIgj9jdLY7R4hrxyfggHsnl6xXPnANXOqm
6/AMLwGo6sNOMIiZlfcMlOBHvGSvYYESuJ6zfYECMxUvu5KtZwmfEeyaYw0ltdQH8IvUqB44Eoc0
fBqq60hMVx5Ct/MtcctHEjulMgs4M8B0IhGXNtGL+6Ytsr4wa/0abqInfvHAdol5g7ogh4k46NC9
NcMQAQ0eiaXx+uYaB97tEM6KoiGS/xtLRX2V/aq+zcEY366H2rfxSkmi0Yo40ROTLNpjAlKXWk/L
9g5QOMaINCIIx3V8qB/3uRjb2z1VAP0F84R0VEJF5xjRHXgeuGxx2EFsOjSvLZfEYCqDSfKC7hDA
z+trj0x8poawayAjGY9YAQ3aGN9rQM0ECWnw4CXLze16gdP3rEPN5HTo7dO6RUcBiwitJ0WnyNgu
3PAb1spqDeEsXumSZhq9xRPz2js0k6OvuUYV35MR8FXY9qWTzGl8dCchezp4jTu4aguJkkl2lo/R
uPfHX3eu4ODLFcOsxhsspb470kX8Tl2hKE8zMlJwLdefu5t/36i0yy5oXCpcRr/s76HTc10kac8E
lIpdeydNbgrQZQeekFWc3GTBAjKHVC+5cpn1ByEIWjAy9kzFePWJ034MwqdXUXS1vY57OoKi6lIT
ZBpyYTENlTvKHB4mg6B8JR5pR9ezjYVNmYfWqX+42/Q13wBmMZudYGD8Egwm1CC/47Rj05CwwxD3
VrIqLTHg0Sz4GbnC4az86cpvZPQlspJupAIs5uwva7s8uhZ/YGx6quZMfCK2TBp8xi1pK4qxfTtk
yyvT6sZKtlrVu0UveJqAPicoIKh96x+azu4rHQ0ipXUrovQ8OppnEyuvqHumiQQVdJlxiuLB44Ij
P/hL4XYHKmii+HpgDXewzNpW8J7lNUI3IvD8HjH8K01ZPX2+jSp6BQ9rCgZSIaAQBdh+RoRFPDiF
n1dXyXMlHyhFYixEr2eU0F2XTZFHjK3SjT7i5bDF0aJMkTcRGBRv+5/5n9XMvu1r9n8Y9Hn7JImo
VGM+izbA6nqtKQW56uZt9IY1v444q0exoxF6DAfXQOK9TArzpNqdZknhzflyCkMr0JQCvqA0Yvjw
bmixSDeXfad5iNleoRp8eB7PI1wgp4q4kVHrZbDPDj+UvpIHia424RXk/UYKabdtXz1nDNqYz2hn
1GT3NDddEhY3OxAk0pv1sQFxmHeceDMKRtTBHO6LSX5LZ4ZX3jip419SckyTN2hkESdAxm8TO4mY
p2nul5a9qsMd35iWFNYkgO4JckN/OvNNY7gf/K/opamEHW1/dHPyoympZ/EMLkX1T+H2fIZGkFge
3Pi8EsbxIggiDlLBbaF9h8SVdLt2CBlwOqZncUBim91rp2oV5sKRshCAihb9U0mv4wQoqw3oA1a2
Nsjl0sT/RSJZ7tUju/oTsaq1ABj6yQmqn+E+ni6YNBms6E1MTe0G/Ys//PNa6rofv6/yCl/5aQgG
YqjL5UfkjYgiCY+CB1khcjgfOyFsrJQQM28lxfQMzoHFzn50dPmDZ8beBSsaRpnFsckdh4VWJAcS
A86g8DzQALfOp/YS3fF3TE8u7QdyH+Bx4deVMXA/R5/j9OwdIvCsaxA8/OtpYQLEtT4uVD6MRUVK
yqZx6x6ARWzr4E1IS3kMDsz0rsQeAMWgAHxjSxdCGsX4Mn2xlmBgjlWh00OSe/JSj9ViHETAkii5
DnH20xUlFv/sJrjavHHf9SpjNRwjOcTGKd9iXBVrKS9N6QoLaBplvwiwONsCuFOKWhZrxkL8IGyQ
vmBgpMEwSS3J1I37s6ucjdC0lf5a+meGTF7IKt+MfsBEN8QDMLPX4rCS8lgHzGhJaB37S2u/TmX2
IyfIPC0as+FQJhV5mw+QcvMKv4vGOZltx0lEcgbzU37Hw5FDMqhAE5z6BkzsAkUzG4RgPLF0HhT5
aZUBU3LQ0Y+98rBfGkzE4zGHYRbtaXxUbnYEbDBHMs66cpMJFqPGdT1OlykO6WL5Z64gzJwfG+XS
8WF3IPC1K00MczeHkuOQfwk6mIgLHsG5SVH7q4jlbRR1lxUrMlWidIQnjgDiB/gbO59fNYulIRB/
ihm1giETNOONd41YksBkpWxmYFS0wVmOiVdzMY2HibncauDltmzNs557KEMqAb89fmDwikDH0Q1A
KtOKYU5UScuzfFhbm21lxheycFfv4mTnACDQxBnhYErDAlYRwHqOFMyETiDr50iTrLeOEIdNoMI3
WBFFSiqOSN8GmztS3ljaWESP7G54nUjoLIxrHPKjwEVxoYgS1525Smnl7zZE/B802P4fb6lEDYdo
dZJV0GvauHswHJQWRPnb16JJfwOoDSOazy860YgUMg4+wK4/grCNIqLMpZoCkCBJildb/J6SHpg5
jRCNbUUgERCtZpyU4BMjvu6b9Ozw8mrDhnv6bfKBE7+dpwANuX39+EuYGNM4ptSwYeG9loreNEui
iApuGY+UEWrsNnLdEGoIH9BwTh+i3SsMJy78qDjtTYdtfL2PMs2RBzVV97VluaikEWGDfMTRhJ8/
8aVyPTtLGS6fuYGpUUX1Z9qolP+h7QDmDi2Mj/XYt6fk4r+8koDEc9+jBg7WQpsh2JkJpKGNPNVe
rGddTald5qdelz3LbkyxPKjLPOoau58oC0g9s9zieqa4bg+8VlLSw0Zh2jNxt9O1GdXLvFwATm/i
I3mXQ1lYpnoYOkPdZYSfOfEgpxzPeF4lIrrA1xDzWMIMWaz7Mg3ZTB2xKHfF1c0P3+fW5/QCNQVA
TqAOR4OpxBX0nHLFIsjrCYqDQQQkO5X5azGLMR1PdvBUKakScOD2mIrGrVEaiy2XicdhZx2dJ8Gs
/syS0XfXUUDlXgmQ1pCrNV2dVnFfXGeWLG9b4P1LLbPJJekSJ02XJ2xpxkJzv+2aUVeeMHh0Yf7v
bYEsEnl7XLnUgWM/+LEbNMUxDqlpM5MmMEUYvUwglsCSeKur7su6+KvHrN/3QXkYEvX1Za4/9Gh/
YbHAd/viktPj9JQXUzsNOV+02udCcZFpk7lVHfRGCg4LM9LfmjqOJrOPcExqLus3TF62lgtedWQO
sA+vF812c3CDzy/ZgOYCEZicMe2Y9dSrKGzoYSQepoMhFcHz/Ny0C3A3LdY2upYKBA6sIWrWeDpO
xQK/FkVURsmCyKWLV7jVS+6POp6wWviknbauaL4KJLunV3T4Ge3vA/pXeSLGPJMrWVYganOhuv1Z
va0gnnlRsCNWBTVBs8PO8lU4WE1hfyMSRyb3wTyXxMojD/4kJLAPHOpOnD4pnFbz+laOKopOR9fb
fo0tgjwgkeVViJ0Qedsr2JkuakddQSyANDzENbJh/fnwZOnc7H8hphQz3nr5stH8fYi+Gj9apAuA
W48DbXtujtOnyM0FgH1qNGHEOaHHS1fjv9BgS2TY3DhzMPtbsSvoBIuiVEYHzN7+riKC9cHCjd9/
p/vkizFiLKJpjpSYUakIawxZClBVgHlLJAqNOcQYlfyty9x/pNjHd/uGZaI+wNZQCvRnCEi6BxKE
H+npqasvWVcyRJxP7+B9nB7Hhm6wvA68b7+qw8Vu6YqJchBxT7dt2l31PnYtgSlKPRjjy5AcDlaL
WiYYG3LgGJ1SlDksQyY5KwNlMtSMeZA86Fcmdh2KVJG2Gthx/782PacmcCyrqtTtvsQlT0+49Cau
41HbeHCpcA4JplRM3cNrdk8SEUXmcyZJoXTR/aK37eCbmDURyCVVHqaN1lIDYTgHiD8BAoPscJx5
ur4sfNbmott9iApzQukXJz597wrp9G+jdrkXAHpfI8UH13toLMy6hHT9qDpux9ZnMaHFmEgYlV5j
3TuvhQC8yaGbi777HrgsMDV0gOAK74dwsPwxi5wKmdDvV73aTi3NF1QITlzrJkShKHaQj3k6r6cN
g9JYOX5Qsw/VSE/UsEmBEYyrKgDnXsdm8Dt6vDIri0zxHOhGLf/qME7R5UjlNiRiC7VgT4NsMoEU
4A8x28O+E+uz02w4nEcfhu0Gx9bZm7MUdp5Ncb33Ek0zpe/4d1MVA0GS1qP60AJEdudAaK4qjBMM
0rNaiM4J+gTzi/P+XKVLfJZ+9dmhhFwBKcxoyBhOrfV8N011gM8V5JNkXOSfEL65HepQZfxuL/J4
p0j4A6uwG7158Zs7oFnPAiCYDqQnuuHOKbOm9GOqk7ahljzrCx5Nl55CbU1K3uzUwGidCoAQd/Pb
qB8+gSm1h0EuK1OFL3CrRSh7NDKRdcSKkOAgT2spjkq0gsNlWdl8rNVrryktUs8Hq5Y8Z+jCB2sm
5deEbw60mHR0eeY+r/RWNTT419qBxpQWPwdkPPlmUARj/EBNS1GYpq/pujZF6tB763BQFhr0Vm6Z
hbAIZuFSZa/6aTU7QDKmIzCEj8hh3Jq0Wv2C7cCx3W/LbX8rbuonT/C2O5/D9HJREcK5i8QBmeg3
swjkHsWizCvltNbmSFsJqm6/RpD509VUHP2rbh2spj+zapJGBsO9zdDouk/zbk6HZj7gRO5cO31b
ox/e3h2ABSQIT4B2X9H/pspZGJIiZdT08mE/8j/WDSTWJWrzNn6CBC4BOAkXcK1NGGSRQLxtcA64
cBwNsIKrnT/JC/HkkIkmKnPz7TZj4T356NLBbByDE36xXUUx5vW+dq25zAicPSbMT2BQ3xIxoauW
gAlkV5Ye4nMjl1feNodoqX1iVeNEVFiTAe1sd5kcpbL9kRswCZkk2FM0GMfgkGiK+f7vbYidHqO4
iHRHXdbCsKhWHFHq/IiTIOjyCBO0IpSXoDug4FY+Dcg0Y5BfrrcfqG2zA6N0ZELqvpFvoLBD/sGq
Rz5BfCB/4GfK/l0+vdNuK251MN5FmsQW/xNAY6Jt6m4JCGR40fok2NWdhnSnMm1Vd8zR5ysrbfU4
8GXeeJUV2jjnTu7pZ6qjCr3HOVleTIiGf89SG/y3RUiIJg9Aa09XuYN1dOWM8KloCdwUJFZgROh4
iRIMaLtEV+wx6yyNtGEtPHMbTUZrr4QhZ6u6q91kN6ENaURyFquhJrR4gGVyP9bx9l5MrRb2nhlY
DD1cbw6LUfe/u8gEwpQzJP1p3vpNtoy4Hk6NDcxlSggdtoVWXhyqcVAK8Cz6PmLfGD/nSCRW1un6
aSx72uks2GOFZQ14M4k1hnd4C7YyfSYBoAATfS+caXYJil6qQ/R2ebBSI2c21YZNb3uWZP5B/QHF
5Eqx9Y4zwyx6rR9lYyTO4uKTLwtmyix7zxwrEHAZqEQk+cRFveBJ1FCdekFfK3QaIfH5YREdYQeP
JgvWOvIOfT0YbO+UJbQp/yJ/yE+whwYyhU2T/YJewQ7nMi9KTfPkIqbnazzvFiNKsaSffJfBYOmF
zEw/XPyxARuK/8Lm2i8yR5Sb8qaV8CnMUY6PynMbZefQVLr9yBDn36v0kSQJoHUjZEBjZYyZ8PTm
v6G+GsV42KF4jpk10YWDDqi9JRsxrIiM01hfsNN/ctg7GfVIL+CkF7Gv3wtEpU98pDma4330zbsp
3bwFWi004uDiaXZFtiHdxhLMIH+72JQCN3ZozjzPTOGjh0WTTT/qmJFzHr6+vmGvIVDRFqFGRL18
k8wkO2nQ/WuKblK5uYvFLp3zJTlQw/P/pbTdwQahl0l//B5KDLbbZOsX/6XyN/ltziEKmsWxXspa
Wage4l2yWiqbF6nagxN7Lwaqd7EPwiZMrV1L/fojRDtmh+W8a0vUcv9igiWNbsfr1ITNLdF9K6XN
zNgqCp0/FlJLurWrHK99vVb3Li36RswsYYB8vgaAV28+3GVVUENBYJXWsVWz6jCo2uN1fd6hiSdA
YVQe5ccUD58F08L/T3t5tQRv8F44WejEV7gtVQDQ0utAZw8mvs9XdWVROrzMbrE+z4CXnfs2918+
lRAVEm8UYnf1bPZUHKqNlcx8M6582sQbK2mMQmbFaW4m1W2nxv8gvrEOLMTUNwjRaI6ecKPnzv7l
/3ezc2bQ/Qx7eqjPhbU7YZd5tFJjg/56fM/8BPimRkVAKpja3iSElUtOt1QxqikV1ctD/9CUEiKR
xK8gxcE/YiepOUyTj/D8ZxPVlY5y/XAgLNJ4gNuLTeQXMCI+feE7DLdlrwl36W0t/yAPvM9VY2Ll
Sf3hv7EAdxkisoYIOtUVmel24m1JUkR7QRGpZXUcGZKX4TZD+oY94ApgqGTSefDKIsetXl4QWo+q
NiM0vysmGVxmtvHRofywyjRAuSxEgHDa2Vs7fxfB0oZZa561ZNoOWbiJt0+FCPgYbXQm8gGPpuYt
wUT5hKb/69YqArKc3FulStLbp2zmlZNGWk8kKBNmHIenPdG2NKc3x6rVg3VjekKkUfk6aBJS2eQJ
cIyneoFAzZd5xaIHOHThCgduMsX0u3c5aW42u59N5znOUexYbfps6rOGNmE/MEqRJ7vWuGWULRja
AS9A8RQGcX5hypceqrMwXXD7gQFHuz9/1gXhsBJ1MVGIppmOXgYtJvOoJ8X763/E+EBlDR/f/n5X
mMc98hcYFlOLUJQ+C7IDkxRzoLBlzypX0+l65uqaSPqpaMC0rPOrAMj/Aj/SD0Fp3JIvreF6kzLF
9ESNoSCJ20FDoHBG5VSvCnA24TByTgU8+13eJgdkBmUJjwHZ/EvWTZ4y1svwHyr8acmrN3Mk8zSv
j0Xl8/cQzQCxFusy6SAdXMDI7P76P0K85P0PlhUWtkU+ae5+Kr9mZjGxzRZDDOjTb3xY/TYB/3u5
CqC3udUjLQZjOIzWXBZM7yzb8VhPqI+Wp/8oC72V/Hdix0ohFhgecDctSa5gT686oGjmNTrImH8H
pf5aNl6uhiZA5n+C5oiQRA96gI//6TwTi/Y0WJq8PbfMstQbDvUB3LOAW3wZ/Ll6M6nAVTB5T/le
lNLBm7wDgvh8TTvdyLdPaTOyG7lRzzC1E2PY9HfgOPLn7eQQv+ghFxeRo3XTvfkDF5CHniHAV4CL
/aXKZQ40WyUqlqdjyZGd+TcwiNo+7nMDLgyf8UdN0cmSnKcD3KQRiks1aidGozvbIyZWw1sYy7D2
c298ek1/W/pTbUyGNx3Qi775psHempjIAALSx+9kbhuLSodGrQXIggmjOtKGNStrTDkGFX5ryoHT
nOtHJVThGrZa6/hleH5ODZgRwvLt8rk572sCuucdKCSjXRe9RyNwfP7du/gPGLS+/FSzNvufywOu
gkz8E5CaxxekDTqzHqEF0H+GorVLorHl1Q2ko7OzfxKB/jV142K4IYsyk4jepGb9Ghh88i+kXJb2
1JucetTql+UH94rTnywIv9ugaidvUapnku/vMCkTbMeHb1zz2Undx8IYm8OrNOrRVCSe/eDW2h4g
G32tcvGqWCZIVqZ/3Zf9jAYTkprT2bNm74zD0WXziH9Y1MQej0nVyfaRlRMjF2LtSj9yzXcWYPVG
6tbL8xJrrOdI6fpjzPHbNX5WAQGdfIiPCpx0t2j8RvxefTamg67rMCbY9RZovIhVriIOIW189Wj6
lGp5u5rURJr6HdXHQOAMiErjsQ5ckfYsaopp40B8pcyzm3D6UScJRjTd9gB/wot3HbqvVsW4Esxg
wqDsSUJGkUpxY9XJoxzE3+zJaCRM83CgqBLc2oL074p/FRuXi7Oi5A9pRCtIM9Z3IBlJdXhvQn/b
yDBpVytmgAwavCygkR+OCkx4a53H8Ay6XWFskoXrimZgk324OwjrLhsYO4RBhSfdlgiMDWgOiuMG
cZo/+nyg8mC+UryAKi/kyHbKipl3AxG6cZDCfqIk89jITvZ6bk6ERkAzr9qkkGqIiMHe0q64L1IO
vkIhzmytkhV9M5XO3fKqZVCw03I7RdawdwK61gFFj1VXmrWeFFqeZ9kKp6gZuaiUsqt3i+9LynhR
eujNQhMsWik4hLtOgI5MiOJEMZJNTL7oaD0nhsBPr55xaz7xjo0LOhkL78P+jA9Aooe5saMsw9Do
/bii6X8bW3ULZ+We+2+VoGq8ui0FN7fevrrE9Ds0/x8nJ55zZoaZorOpymf8xqvvYbkCSGVePne0
0H/PsVixvsgQIL0dQWWPobJfuwIWajPPmt/mYZ6SIAzPMxHLN8UPPVO2MuELbzCUTDoBlRIP9W4X
pP7J7W+Zwzdm/U42rfEuJ+ejQj5kH1/kUUgEqtGGk3WghlREpg8LmlDUWY5zcPXQSr83JC/0PlzT
w6nGwKv/dHLUtSIUMsji2dFddO/FCvRkGS/Pjt7y0rSyJ5p+WpmyJMcw2snNrT3bFrZV98D5P1jF
U1HIRIGMBpNj1Y0HW6vAFupGBc2X7kIPvSCILj4OdqCmGJeIE50EKLTdQVCP5UqvYTDh1Td7W5JY
TW6FbK4evKRgJgfnickP0lWFgt/4LHmekufuZ4Y8IHPcPwGcVDPR048jNZaJPo43ydwSiKC9ccKg
s3wGyxVOU6czqZ/1Nw0oYTQacnxJjMoprh7Pq8YOGUzaFQZJuju9o2dLg6tPACM6xr9j7Nq5uCN2
hdxqm5ZpBvhMaNGNwKnS/5DG38LJPRNdbdAGx/PnhfbjxvpruqiXUeGWdxzk1mBMKcInI5BzW9Rs
m6t9kOrHrsEBwu1YynNIyMn2YSC+OERrEwiGnZ60SGRx/TaL6wTHBYqSI+Cqy6lNxE2WBwIa7uLK
VCaZDeE9+Q2NzScbcrw2bx33QOGdywcqES3tU7+VzCJ5+yBHFlMVQ6xEBFX7q3QtYQwFJiPuJaOD
M5cMnfDHlGJNDcyBZJSkqAn3K0szmFsSwN+OdiEce4hwp1022ZHy59zxCBSp35EWEflqmfhxR0d1
33fW9maweYir4p9b/+HDsiqCugM3Ij6jHXHM2YYdVUBhuH4sZCatBsbsc0Z9dc5F7W+CqS+Up1CU
j1kNiFu8qGqCcrmK9VgXqKtImid6H5DjpRdJb80gypahhf8Et6fItUKcVF+SZjecDyERll1QUHT9
/gy+YiHc3GgjyqZQLsbyGQ5R3jQGutk8I8MpDUNgV9xdmHhZGIwYFSqEgHFzme5beYgwjVGkcdXP
YWTuIpYBtC0c3r18wAWpbdCoAS0UlzjhaRQIdjG3ltaZocDuXsmmHRLMR1poHdsKDgn8mdH5bAWA
f8B3mQuSyDjnAz5f9IDLmKPcfPW0rj9ei/bYBX5LI4u3JzsoFVieLIGFoTQroGdJ+vO0Q7+IUc9n
Onga2GfaKStCz/LdnmXszmYRtJXoPVO31hYSMaYdJN59WJvLpxBGVBS1oe/GsLenAf99hptQburY
itlPvVpncijaMX3J3aDbqaEJZ8+ujEBIFo9xhkA/OfmhOWe1W2M9gE+OxX03jk8D9Qd+yEtg+ygU
APIdVsoc5/oRwmubVfbzyNaKVX8XgSHPlOpCjSyq8bAhv/1UH4GH7V0jvOojN96jdP/yCcR1u9Bs
ESWAoQDOmYAl4xYIR7NgecZWzGowQp2dZsfgHQ6MvFJLX11zGVfBq+9DNByTT2MDlUsmtCdJ5KyX
S7g7xYUjOqbxDp27MBgh6tkd3v8MVGRylnF0oYqjmlRw5uh8thN81oMn3WqcTXrXbL32KgZYNNQv
PZ54dMEKxfY4q43mzg+GhqoMhaCbyLnr+6ITzIelm2HjqugMQYz60pKTZdqbOoSIwOzyKx/T/WWN
ysyTW4w3NfipZvDheGazuqH/tuMQHw0SF5VSaUTLyVec9g8B+SZJNOP3bTc7r/3WVca/bY5SwIjl
7wcYHpStEbIM+BBIuO2rZ9ivtFJZNW3YVkQU9oigNMiufgpUYTRvuEzjv2pyBK7PS8kntoo9GTm4
g/UU8kUYRvM8B2y/PeoRx+e4cvF4zqjE4pPmW84GLr/UCRKDYN9LgDyFls+VINkFSFiIWlN6iwkz
6GwL2y7D8WsExJzAo1PLIBAyJYQ48mnGz7nwEH5teXoKowZeNsvwtviI6W1v/s+KBNOQGxe04kOA
ds/o27wcDctWlPIOHFX08xwnM1EIOd0XNjmLhnCv57TjqOU4FnwIng0sqLIoIat+pKY59SVU2GMy
3ZIUB5uy71wiUWO8yCIqRwS/dvJ9jQwy8IS7+iPZluWaq7hjBQiTukHOGtnuXsFVMauBVW0Wtvci
QJlGzOfVO+G3reayLWhvBAiz0qDAAChwmUPXgfGxK6J+NuxDgjTlP5IkQ4xfhqItTr77Ysxg4XuO
rc07BpTIfpta6lvWkZtB7HUI8Ob3QTs2sNOGP5gU/i1DHQHjAaAGoMmPtur3+nsfnDQdDTl44JYd
vSygpxkUT7tvoeSzDCril/z2c8tXa0lOfpbcbcp1lvjPvMqzqSqqDrVWK0WX3NEW6gT1RTj8uz6S
jkbMzSV/IbwBEn61EevCO1Z1xV0mPQEnkVXQ20s0sqmZbSfPPf6Z9tUs+gJ6OAomUGTzJ7I5da8p
u0UiMk5c/r19LuCi5IeU85a+B2zFjKK4yfUKAVAD920YJ1R6tp49Tzn84iA/CMqc5MCjchMSNcqz
uyJLenMEBQrZ01mV2Y/fyOdsa3Cpk+B5fSYP4VbgtYCant8UOj5Dy4YPBeMCJJc9+MuySAYqF8fe
IqDC0haKoAaRXbleVSEvC+I1CvcUddK2DAFd7ANUBkyGvg8ICCPRak7jfsdSbt2o372Eu7IwDqWj
Xf4Kqy69MCXFNmWn5735IoXFJ+7Jm48Fjsg8jjlEVuE0ierGg349WaaAo1a5hCM4kkXw1Nh8rYg1
lIxMywCL+1xSL7CmXpxufWhXQ1i+YLIxI2WBWVOeN5n4ku/CGkjZg6iPe7YDpyv7jZtUnHh2lax1
R/e1GSdchcrpxL4/zyu8RlcqJSGrdRNJiXfDRkCyyv9dlTw3h9CzJ8JzjjWGaVBrDVnmJfdNlqBG
WtcJRnt9TGjezzSbk47cMdksWFXtQ4hzSDYjra1PLhoPSjyznp0tvOKUMc0aM9KW4eucV62UJ+34
mfXioIUBobi7QJq7GphKpkJ6itK58f1tbebPX8CuPRcgwt0q0uQjrOXYtpbWt1i8ZkWsq+POedeP
3E33XFOfdB9sMMJnN9YpGRyhMobgQqf4xCHFI89F324m8dqmPhselTd/Swfk0luBjbzjWT2jp6+f
fxdYTaOUK+ImLTBLvoNNb5hJYFjv+5Ed0XDqWSExt5CW01I+8N86vX+36k7dFzsSoOGk4Rq/vXP0
xlY+cOviIi7UAO2qm8dlQh0K2k9TWKpnvfsaFaFVjf6MLDMyDNMtYp6j6SVWHd6IHQpTHqwkRGku
5HJjeLJtxi9V8BPm0BpzciIy5Z4z24pk8AOR5z15SxHHcXMawVlPIiQ4XYI7fgPhf/INIz8wBpac
mnWN1zPrz/UYK7QNciwWXIFjYoAat6bd3AQp6oKIOHjkOBytep4mFwGYUVExaUYb7WHTmzPqiUSq
9VRXFp3dI2exj//X9L2Fmth8wV/V9voT284tlngphv7gleFoxE6qeiZjDhNeOANYB3xCAotQkJXz
fD6y+COPaScD2B7Fm93zoZ2PHqGNGBUsVZyKv386v7aX7J796sZqhdhItKMOGD5KOnMT8mO62nPA
mYwW5o27As3cKOvEku8qUzWeaaJkeso/NZUfneVB3A6EygPCVwfN2GmN+gVe9hw+TcUg7OX8n2UJ
zr9XGwrrn8oXOYaWyYajAoU48KPlFD1vkJmyDw8u6BmopnZKlxrvio4Pwmg9cqiQDIrYth6qpeDE
4DzvbjTsIpTsRgn6bA6YV6rVciJJncSTcq05fG+aIHV1xmHOliQZq4srgexLeQP9QikPRebWs6a/
Y37GCEA3I0k/TqMhbKvfMf9rlYX4S3GKxehGu/PuWtHIMRQ9Jj2/HToYXRAzJdi+RH0XiGtExidk
UFzU4n+4lpBTKjw4SP3o7m8fx36/bdyvqQutFY5AsXkl9UwjHpu2BKt9I2hdwVbbL5gSFRPCHDKz
bXvYLsjF6LexzRdML65r5PmhCO4Wl7/tQdbpviksVvjHHRPMHQF6oA+jpjFmdCYN532L8gpZGSy/
mQ+MEliRzVs5acV+Lfq3kRXWDMIvGoFexCMT94BZVqDTSig/yt5pJzDJjwJqweRJ/1ofQDHY95ub
uMQ2eSBhLxND79WXnFN0oweBBXm8CSikM6RXxmPILZ1TF1R3tInxwVGRh0DSxo8aLiDu4Aa0Kwrv
Tr3/fgeFYaeLVODRy9HF4/mCbCVzyPOqhzQozOCpVNgindGZ/AXEJqGiNl7QVsKZLTrt9mYt+pU2
J9iP2V769DErLL1X6traSn0PZohzLm7U//Ii23qUtcrHFh8iDR9itamZADhyCbBu2/HB8v1358Fz
Tc3oYbCTVGtCU12DvKH/s7fN073SpJVpoi2m/jGflItepgmZhIPwt5Gfa61dTEpbuu3azKI62DI4
1ahBlIc5COv8z+BZLvzIt1ybxT/mXfWkE9VnNwaOhQpgDL+j8hcJb9Gb614GVz1b5r2PqiUH0A4k
M8dbMHNQ2qbFsU7TJgROg2qgs3cm3ovmMmeHQmEqFpOczA2wwJD0Zz5qNmy8kfy1AcC8sKNmLD6n
9EscIto/vTcAw1CsO1lO6yfM9M8+fgk5Ga6cAQSbfUXNdEywtAPhY3ZOhKHlxnraPXXsdnsIS7NX
BO+78+TmGjjHfzKWuWAYuPDNFyHyt5BtNranPHoCjjTsp8oe6wUNYZdRh+BiWdbUrTqdNIulcfEP
xBqFoKpXcbVJfqmpFJW7FxVS8fVhPf5x0titp1/KbAyun7JXJejKi1gqmueDoHQuNgnXzcC9sdGY
VHE9VKE8yW51navf049aeHPl+CRAlBU9qComSt4KJHPUu+AZePsBZNnp2mjzKVfVhj8G2phDV5Hy
wvNgGnuocytJXilYBuXxrPy78nFfwhlOFsHa1xI7B91Yr2fcbByxVVWaDUbhzw8PZuOMwnI+Coq1
Z9Fut0d0fPsuSau13+IlIl469TmGvMNEtskRwagPsivNgWG62QHUH6qGkKndmjQq3hyQlu53ird6
GsoE3jkrk7FR+B3ugaezmfdMsmA3TTb/QvLKle+DerTkrjoF2frYYHs8h3dgWp6l94HlR3eMv/Im
ShnvsMa5iuccM6o/9Xq6SCpXQWk/7nl9qUlHMDc2cLjKU31j4rzzEwP0JghSeyvhAJfOS0mTjOzg
GSrt040tkY7Hh20LMD7VQi9vfMV2RRrXQRQ2ho3A8NM75/jIT9m/vi1sNWVCMh1t2+8T+QfERByT
hkiDpgVmegPzrUlsmfxqCesqZxGGvwuRyuyPllIbwP2Uzy9Cr9LjosmuQASZvkj579b0kQOvu+ZM
fQGqjK78T/3wn+3tVg4FR6otLYJsK4s5HgLh8u5riKBhT7yztn02+Z4hGX1B21Y9JvJspIQEGpVA
OiHYUx/pegofEuWKUnEaZgpm0qUkoFrvCskdVCyK5vqDzqm928QENc0KzZoWhYZHxgCozgPVHxEi
FOBzmLaKBQul7e2Iw64rXlrAyalJGSxNmxg1qWX31AP74Ggf0zypkVNDZ3HFBjsYXiFfucDdnDup
JJhtmqkSErIF993v09y8miiFsPjfwRtqf2UvxaofMVkdLr0a4htmqKF/+XW1Q1Kf4LovPlhUaAWd
mfOUl2gRQ5ZbtSurDJN/wCTN1i0cim6y+Bivyr2aMH4xMDVGT7w/IRUJxC5znk4Lvw555NrEkCPW
S69gjzGgwhQm+ju8+IqrN30RuDByNCMxk320pvefwHuukdjMN5eN33Xg2heIw3rtQPB/P7sjxAbz
VzSwPc217s+DyW6SJFP1KvMLHkji9fjRYSbvfF5j0YeHHphQRGl/oSvuv36Lw3AtQckzn2A1ypu4
ZKJW4tjxVG0b2cHwt+jbGg1cM2B6NUpq1H08rBmOT/Ogb5dofRod6WbCOaLOcrokueOwcZ6hguEe
xXkyfZXkoGPlYizeqGFBFx1+3M+IEuAneFSzmLDGXFdz5H+nkSpdTtJp6NZj4IrgMC/KDDpH44g4
dwQK84UpYdReuAQ+SGV/9dheiuL3TyD99SvC+ZRpMbvMije/Zx/GXNtzp9ZYbziniTuh+mUJisy8
eZ3Z06Jx6voJ/xRVUb2b/1j5VOn8ZXmUhLMKM6NVWSp487zhV3F+pO5x30kflMK9uCkOukFFd16n
kra/8TivEdy5zmZlTbrA/kAGKezPeFdddbRwM2VzU5QVzM7rJkGz15O3DO6JiKET7zaoTksvzWgZ
oJeIwEf5yOHCF4AF8NLobNQchLNtq30HM9YGJ7dg8qfjDiZTROBlku2qXGCyiWHUgfrvJnMeJtCL
HWwVufZZ2nbd1JPFSiGz1GPLgr9iW+xC1s7ZnEh4E5CAzBv9f47JNUzfTIiDKhahwBodV1HNC8OV
OcEY3ULL8jVaFa9Mqpq6o03Rw+A7D1KBS8lVdnQEMokx0yHk9clTCRtUfXeZwDPPEU0+JrrcPoRH
Nn8/e26TrZP78b6xqEle8aZKZ3eWg1e3qqrhapuei/aYkJWshEe4cPw9Tv3F3BuMaUSxulAEdO6z
PcJLHBOlztT+OX5WzvtSa6jlDIpzlW5W5O0XYP+7zDvpSzRR19jC6QB0kOJ3j+Y0hGkei/6z4XgL
pyNYoiHAADv/idqTR4f4tLpWJCdG8dHU/CIu5yXLgIWJC5zu42/AXrkMRNCJqRG4HxCXnZW7xbBR
qZ/k8wOUm5t/MN0s4xzPfmhv8ypAzFuAYEBl/K59WYdhMdD9cu5yXSIkHH13mwFk4lWysbrj7EzX
91QVKg6vKP+Q3VV9JhS1ctCQDXvGgJFRQKAcsUNiGxs+togJe3YJAjnWo3b1F1lZz6FGyFYJWJzj
nLhcAvvFEouKi9te2QEtznmGLKWEn6Aylb/3rthlCpAcOU6rorPkV0iKSv/Ko4BeTD8uVH/hVq9e
PGqnNbRct7QZexL70TGsdMM0j4s1p/8bU3Q7wDmAszTFfe/pzTNLSMcBQ/Ks0ErNYxnA4/JoRUnY
dRM+GQrdgrH7SHpDPzZ893c2qcM7sUjPayG1KfMmGAWR8NEz0ZsFDP2SOoWX4VbfKGkka1OR20bs
061H8Z6hAuUZmNCBW1/bf76d+pe4TCZuIk5ck2KpVS9F64DPa0Opopsrj5WjhxCs16iSfeiuhwW7
vuxWJierD5zZ+v/EDn15BV/LPG7/q2PkMxBVqwacn/PaAgpDoGL94SMY1/WiXoOlOV5oE2i8UnOJ
g+Wb16p030aSWXJLWJqagEjAYpIoTGG3qKolOYXKP9rCd0NKJBi7HycVIDXuF7bo/um5Zf6uowFC
c6yoyyOIR4LJvxE5Kr8y5C4oPW2BrPviFVJHb02tuL0HyRq5zzPiruYW8QSE0TIWjO364pzqUuYp
WekHxQDJBpA8L2bNJpgjrKvxP7vBWl5ZZhvPyTRuKPxFRU8mtMa0GTBms3VrzniO/C/omrbgfz+O
6sp0wCQ9LFQO/KbLmWMcHtnbnRx0fkcoXkNwm62ZDpfjWNKNcX0rMxRa0pzjNvfZ3yV2cokUMQgq
+JCKOg5dc8MJfcqiVtF8UaUOKL/XEkVp6yZqSmwok7Ubmtmd8h59EHIlVao2VfLlO3pe6iP9DomN
Qwt1P7UKwkkw6nnVJ1jlHRWlnEGq///3Npwxa49kSJkBndOHb6vF3qS/x9AXI3FOiAZAlHBbyU2P
HFEqo4ZRjOkDxyTMqkrrFapJduHyZOPLRHt+xa7otlgXhQhMfkuBi4PexsKoTM25BPdC882lde7I
U7jFSpmku9kUPJggyuvP3ZvZTcRWAHH3nvVuc60IIIewPDHjpaXRNhEaTz/idC6dYcNa8sGV9fQ3
KZoZTQKJ9E5gaXXkQ8LajoR501Fnl/DBAdtgU7tVCXFU6JfzH7GZL36Amk1Hyn+ZBafv01IRNvul
J04REsPMQyv35tdFmGeu/S4xTek/7xajLNMzPe0oKqrmQNHmB5SV58BEu8DwV80Or0PuwH18oA9V
t14/7x/+PJPa4ji7E9kEp0LFtv49GlrhXXkSYV2ijw2G0lY2rnrAbbY+V5Ssoxjt7CTRkCo19gJR
e2usnAfkcBDBclzkYQZWT0uEaA+Da2t8M9DS1+wxvIxKTo6YGHJspyK6SXzlre/OOoJNalGvmZKE
PdcwBT5c1/051Qz3zC8GnNuQ2XDDNV+vtZaqcOZ0bvWq7iY6c20NBWs6jmJpWV6MzQzDLV10Diqb
8OL+KUfruVORXw==
`protect end_protected

