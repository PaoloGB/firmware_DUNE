

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
HSlhxG+nGNeb6BdO4J7IkitJYIbtBbsWDmFZ1spjjwtBOyAIYqwLzJC1ig+SAcTTmNsfCsz9Y5nl
2hGf4jr8fycEIdacpU8O0uNhXLUNHJ2EY11kYhag4WTmIbfP2Q5+C8Zn1fmsXm+S/Zj7B+FEo5ma
PLMSuCWk5Ke8lR8f6kyq0AkK2MMkDcuPhBPGcEHRyYiZsHcWKdcqWJK6R9m6lhT/VPUv/bqpTXDl
w9kuhcpMrpYrilDExzRYqxzQrLadCLQ2Ssow0FEQEA3AZVkqrFF3RRrB3Gz2LXMiTfbUAxlbWG/5
CVMM8+gNpiFlgERhmZi0j+uhwJdQ64Pt2AHj96nB6aFfylzGiRXADgb9xykhL7d7TQVCONah9kxU
v1o/gVc06zz2Hewt+BP5N/nt/Is2MVfSJiDnSMq6s05Mo+F/5WlHHhs8Ufi4arMlaGbJ8hVM5yk/
ljQvkdiA5bMXlgBsaxt1SIIyQObdYpSgofmynKqLVkzSfIujfjYMQ7RhaRMZBmd2dSyvjexw58KM
n7TRMo3p2ae6CXUyHNgEz70ALV0ee6Hx18W4Zs+U09WVNRlh43iWvLlCo9v08WSFdFo8ArExBPNw
MkxqSU5dLyRIfdto152bVfrafb6WG+SlyRUftkU3d4g9cK7M2TX0QDPQIyo3SWJyc6nLqQNG0SsN
O7kE7JSFQ8E7/Kd7yg1rK8MYmzOa1yg1HqITTBISLZxoJmhVTPKDV8GUa2NgZLeqZyT3GPm6hxB5
Wpo71hftXtxDTLCB8WQX9DEJPmH/c4x30RPEyun/AED1ih7tU6Sb9Rx8+xuBFl8GEkXIFxA/GEVd
yWtelD1gfST5PF3/VivWWZCz71wJIq9XzxMvs4HVY4yI0PZGuDeyBrJpn0jeOhk2YOfG+Xnjx1y3
p51YP6+yt877yl8q6yUMh4yPmOxpsJ90Vh/zyRvfjzXd22Fw+A6RM06kNXQhobN/Jhu1jG8lvMwP
yv/xrI3YvRdFjjmTf7kEIOhCErufGWgiLSOLoR1sdSgiiFXNma2+PV0NHHBiWailqnmgYJjPT0NS
Xl9UaZVM9jBO4SapN94uy39aIkcltkl0UEIj/J2TzPd4MrhSq1xXBsU9sJj4TvG1YLTFzW8T/NgT
MSkV7Ttc/rW2lcOgIA4u2nnwOKTFILd73RT+T7+lXx8kBvI2JJG8P4EVaO6UWL/n6cnZG0n44qHZ
R2MFLV98hAc815WIMeQz7sSwbLp6mH2Izljkb1QiDk2o3jYdEp3kvsU+mWQmssjhbBYx81XX56yY
+YYRP26FfaUjxVvhdYwOWlkJbpJH7JFIS+jbvAH659Kyu7XqLxJuEadwc5HJRNvmLvOPEvClwZcm
2EJOslJMRIAuMHDNIZTvVy2DEEL+bhF/ql5NgSLVBjRciFijuKe3MjG1paKm2ITPcKRr+OSm47SS
A6LfDGC8nCNk8LXeOUiTT+36BqIMsRP0IYuKFU6RM8udUkEO9Gfi1V9argAxzokXEaRCCFfDkRjX
JgRaTBeE2KmELDSiCdSzhm0wdUoaqCwfGiIRkt6OcNK2eq1hD14I2pOG2bVFUu9v+98Cozc8n9hp
YIArvR3+e40mRzr7OOkP5kuVJN5DXLbu03sgIlznzR7mp98ZZxQVTqYBx7Yp6AA5keOe509HvAqs
w63hT+Jr1zCNpcxf23mruawMhnVU1MOcnenVdK1NyLaYSS9e6SD9mD3IYWVRO7++xgojbe8YQER3
C8Ysa0kDFmpEuE/HlYUMIT9OpNeV6XH+1JDCJItS2wpX6YkeNITrU0w1KDe1y/cfULaGoZB8Qpxo
EZW/TveWAxuFVgA6SsM3LXG0si79E7uAvnDs3O/5ev3raYMRx3UIL+f1O4+yeuwOWbcTQ0kJ89S7
8uTn4yQxivnwsn0xCTxks+vJy7NCyiVPBxXtEsL0kfxhsfylX6ShnbwgL+9RBbjNuauvFeTzILhl
xF0IFf+Di1sRdVpqLeemEeiH+gAPe+AjiN3asiugzY9W1ob4n7clRCBGju1Ws9KcVgpjImbWtXCb
kRuRJVFVxiEi78zILTKrieZBETscZLY9W4xxavrimJEyvERhCCEHk9ALYcem+zvBA8Gr23ffQ84t
Ew78t4J8gaOCBUaAGzfbBMrHaqWu3/TDeNSLZh2vAwkg+DMw76pv9QKYIHcs5soxYbzbghMNQLGF
O6cbeuniRZhx3arQ0wubJULdkYDxohqiQNf0LAIPaBpum/XXxmxs/BS0B99AEYl60+usVrLMSwHK
FiP2jItbtsE3QMQJV2pnGg1JQQcHl4VByzXGlPM6a9jSyQWunEWUWf7TadpdN5cvjM9yJeCQiHmW
nKTL9akEBVMIpoHLBhcGsQsoNWcn/U9eKsE2z6XB4pMU4zwUoToNNvMYVwz2Ovf0/s9A/dN9f1GU
xWTKcBEDXGXUwBMqUXwiQLgoPg4ebysjJm41VqOiHtppjoM0jGTQJJSAM89Z/P0D8FjQHz3W2Gxf
MOCF62y7YY5Hpe3bHWZ9TBXnU1tSFGeDvVhHWuAbs3JySsVONL+OOg+/AnzvS7TUvq5OJ7raCm1L
JV3rXIP0Q4bqos6ieCGM+SNr7pxPAVLI8hoM3yPMykTVWqYAeex38shAT+zPmc+R7vIjqQ3Hjh5c
VDUlW1MATHB9j1VOFTQ5gpVSjfGYLzpTCWl60Dm+GaniD4dFr7KRN51ob79mdPzOD9XDRAsgAs3O
3oTYK1CR7wnMeCKCehm7Tx5XFM7FGtdTiiLtJaS73lwVI5onWIySlU25kEeW57N2Qx1NUcgfcZzY
hOsO6/8UuW8kxJCWTmNeQfLFsKp/BeagNHNzI3L+CfaK8EbWbaxQBRZtIe/VX17Rl+RDaG/2SU7i
UFCj2xiT1Nu1YI6FEkvafVTOSVMa6g+zbLPuQSJdkLYb0v1LHYhk81LKb4uDCDVfJ7VDPz4LJeOU
XXr9hqbf5vYajNb4rc1VeyqRaWd2KMQQqFvI4RcexnbE1UEhjjRDgrHOwe6WPMfGkO7p711WbBwF
k9oQZlzdxzUHNOsRv7G7VGdMtv3+RGyW8Btmo8iWZfFE7nASKEldPMB8/RqruAmDiAMxSDyL4yrh
W4F3om/dKHjYlx9NxulfIZWU84AA7uKLFcXHIpQ+TBBmQn15f71fCeCbnZb5kEfPwZ93DVuZyDMA
/QyR+AUsxODwAkl/TZ7BTL/2y3/j+I+aySU2Pw5DC1W2o+1AH9UT3fbv14lYpdxFNcViCb7sCZI8
E031RTJPlz0Igg67SudDgNqLZ11c6JOjegvWFR/Orsj38qG7h+6lKA6FOLT+LUT73KCPiwHGcofh
NaB+opxoyo+ZO0Puw7F8lYP2u5ccIEaH6rSabP+ZsVxgWD3WroVkRQPOGbax+NLWVgRpRRhYXEB2
Du/EjfACWhm8grw6SVutd1Md650+I8hIoNd0dAbAI3FcyzJ4CVpMAVG5rDgaJrh7TM6XKmUJ7CoN
9BZsUJ3fSobuJ0Y9aPDeGNmGt9E5l2uGJTdlHv38TIONaR79k7fi0hs7P05U5CZAU7kgSbgKCL27
YyRVBb7ijatyj4wrRfPBYRgypf+fA3aNiRZb5m2n8ZhP1awdW2j1wWkfYKZvlQcKX4fkx+XX9zDT
g86jOB+wmEAJGib1gkCZoefh0Aqgkkpd/qTAe5bdsF7wwN7upsy73RY4X+Haxtu/9bEtir0Dpu6e
QYzbKqt836FU+E9PYxPkitP/w01xBBHyfgtY47xPAQIFWGZ1LI6ofrRmv9YLnUJ1em3Ct4NS1pQE
RdhNHaIcAEqEqxQ7ZJVZg7YU0zApxYMxMyQxFGHUZ0APSUyEh9E+kY4Y4FuHl+0KqhxWmqJHlGwp
Hoei3uNg1qgUl3azpTjgd09NUfXMdJ/jT6S4IhOYVa9H+v6Kte+ur8PLHKcnRsvZ6m3dmOeVKQAy
GGma3O2PMwW2DqsSe836Pylw0BQ4S3P4OCeB7vkp28/pwZVR8AaDZNHpWiSL3omWoDiFmVsIIxgs
cPNbS+2h9rsM4Ow5wvA0cqwi1HFfkROaFnklnNBgP5+vQ5SHe/jy2L5E6FhAK7XonIR6KJ6OjIqp
0McsFuF2y0AtZJftjS50aI08t+SqRfJdiNufHMzeZeFzgCzWQvj1dPuNY5EWI00cjirxFnSlINf8
I9bEJEmgpA8POfjE8KGb63LDPlhyS7bofZDqBz3EPSBBNeJMVu3CmKWZEfTaVyzMY+kk0l/33nks
2PxvZ6ojT1SI4xloPlOkYxdl4XjwbJ1v5kKCywjxwb8XgsPn0bNnkTanMMDH2g7NNuO7+yNvzAig
zdag+XwkTIFAinxXIWxyYU06HkWZ0at5xtCiZYBgb67FlyQga8DnR1gwOF2LBBznCnkomJqXIlG+
tJb2vreqaInygbYxCfHBK/eHztSTQxtP/rBNWzuZvwKgnXuvaIEzj2O9Ox+mE4NjjQH0GKZegnw6
p6sItRoTtyecAKXPmnhUNWrMh4ulRJWD48wuY2R5tRlDDn6/n3KXH4MD5jW090GFyAtj12/yC6+H
SyIAyQWvFy9zQsAEqyXaLL0Lj02+8AIE49/XOiSAqSsbpzvBSozoZhc/CFtocHBKz5gfOPOV8EJa
y8zqADUTblLAiyis2Pf6dhBZUI8FPHhLLR+/kjNkgCCAyGp0wJMt+CJrtMa96XFVi87FTj+V/OuP
YXpV4wxI8W0ahT0jyGvyKzzOq1nlih4+R7/mipIXe+Hk0Voigr6FPRqZvmXfmVS70sLt83SShyks
LtaRBaizMRQRv4TtpMD/omz+huPE6kWCLzpr0FcjMwcn4ZOOTz+xLLeaTnLkc52g452/wFgJuaPG
kaT8HkfXy1NrBChK72YPiVaaIvJGLn6xNqiaRb/rqP2xc2cYMSmyLWoQCifbSfovBIuTqrCtEY2k
ieFVS49IjGxopBfsFfkkOGFVmZVFBD/7aA7L1G8SFx9ILul1N0XQiM5asZgdKLfUMD7Pespu68bg
BNTcc49yrpzhvGcOYnv5Wbn91KfOhOPqIHFOhdY4uCZftI4ekTeYf0M7w18rbE3WkzzU2cigX52F
4J5SEVo5MdG5jUutsoRMBJ3NHPlHL/mDZDi27yC5TB3lkD5dXmFWkpYPFFAOVwI45GTKGDMpsnpE
wKuGVrpIgnUO+f4xv0u+VtIAabe+mkVdxiH6mygxTHrF+NYAvDbQ++6ABuNctMyXXjDOTxCIAUz8
I8ZRXxM/C0/dgisv9N7hlm5E30bfW2SArEljhiGosTVjzys5YI/8JGqa+Dr0LfoNTz1nY83vj0c5
LulDaO8pbNDSYPr3hZ61fcDlQ36Ko+zPK+B2OyR6kGovUITvHhvitHFkGo1pmi76zVr9449EtZ/m
9ec2wqDOaWbEJ/N48p3fHvLblodPDBGs+BjaDh5/H4iEfpJ0xM5bm/NprwdC6EeMZS3kvSJQfme/
/CMmLBxlVLicQbei8Xu9nygPgNv1ONQdDlF/TLI6is3YCWLxvgP0sFHeWFPfEPkHi6505y5FoUjt
ylof6uV4tGltq4VM1DP1nJxuYxu3akC/5K7Hz3I2ktxHAROYYAG6PvIyO9Phrl0JR1fNlaRS5xlE
MarGxfUsd3oYpbIZ+U0XR5yzslRqMf2/Nrqny6RQ8VhqdBUlJ7jVS5rWm2lDfaTeC/HPKOLPteFL
nB0f19F8PZAin2a3PTw/X2lU4J208MlIX7yf2XSkxtZPdP+gVjR78smuSXvCOAtNC1PrkZe6joE+
8i2DBe4OJd/8CWmQJW3Mihp9R3M3wJydINc02hzMBnf7e+7zpLg4dD187Bt6LB6t8DDw5waAXgoL
dX2wX1WqBM5FtdMNjtMF/O+pvzFev+3JknmY79H/acNigyjR6bwuP1E97/Fhzbu1Cl2k/kq0Bxzn
slLvI7rSB/dcnfQ/MfPQvF8A6s3Hx+zp+MmE3ChoXkv7XmEXKHtyaW/5Aore3L7a/oCBIhM5tF/r
Is1vz/x3e2QHOwGtp6c0qfSxSLn/j8x5+4JGUny0zgeRQIdyfI8lz9WdMj4kGY59ludP7U9SHKS/
59NKaRPTqfs0C+Dx1RurXzeu+DXO7kIQb0BBXu998Voc4fIGzhUnYHeA9Xnb+qT+vG6Ux0HYuBiT
k/h0xBfO4eP+czzldYPH630B/zpxzSGq+iCmKJV7OG95YHWyJqqc2ZQ/9vRY8WVglx5sZP1XQRqH
OtEeyWfFZNiGUEp9HmRIg3zLi4yuztP9CVWIXyxM6J9llCa4MOnJRRcwcxflXsfv/Q1EP6t/jHcc
LTLBjwCJHjhqJW7GTQMtrSehnKlOnKIfyl18Q4q4C8ziamo0Ybm4Jh8u2IrAcdv9j52JdFXN8fMx
GL+EghQZ5iw4+61FnUdvrcOM652AQju9Jyd+SXdUU3j0iA0ZwFK3GuHWhuK10eLkZE5CE9joUn7a
np0N3IgzAV2KVohYfCtAbX/ei503AKLbJy7wZj5nLb/pzLt/+QdsM0bfMqP9Fkl6l+vKIBctDIZB
AO0abX9ApSrfu/kKIZWaf3C9LXtXMM/eCuOJmWPcJKRGuvB7QyN93VBcZhx8OXeChsvX0apxej8G
U4NF4BgRl7Y7UuB+GMY+fBaryPDZLuINUdCn1OYVx45SgE+a6IAXQ/5hszYiEVn/eRoTX6YrHeNk
gQivdpoz9tDHdml8qcVFNXEZCXuIPjMaPWSX7OnJqq7qWFLwgGiFCepHIeUueYtHBAEgLwvCkUEW
6f+OYuGaqp9p8tAwTbjWmXSA3EPguYigG1nPGcjfkORt6h84eKyJAY8TiHhVdlltDAV9KOPmDXnG
iwXHClmwTJq5gwdyN2Yk99gW0v6TaKCB//8ly3Nz9gBSxi/LZNfLPe7BZF/4W1IzMgA8i4Cd3wki
DjdrzYV+HvCTCVeTClK7HyFQYbVOziUENOPdZzl/mBDT21TCJhdCXD1ND/C/7akxqqbGSSAnZZVJ
UhWTb92Bklsijwwi8E2NCvYrYYPDh77uotrIJ0UPJN5jfDoWEx/V5YMRZV0IDk3Y6bFojfG2hVJ+
Dosa95SxHv0nr29EjEqwFcDOX7kT4cQLi+CNiGtE07ADHuiJNccUEQFJKopUeoljDBr0RCP79BeO
irk2EJz235t3lPqT1clPrhyzcilPYg/q2W2s2uumB61Qc1IbGYiJNcHF6jEmvXAjhgq3lZygHKNF
zAtPfEH5TjYEOmgzgUazgI2VLJY7JHIY8IxcLZW42NuKRv1WmnJofL1YZbttgcksvDJBxANQFuPr
72pvTGU91Qs3dNFZ2QC5M87bhCWk37ioJm+QwrUwibV18esa84KDetFBSHtX6oSK7/e7nLLsI1uC
HtGuH8xca242en2RljpRdFIfxlgcZw3d2XawfzOLuwp7+wti8mxauWTWzFEP6FEO5eRfLkGgqxiQ
zdgBdqiyD4f5jm6A6yfZ24sTGh3FopVCLjdfCeKCtvrRjXT7Xb4BPpytLEXFN2pY0GTX7oynapB1
ZSxx+1IZDKhSLY2cRrXAzS/BWyA9LIMlDGlDZFvdQ0RjT3uJE1U/5/XMcJJBGVRIijFQdrMBu01g
vkVvvreCIQoH0jzz65nXHtL7GPUpnQkX+KaNCnG/CPQoL9IJg9Yyy2dcZBnedZ5jfVkkPWm5hr35
TV1dyE3x8BAUiHxlXlzkTKEyeobpxuP6e7yBIPHBI0coM38FUCrmSy7GOm97ISPaBsH7bTOPr2JV
t0ANm33zMCh4m2fWd4fZp7MkuiS+SLSNC+7ciLecz8viUxOcreV3w2DNhYJ0flGt1Xv13lxNVFro
S6L+w1ReFMBHshGlVNukwpZlCti2pCDSygosuVKBgs2rYpy1zGUwokEEeml32uNoypAFWBfYDpRh
BucImuVmJ31fUJrMqQhVUTnFvwHwpqetVvRWxtBsEh8pfmGJlgk17uRFhZo1l0hc9wFGrdJ5SPjR
nD5COZP94GLrrW4b9HXXXkv0MjDRhDIMsJtxNjA+gtt0Kb1Om2tVC696O5gWlUl9WznURBxUZzoj
8RVAPlNLnBHMF5V0ALxWWlXK3urRNnhiiEDMjp+cILMVOpx4zQbWILJlnURm27ul7lCWLE06MmiV
1dHWcTFtJ7uE0vrEtG1u3kqoglt4B9muNlkEIn4Xb89LkTdYgYiXULadZdZgf1BbCLeDS4Zz5Y39
zXRFJYm0Ab54vljlnwOTj/o7XQlkh1MvkA+cXGRVmAZs0Mr+0z1A7o06vZTfBzqT5oHG8eiBQ24I
pNbTMLclGoj/HYE2qE2Xi7GK7xiZaTNHWdFHUbJqXDysVObSAYndR7SstBni3j3c698it6AKKEpp
I4TPaB4YuFDM59S6UqxEn11sBmy7eJi1WsqZUST5SiqMtQkXBdW3oQEkicDio0bEBhaAMLeeiuag
vCpHxlCxpSiOJuq9uosGWNHUOBDe0tnVCRTzLam56wRIrXhukAvlUHJPugw3n7TKu9wkwCL4VtP7
nn9IJk10N4v3OLzPRAEXoo7Vu9bbiPSfCtr0sD48C6wnlbtduQpH6H7nFzsF/FuCBuknXES7BZwV
Dv2NgJ5O5kWEf7M8EbT7qWyyrjQjo6msBkJTzPZpxYcPrMIwRQqlCt1GA81QI8lzyhpfxHeSBizI
UUlnXduXRbnGFIeQLOJNgAuX89ZNtWists87SsnuxBbWI6NfYctCt4Vwg95IYO8roUP2lZpHb3+O
wTy0Z0kopsQ7hg7OBZjxlrXjKScOcUNzXrTklNO04PNpo7Zhu1OBQccy9FiSe5QfAMZUJCG5ANU8
HZ+maKVxhKIyOVsS2e04eBCJMHzApF2XNPELFWAcRJPaUIqXBqeXrjQ6VRCwNbwtqWfndXDzgF2S
ICh7slnz/5MPQpRvskkUglK7MeMpUvz1vAiG7dSHt6Rp9o/+MwWPfueJcis/2GVQf80TEYjfKuqd
1A5EarXnmWcTjwZP52BziZaBEmo7R56IR1p71syVBqfHf/pAb4iJHyN+JBMo1HtjZqIZypoXCRLT
vsGAexikwHU8ViL6tWDmQ/SWAw0JKaraFYw7WSRbBsj9b57PgN2+MrsAv+7/neNdMyfXT7mJ7FvL
Es2c0nw6e/UuOq0ENgz3x5AJo7NXDKwBLfjUd1WyT8WqTWb0jAxSB5Cia3irmqa4oDAAtxuwzDjp
wvC+YTyMvsrApIBz0hSA8zYvBQK5yqQbN5rGLOYzAan8BDpNmYdM9R9eGj2HLSRe+QhDMqcVNnA3
wFVnS/b5Gm8uErRXQ+iThlCZ9sDHcQ+YoizS5PjSbCNdTvWta3m8toxFTPJ5fryFPdDYYTH/0mmI
CJmk56plXGSgPtcCjfzs3/KJElxjrytcK8CHrEYKTPIXREf1eJOMoT3cMuUmjttX5LG/lNEQYfLN
LLe5jfJ+Mel/sw4nM1ik+GWeMOAcY9pHGYaE9ilRw/uyxYEnBsUWGkb88pNzh7f0nxg12v2JfVTG
8Bu7LE8i78M+vcj6amQ9gwexOf4foqvujpxn25FdRgV8bEsQDt2DPMt8Sud8YO5aJVjz9MwcJVWP
JQwc8WDBVJbx5gaN6zw4TwoJiDpRYB5FToCQf+9qaCDlsbU2BNSpQYSuXh6weKVUQV3ykyZcBx1p
mqgpcodUfEdetoTNvlqU60OMJqOUhbsaPUguHchWagVuFaKdJrt5zmvoZoN3BZimx3p5m1c+7k/5
hHJtRyz9WVeMN23m1Ul/YACjWf1ApPf1RKkgejni2gC8uOn22GIkuFv6R8LEMOX2nE81vcyXFtS7
d9fCVc6DqQy8nM97pS65SxzJDgGTYOq+9kRfokLIqxTWwr4Brly4tU7Y9VwidWB6J75E7WiMyksO
0dRogPxE2Q1xQLSfII9d2zxIxjofN0RwzNnV7d4vyVPen9jQkVXcPT3UGdJj8DKFs4TeM3VUqiWM
jRQDzIDoY29UA8ZRmTMdv4HSqyU7BSDpVBUv2vr8z3aWXFis0IGMTYOKfykNqeZBbQ5s1FNJbZB2
mEXYJZZbgpEUjX0pRwBbRp8JOURGIUlgp+U0NC98INnHmmn/1eg2r+aJHYPZD8wAhhrcSm//T8Y9
dQTn37z/pic9hZ49mbY+CB11bf4aP2oDE2QaGqda3Edm/hNitp0HI8frl9v5DNsl+tOP42A05wRn
bIzplv27hrMJzE9WQnPF0MzLUfdymND8LKhyD46/uf58Q1vbBvVHv6peI4Pr1dj6/iju8qoR5lQf
ztgZAoZJ7T6E/7qPAxCZ6X6lBeJiLATp4UGaNBv4lFSAw4m9HLotU2t0IR+++a/Bf/TSAB9gb35M
0j8COiuSTMJvHJRFBwWa7O3Kk1jwITm8qVFL+/E8VYOGeA2i+PYKeMrHeml47sbUpWnskNiUCKtI
iJhybjKnO9c9zf1gc6wfDEG03aAqVafBvjdw2yJW5gWKroSrSpz8ADwyo2jM8ieOkPBTbemGZEwC
u5PUJ+IRMgL387iAfvbFZlRhuPrIT9b5J/axMFJqmHEmdFu1lwF0qNfhiDWZXbGGSzFrCZMUqpsV
9EFdhL1bC3bOeNNJVudolr9NoWqEN6RiyBpuxHCVoFr1+mCgsf4j7Y+1cPZG6CoshfYPX/SDQp0/
Mn5tMTISlxlBaxsNNjg4/R+t/sRzWD/I1DW1eO7Ik3eerqT0QRAcar0QPgoR+SP2ykomum0WZ+n7
lUAT8aFBkr2udrY10/YXpBWcHCneixOf6iuhDPStBkEkWNWp2DmKXQaDknyA2wfwTGXykrhEfZ2m
++zYU1lMMDx9ZpVeK3fk4zt9+b3RwN0ZVcBoP7uetBo3sScrUqQ7bWjdj1DsBpw02KGrW7fDaVU0
LjjXeNXIEc7fZAmW7CGImDKH2ALUE9Aexb2+/65XFdCwemy/RN4OTNb05bFbG4sCpuShbT8j7WMD
1Y1MwR/mSIp124I2F4K9e1b2rpuW5DjH7FattVqkMWkAbXGIL4ZaAEXCjThcXM5vwfaKG8M5nUou
lgLazYlWwiMpkt+WNt4Atmb0pJATS+gfFyA1wLkATPznSlwqg8Rbu0Z8oS2KFvXZwoqNmSHoRe8n
IQ2hJF4h/zuD4ziP/hl3ZGEFbGVtuXyi9jmUOiiQvCkcV9ZVgU3jdydQSXm3Ldk/SNyXTw4zjt1E
OhBrvzlPp9FU6cTfz8Sl2SGuVK/Hy4w/b1hWq7Nva9yku8zXNbHUbCu3AaD0vVMODHdCmDSvIpEr
fo5IzviTXhjl3UIRMy6LU75KUEfNuzryUiyE72fR7tB3uIIpiY3eOJrsIqbRcLPS4ARmu8Fe6Z0U
P/ku7am4etm4yspA7BGxE4sFknerZIZvr5akOiILYdHfeF0jucCkhkPsScJeXP/6Z16yqMrD2lo7
4FR7MaFhQgNT0cWPEBOffDgKJUpUNOD/ZuWZzdHnfeJcl0etFCILpQSfmhHiACQAhe3JwHfZWj+E
hZndZzONJscTK0ooebDGnV5IRzd9202OJS+CybvvKAs8iUwmvyA6PAZbZcNmp/a27nO2xz1Xzpzw
xJk3T8hI6oSsMGLyQ3NV6EoI/AJ82u9q2f3yWm8w5UMJdI+2z1A/6L22/ehDGh5PAqQq//52OrRA
TirrK+2DnuhS7I435yStlRqoBe279N+BsNTLUMSChtKmFr9utFracA5ply52fKMgjlTQD5O1Qp1Q
YpHSgwR0WQ+uz1Zu/ko7P4Eht1RIvXtzRXRB8hRmIfAjvHGMUI64z0HWTZfLxTeoW9dsrwxTzo4N
ayVhILIAhwjzyM42aS9MvTCLew4lcGHQO2Uxt75iZg+6YcbfgCUGw1YPn64L5ryf6cuqi3vZmwnh
ZUxsMcpATjnE19vAQp9pxl+1hBkz6Jh3Ua2a/MvkU4io5Rjwz/wem95FkQEyD7oXxKwW1BUmZoph
gnBjBcYDm3A0oTsxjusdGggnbU6y9yQLbyPWNkkntcnx44tYfx+/zIeU+Am9AMQao028qHtsxr+C
9+Z/ezHdBeQm7Qc3cF698LbVJ676rRyWhdVhYXzklbxednxTELeCxOVy+0eGy/8Uldvx2zzjkBIa
SjCriaFLaAiaYj0+svrUsd8GWGexHMEywzaOmWPs2vpkDg46TzwOAWqIPMu7wzoB/6PwY9LGWHK+
VaNOzpTP1elgjIssnYNaZ/yPn1B2nBRjbB9I59S+2TH57brXCIV0ypvLUKceqz+xU9YbSeht+15g
Te4Gh6AfFIaOiRRoiNjMgtfMu6KHdJjHHPu+8dWkOHUp5emmgrd8EEG1rfglOVSnQSmo2C8GLxO0
KmuzDN/nCp9mmJrPcrAAjW26a0xkjrnLvAsCFhHnyEXoSMpO8DeDiiEkqR2OCLjl+jeG+DHixnmG
L4IDxAgMM9eoOAkplsYLpS155Lu1AAdiqnPKw5NkwuAFKoLnJFnAPqw4AKjfusOJEUZAtdMmCE1O
W2I8a/Ov0Om6EbCN6Ymm1gkVFlvbjjkYwwVV6RT283DosIqxFwQeaW9c+7NxyLPW1HW7FWAvokBn
QMHO8CxYD8qUkk/L8Ydje36jzJWJZWrKhfotPYiCTZURlKwExubbGvc4A8Wi+4/KKlrmSXz3KUPT
r20OmlkFReotvgB3G1DlqxXWI6BXm2VxqSlBzUOpUgUGoOQLodZP9Bvanz93/DSAYh80q6AYxFFr
Bs2XhyAkmkZ8ej9fY2AYIKunhpQo6bDXlOqM4iCL0XuCw8NXvEeaSbmcPJLgFwIcOi88nm3tYjxX
XejutDb48d4XPRJaitJ1LLK/lLyQWclCuWvA8PyqnBrWZtc4b4SiCTAg4zdeC5ms88DeweWzTpsh
alvJ0sBtv7xWAWtgJeYX6QaTkbVAqxIo6wyAyu848PK8jgLC6jgMz8/Wqw0s3DxonrWMeaGYBM4u
uDevhYqObMGcDfipRViph2l/UB8mJGl5jmxHsBkPbD+t6haDq+MrjHQKRYNHYMhLLNoLMNqovjZi
hcj84Jf9Qa+gmOHG0j4mKijWgdX43VtDxqwkCQ9gAu+HRciQ4cHuS0PuDZtVLW2ZDN6aLe3IWMyN
1NbDq440s31E74SVd1UgcW5PTEtu3MASJ9TplujSNsUQEBEAcb5SArcDoyyMu2ei3gC3jfxI+Z2C
BNxUbAVl7mMuuThVUj7ksXkB1ajrhoxNzvAFnJ61t/PkK367tQAnG1PMsbnJelDApCaHBS3N6N0H
OY599HZdo1Osk3mKLHI0GeeFnhhgOjBBHIBeon4paZLP/G522XDGBKxanwZ30b2IPcm6h7bmt2/F
sKnxHeed8xtdig8AsWAu0fsDg3H7N/OJJ3uA66pskY55t6Fw96IXcEjBlaa9Ol4Ziiwgt2shJsie
mjag/vpzml7RmZE6iv4075lbB5d4QrxzP7iJh4vChGY6s0CBnMpMyD7MP8ZfsLlQGj+KaI1sLjPG
PXYrngmxjRfk26H9HB4hX0MjeFGTeD7BtKHOxTjaZgFSIcH4/HUBpSKArF4fma3v7Ohb3ceRX33r
7p28KfFeDFr2z+XoHfHnAMKGGCchnQicfbALM0VRdVubNMC9LuVwkOykLSCWHQjmc5agrmv2zFoR
31qDC2PTkpMGvjLADigAxHnHtzrUuFUzSn/kfS3F18bXyQCqjCF0+y8Z2mHAg8HBgVI60q6OIXyQ
7ej6asORq7O2QRQtEvSyazNkFOQXDL8jVkISpYV8rsVOf6fVLpZiEkksRZajZAX0hgdbQDhCS9FP
UF7cGUN36PFXZOWAP6pysNO5wXQhwjZETiwwq9uv4gnjiSQNhKQnpAhEdfEYFqci/6pWAVZCQvbM
GKJZeBBW8wSAcIttNnxLrSHiZAps3C3CirvsNwUD2Rx51PV542DJbYU2OGJG+ewE/rIzRVGjy2rh
313iX/RE7JOJykMLG7u0wLpmTWsMAGjn0sz6MBk4N3zUtapcmtDkaHn1uapdH12LdfWQR7txXd3J
lWcB8dY0TclYEh2D8AreWfzuWqOpC0eh0as+xCTvB7GY4vufBX2S1StFlyJTPm4zfXtzawU7QynT
A46+RcXfJ4FveO1yRCsAMGx92Rqaz/3tx466q8mw2zgBbpuTF2aZ08YWaoJ5bDFp4wKGxL9ISCcO
eFdd5m2wuUUMnDBX9zrvczpa5nbZqhe3OWPUFSoGaoURXP7HkQ6L736/uBx84EdW35Q07ascsLb/
94FXn2jDM4dv6XoYcBw2GECGFWQ/XztpZ9psVFSswN/tAQkvGnJzhdgwZQgcS1nnn3mE6PRTDifT
au/H4daRDUy2gTk9CNFqKlgqVfEGKn4sQnlf4GSXtE8UX9G3koavNjJwJ3rXaV4Pj2sI7nbxcqhm
G+1NE2Q/b2iA8f62F7euFTrcT6w4LDou/10wZbV3hSYZpvsjR3E4QwnWF52Y71fncW7SKPf95KjL
8/jl7d/1fnE74Zww1fbxh/rP++qZC4pZTfVVCp05c43qsRK2YjpyqE4cVokr5ps0PRhZmxWF5fMT
Qvpz6yQVGHkxgiccQ5KBxPm9/yF8+tPHDYYHe4zpgyawV16kSejZE33zAcNRB0RKtYn/pU7DG0uy
IfcchbQyYkCIx/HciZlsnXKlvN6ZSN5kxpxEQsPPK4UF07yKSh7euBsvFEo3qFmMVv6BRBfpb1Sg
GrD7v6EvHRStY0vVBUkQleDy2rkWc/YZt5SYKtcqLsUfUg4ZyYoQMI96c7kWlrxLYpDIah1hM25K
pzyGTVB2IYCfA9eSM8K8WJcX++3VDTTFMPFgH6ZFs7jqwTHwQ47Lk6OLzqkx2OkTgpZeQ7CMaeh4
yrowu9T71xvGiuppWHoa4ZxGJVAg0Oznw3/gwPYMFGi3uOCQFcYsqmVKlQyl6sD04K3XSn73EVP6
HXfrUYvKlu0lNOLmH0iObo4pXaloe6kOS7CfpUu7D3R1y1uoKmUHBUi5EZ0z0Wr48MZgsuLVwOxo
u75/N0LRMyfbhR8mCU9IEBv7NJgcnHyAwWq8QGkFjIQftivf1Eed90tP/bQSLddhjsmpubIQC/zA
wRQ0G7wkp6IkazhM914El2Xyz+ue3ZDOQiHeIbcWfDvT+eAGGVWSGC+Oc8Zeo8RYa8v/Aaf+vXij
GmCV1oZO4IQaECbrkSC5ZP+A2E+3ml+mfuZFTZuNap6hjCPcdcqxStHx161b9q/ZEzrMuQwdefli
L08QvXf+oyEHgqSYmEqUUYiVkQLLiq2tuDhWyvFIc+itSDK8Rqj3DzqHsuTiYbvlEh+W4m1peZs9
df+KPM5pr2nQOVI+tZyHR/ui8cUwPGHdVsrIEtZwPQrR7fNY2BMPG6TAmki/tmnVd94RaM9RkNY2
Ahvu8xU3SdEArdsC8MWBWZleCVavGj7Cfdl3aju0n0tHNHS+WAVLlOZshkOA9CcHLkNkCqH1I7T1
aEujOwKhafWNv9Tr78f5vEZPcAo983oPjn2+bL0oh2OzO6DKGXyPLQ1dZCHq3n/Bi0zByStiJ2iO
JdZN9dSJQuk/tFY8qoUaqb9DjWLFsJHCyfabL+txoJB63rK5gK+L79fJX4PORMNQcElnNyqC/9Tf
hYep0PeZwIaINcAyBPFWSlFiFSzgFihjYZ+NvJ3j1ojg1N31LlAOfnPtO/lr27woXgHKNyatfdGt
ZupGu8s76H/39bFFnJp8pNncPzrfbnaB3c0m9NYDg3GBVtsB6sN0YzbCh4SI0Jj1zZGjEV4SSn6I
9bzMAeAoR/itNAQ/DEf5u+ypz/R3VegtrtAM3pNExsLTIMdbsX7PK1v507ipURA3HgFuackRB3TL
37HRa+w/kkDhcFmQjM05mr7DjoLduMgdDseCvndxGLqN+gv+zP97idP/Ujj7vnMymuAFshiUIZMj
IqpV/7JZxM+dae9vVWmCICobqDx7tcE7RI0sb5QkhSlinPYyGxKHcQbyBH2fMyBA8lVLswJZE+XA
qCvqUxhLYCtVnxzQfYYq+gDykyogUv4//9jxznt8C4nH2TY06HnSuZFvVEiKKR12FhZ97iMoTSx9
6e8prv07+IE9iI/OlTFYnoSehvsggAx6ZNvtmOGcJJkRhCs198Hxs3mMMLRQoACoioWGVfHRtoPL
M3+Z65MZQJNtfmbLKPQLIejNp5iyeJztJ3o7D2oWTYD1t1vczp3lehnhPEl/uHdDPc4uzvRvqu13
tlUuorK3EeKYJz6ocr87W1ANGVtA94ZYvW5rn2+tX0DoRrVCRsQHyg+rQ6Po6t4XijY7PcKDzG0W
BpbFx6KYHO4Sglvk2zFkZONj1rotMyUPU/od8QURudzjfw3z7P7XcoJWOWmtETZDTN5nQVuo5bLd
0Lx5qEnQEbEEW+5mOeN0l71r0YtR/c5VA+eCMSQuCHCB6XNPyckpbBjGLmnD0egGzYSVh1XI34AQ
VCVhoxG4iwaFTkhk9Ds6t+/H8YwPmGkwtE0gAqlRuzNdgp2LarbTHg9qwQDemtXV+V1ChzW9bPFs
8w/odncov+4t8nocZ1JSVc0qW7Tx8m4f1JQsgJXs5AhgUHurU2OwX8unsd0ePdcIpRigp7pnPovy
DycpMpx2gV7NMkjXuKtYVLtgkqPDpy/xft3lB+2cjuCXuQBKOLAuCwNrXj05ZeHS0i7eg5ABPhdR
TO/JQgwwBYYHm/QQHwZYBe5ADFJNK89zIPW4ZLBz5VIxONq/0H2P2rQf5m2VhNdg4PN5UsyFIeuL
TFpoUebo0V9uWAdQT6EkPC5A8Ka8g/KMdYGXce0rOthpbRJTqLCxRwPQAkAYWiGkuBjE+ho0p7Bk
ZALCm1HOwlHWY7dM0YKCg47In1F6vsiH0SHLnlhPZibCAMYDQMmUsvQnzZfsNntSN4jkX0pAnOhp
IfCsJdOVXzmVDbpUrKaSgHxvj1dvCdniUtsko4emIxuu0bFLCPTNm/5EdAr9UheGzCLwOUSdCWjZ
Rtc9i+uS//KdD+QIUvYW0wbXAGqHPaiuvXXmUcCMOZ/qPVirb4G4DMB+RbVVQeQKRJIeLy98dIIq
pClNYfws9/C5eKJKJUDiZsQt7r2vjR9JSURxv964A5jYSx7Z1fAHCbaCFeNhOmBIQxvxivQm6KGc
NGXhUmrU2hRSIolKT0F3dteIPOkUqVbNKNJGdrdN0yE9qSVPj3RxKG8R+J85wYS/ewbVQW4BBqOt
+aOv3XtGKlYs4B/d5tedGiOd9L6lOS6cRg6lIIRxfdn5LZfC2BlNJxY6GUN0zsJfzahEF/1aRYGa
u4FaN/86+sqAuyfhFHJkr7CfZtVEVDQXHtK525oE0UMmAgCtBvKF25e2BzuV2paoeZ3o0AYqQ171
9n2v/DvgBqSFmZ3pUOeOxRuL57VRStigE+Jg9ABVfKi/iSVkc/3V2Z065npHSvkAU9R8lK29cv3J
ai6sbTfgq/IMqAPoUo9KZJGjy6QolveCEsAST/rJC3PQZh1EzKJW2ESJu8oXVYWHDmJtMS3m4aAP
J+SF/1mDevqqtgBlz60WjJJcDb0q3fN8ddW4jwjNl0HV3OrPzpqhWCl4aEJRtig81ByVBg/OMpJ8
zirdtGr32l69KiRLC3Q36WnlYKhsIjJ/eyFXCyNHbFITXJ6z5UWH8kF9ojVYfvsW83KuuOcXxV/a
Y09SkbOv48QSbb+JmBRRzjkO9tx9GrGgD7nb5zt1f1ewBVjdL0Rz+lUuRX+djEoixTJp3bMj6Jpl
Lt5PKM3XI9PiR7K52XuXFLDioaTdwWxvLgYneLYfxSY1D2s/SR1FCIk6IxQjlM2vnIv91uND3aJh
EIvhBy3AlK/bVbrYFVfxX2hT9i0lfxGAktgSq5HZPbxN0i2vMR/KEmHjyfpwnQUhr1rWTO/rH8V4
vTjp7NJQaeMu61ml/UpC9k91iUnZbM09hO5t7CThPwCZcUSBejyf1rc+5S6xYcgQeESqWoH/9pi/
rEB0ZhzniU2ISHMg9oGflKtpfFvaghP6i/YvvE1Fe0MReyO2GE4HZt1YI/fF2PBKBzmXGoSMGI4z
YJdUZ3swwki2gf6Wzo6Oszzu0Wb9z9Rfl9tBM8ieXFzPe1hj874kHTPJspUum3Zg8oqrSnyZr34D
pByfIRHjjeQqVLmD08Vt85FufP1JpPad8wc8zZZoLBM95d+dmmfoRf64fZtVkLOTWP1axbAGFW6K
rgcQcEgRk9c84kLpHgG1ya4BkYV/v8DMPdogMcPG95j0JDBL9hyuny0nY0MGBc3lSkrkzg09UCh5
yYzW5BIeS4Fy4WG6EpmVGbJm2Hk+2Lw0SP3XYuujb0RV4gQn9FvBZNntRPC28L76wuKmjP841igg
fuqkDSmw14FpaqaTeSaxJEUJbXX76XTRWh6Pan58zAfjo8sxbHAgUsiiyO1t8BwPuc63TYmiCy43
m7ml+E94IbrAMoUdlZnPrnb55MxslbTY3HNqUVPxvKIeBMGcm3+dlntcQgNtUG5ssclRuDcYMbVd
BjqHxo4bQioRoYUAXrEBnY+3gxhZwNAuHrVy5MFvYMhuTEKRyxXHKcrP67Xbi+xsfOenR4VV+wjW
feDyi7syAQ9p1US26Jnjy7GeZOV10DTfA76QZSfc24+fhMPBJN/aKnzSXuwIPSNN/PmnZbQTweKr
YMenxwLHYGYmueKgkGEvBg+vCNRjjo2Dhk5cjgjlYjDPYEJGGBny1GUWH+s820qgw4TupSnzYDXt
XyO+qBkO83i9dqTzK2sCvbyeSe2BJS7qOhFuDdXjZls7Bhz5jSyTZLnSOVrlh55xnFpW5wr+ntMZ
uid+zIUx79qFPZplXJLblQ/vTmT4zjYMDZCgGF0bewE66jLipRYcMvG3RxS1AMuKdUfz4eYUAhaG
8jMlAYQkUlzg81BN9bFHoBTEuygr3yC+Qx1u1KFx0nHMClX+T3NuaHcnAFkQcqVSf/+Ck2vHUNHc
pLBqQyDU+yheatMVRjmJImk2rPde4VAcd9VdDuPpDRdW/QlnsacfQKUmzR2M9JxdyzUsxXeEM48U
DeSkAEA/imaqov/BI/FxeD7jfc2UKhVvZBFhdBrh2cVQwU/0d1i0US/jzQRkh6fZe72UXABK+2CY
aVj4sYxhnjjstdQTfDyZNa8nI6EZv2saC4U7Y4uneFvMGhkvIqTiey6GEUYSqB5xuCRYSN0lDizk
3gb9AfnqnIxH4cxaNYNPu721+vwpDrRvmFgq4ghnCjkSXA2yGxaXxhYNSKOpMHPKimhdNCHkf5u/
X2gdQNwFBqfuaK/MBFK8Fl3vMq9VVTFgrIb+iKDVqCmGAdQnyrrOdI09QVtl1L/HXDAeV2MSGUjn
kWyhn0c75Uo+CEe1GUZD18L6uP1LVuciLXVsziAGa4IJ6StHinstdCxbLDurTxduy9tYKj+0RLvQ
4uK0yLkL3CTKKWnBWi0xL/32BuzK3NrsMHDGcH4z8koikj9FnZNwDW1jcbNdBz9baecnmableUVu
YN5XYhKFXd7NjGG7lDgNOD8UBoeDkGy2C5Hkk29CcrF8X+grbHnxMUcVIB5NCSDzCq5I7WcoRj9V
dBwlE33cxn5z/OMi+qK4jZpb1tbOUMhoj2v6XR3wakX1Px6wI9OuN7PLePDS6IiQLGzvgkGV00z2
xFaxuv/D1jmiuwAWMf3AQyL8tjehHrOE4J2V78F+nX87REUOWq2v5lWPb5/Xf7HsTvBFNLyDOsyB
1tJieBD5qEW/KUfJZwL73xs60PyZuq4X6SM1vLGXCj3s2JNHvBfBG+N2SNKupZh46s65yxSoopJS
eGc5LSp5CdE3hfLLTwqevBXMP/xTxFErWGMoafJv6hSeJWVZNx/An3oOa9FRfpjwuq7Ovqtu91EL
tSQ/uDUX2MAYAHS/lJlTtXTX+vgEqbnyq7WBLpidN8fyZbKTJZG9wtflCqBw5oXAMPE1x7r+00t+
JkVK5igmH+OLQI0B4E2DLHZleXvqPGasyDsw+Ao+SXSNTY6dPSUZgft9vYab4O1CdiYGEdgOyBMU
UviJ7MFb9pW5CBa88Ih12z5dRQ5+lC08qZpHSk8EES16w9Kfk4ThXGJPOcW0VgrfSV2ASQUSwhmK
Uy3fJUJH/dcE50omd8HeV6wndV6mmnSW28qy6lVMCcWL2rXbXvdlpqtOuNrDfq2F0dtn25xXc6Ok
wj1EyMCKIGh+lFRcxeCeeMGjzB1OKlZ5Y0EIueIdfZxfFSRZqP+Ku4S6MxebEyxLLfYOSUZUFFSB
jhfrMwERfVROjmX+EZXD6Fslkm1doFxJr1nHJPAlLg0exxupPDSglobPq42h00iKI86PjyCCbR/g
o/HC4wTWHfN9N2pDi+fY1PgdzxUy/34cM33x2UGFGgypHOJFQoHOAZTiT1vwsFZYelZ3XVjp7s5U
/pyiTwlqpB8jE2pLXcemykCHxZo++EMIzvDLYnyBoqXUq93LQ/X3D5kodm8F41+mfoaeYM24aKa1
NazuS5XsHwEo6X8p57v8B2Nnz/1Qf9Zu6GKnLHL74Jy+s43n5Ct4mhxOpoC25RhIb3kWTMW16OZR
o8k3guHldTy98yN60UorNLxYigX6oEsUlDDs2qCQWlgp9tmgRvu7L3NgMgnM1v3y95b4aAjeaN23
2T5PLaRvWjVPWQWw2jo/AmfdAXR8F3MLkGiCmqU0UelACBh05YwedLSbnMyqagmX2G6Bcc4dW97h
GEtaqHhh6LN0E+P1JfkIxSt7fLiMIH2ZoSE2rI4X6ilUUxw/jLjl0AWUZWb1qxlRJiYAwxERXR4E
CU+YYZUkh+07jDcp0pCwfzT1nfYg3LbZC/8zs4q2Q19zZ5OWyWdHwCyi2YgWO9k8KiBvfkHWRgtH
2F1KdSMUsNjMugpjqwhyyKr3XoBxdHIq408ad49eolLrQn7y5Iua7NMa8x7rMmNI56+pI0bPNF7l
jjJUaLBwjYxIYc3+AMwK6USjc7NH2nXNlV4xrk/6Q1VKbfMtIMjcLuQ7W5ivxBDKam82QjXVA/vD
i3bisqJIrvuJxFwA41CYmnA5UamDoklceYsXnDWj3g0h6a9udBZgHp2pRhXt5/4l/gcTPFNKSvxJ
C1zFbiFzqUaBhNT892HEDav9KOxNs9lYBqMi/PNQZYv81nEQ5EKI9bel5SCqbVb/imZIxWU9My7l
QD1lZEUB8Os+vj1RY9EAMSrvNvMMwnCF1BatoFlDhSKhVroN2G4oLqNHlbZ27rsLpfwf7auR1+LB
jKFBMftTjOG3I3BR4XP3OuO/uCOmmegBt67hh5LOMea7FPEWZhzLZXC6/lRKw14nBaRDfL/ef0MO
MXYOwxc/cxBOFzEpQmruDCR9RB8TCUXHAri03a3RluyIxqDSGCAuCKS5AS6K8g6HATQ9QTgimx+w
qPkRfWklxz9c9+lcUa0nbSkw/i7Ao7KfpGuQhSERJ5wb9szg2N3ZT8l1IVS3G0E5r646dENwzuI4
WjCLosW5XkGJc9yApThkjnV3Ovsn7b2vlPhnvTwAJ8eIHJabF+JlpU4qZ6YCvuvrwPEfO5qDaHpO
cPKfDCb8QPBOhN/mwmA6fEwK85aeEcuclWvTtU2jLZT7dc1NQx7nomrd1ZzJcZLOAtJCrLVGqZwk
MbYp4pLMXpPtC28g3ZZAPOMFXERQbteD+1TYCXKKe81kL3b65eYGQnhHQsQ8Jon9mr0usE0kG0oz
TjQWHjUQk+bnnkybMqJJax+rP58Gue3xE/aSY3zx2asE7HILT79NcYQ/Dq/Hmfhx0czCgnaIylOh
x2jwBT78FNQ96CBwsHA6qKCsJAUHJinCJvYbXeCvvMRcj9YuynIdO2lFyjTJLmegmEnx698zcR0n
NOTwxZz5cx820tH2nvknGpCwfbUw0J06oXZSL3o5LP6d8EmfhCZo+r3iChXAZIz1XH84WGHK7uP6
VMBjU3pDckTCjdBcfcGdDYHIq/3t6/VsRGYrWfc5Gv/yZQLm3DpLnNFWKW3glrc9dkSGkxJaohSj
ZSAJLAiQVqpnxusegrRJHX0JVIFXWuky5m+LywY3/gGhAK1deJ33/nyX6IEk1XsmcKt6Hfe9yWm+
NCcaQtX4jxsheavYjUa1Yr5Qj6K+opRmgxww39dRKpfLz2zbWbpKQmzhZe2vKi4lXsJ8fsP/Cr3B
zm7l2eTqDTU8hOPPu0/fBwp3FrBFfLooSBARyqfQVpfg8swuABgo3wGBUA73fVZWBLxCrn23xllp
Urm1tMJBZ9M1yW7ox12JQedXmhj6cFpM62LwpCmX0Mt1zkaep5W2O1CYo8McI2ioHi5VL3rQaoBj
OfJLD/FvPbzyBU3vjeieJ25myy7q6k8PfPZd/3oMlMIkFtZuxO98tXOG69/AYKNzC9faihhPsEI7
SRv73y3KvZQDilqueu39rraf0X6dlXCMmRK9W72uK81wpaNhkhQBIyI0dV9uXg1DyIsqpOPW67Qc
7nkMrkdb7oCbelhQNxWOfeXACzWu64lPkMc2cDXU47cIcm53qXgRU/nC6BXL+sgXgXeg063+mo2t
GKGORAmKEJbNb8GUJzyRBC/FCNcEbZngv87bhr5+ayun8TI5mvJZwANqS555HS28ayLqXXt7dBp7
saIBHxsURV0aDgNrw7tDetBSxl1JKtJ7v9Dvdiq/Oen4RwUQ18QvMhed/pFtoVMV6kE3KKpin41d
zb8l6GjFpw0v/LQ2IpcCOzmyZXNLmphHw7zvZZRGk+rLpcO/OJfTcNk9hMZ/aPadW1GEmJQ2HcUS
gdEMknxxprKEhddtpfYdQMznASAz6haHpFOj083oGUfa231MwQ2pCBH7dUsHwS5v+8F/GeB4yo1W
HU3h8Ro2byu+Zh5j0YozeBmGWTs7Bk4mg8O/JPMFG20u5Do5HZWg6UbbL/SMkpIFvxnUSNK2hVIf
1uDf5BwDYUXMsvKXGNsRRzC+ho/KDISC3iC9w1sZR6Kd+YuMxEBWVb5eYYye2spOB+Ly2ysAIO8k
ziE/S0+JsvtYUi5UpY7kKaAF7IXBXU5ViA76gteXyduWopMy0b76RjWTepOXlSc0maybCJa+jjx0
k/02KET2LjYZWnHIMU1gDl4xV8CJxCkdpNHfecNJBs+KCVosVxb5ZVlF/e0S5hAHajsIx66fyZBn
iunUFRFoe0YjGy4Xy1YC1bDm6U29OJQlfe4JdmZCZqrWq3RFxvmHQ0ueEXmHLDHg+XyhpquJHtdk
qT1l/R1WFvABGEFRviNzmcqvSOnN4qqahjQgXbr4rmbpzo0l7PCOJJSJu56yPULVivmcQYjdK0RC
Ml+Q+M4sC1xa6ILlYIx0OB8On/ngWsvSrs5NFVfcbfQ5nLZyeyl9bRnDezNORsCOIN49iLOeEr9E
+jxC9mkwXCWNfMyVaatBOtSHbbd1SVfYKXNl1euTlKmQlFYCOfY0J6pwOjFkSV1O5BsbO07ozO59
2D23qNAW5z08taaYAICK8jfql449vRgU7zkCSewKkiJnNa6+8S7TR5rvMBdcoqxS/W9Os+VCnsmU
KrPEB7KDVMIAlNl/0nXXQ9KDlOSyyW9OUYXxZanFRnwA60T6sYgRMiLE5ImqyXjKwqPFecNprbJ3
KemSCPCC07Wo3rUVOHmQdO5Mb6MmacO/R8gnFezP8FV7dIbDO9SpoI/DKSI2Cwh2Qk1ZhOPUF2qI
jqaPpQSR4P71NNT3KmZ+e9y34SNLpA3oMgXNQqdtPXkTZB94Lfw/SZcbjIpf4gYXyMNApZAvMTsQ
ZfVN4+Xsotq9RQ3O46pt4atLxccpaex721USMTzAqULUWHw7hi2IWr28T8X1GZN9z7E2pYEzgWS4
Gjw9Dl7pDfWCoBumqziALHmzv2IrPjTu5pH3wLmh2d2pSz0RLezBZFv/v1MbX7YL1PE7H5qrEznj
Ys0/2Gaqgr7Nb7BiYPQ++Oia5ma4K+pILZElxvvwpimKqRmTciu/+62JwWJ+sjRhQvz7aU7aRi5e
fFfcR+EwNDkox4fMj5EbP4V80euY5ubkWMN68dAtLvzW6z45Mza6RVs6NKsFweoClwnxpCvB5f+F
ZwKkHuKlzaVGnn36yagQ3XEPRkOwvbLw9uQoJWgEkzGZdO2L3LQtxoEbRv72VIfyKnMf1QNUD35M
uG9XGkvyCCxHksg9Jjj9P6O8MUW3da6/4kE2tyPFu57iUmU2sC9asQFXqrhEnK8psF+2Uuj8MrSA
rW7+2ReidM9cPhju4LjlYtFPqhyh38Vbki/mH8clfNM92MckglbU5+CiLl1GFVbPJQ93UjeAIx9v
Cnne0opWLk7ZvUfhFIDrqFZ0i7vnC1uHxJpqJegK42V95zDqWeU2G36iQEVVidaPkwUwPqYzhzWd
48OKRGlqDPwsfOx+TI89/zIDxU2OsLQcGHpXLAlYbXTU4bdv9RLXLM/WZcLyI7bF4afThDERZwg3
QHnc2XDdYwI5MbjXQeAHFzoBD417Ie96OliXp0IHe2jKo5Z5TESWOY4mWK3ncVpwPE1V7y4/8+Vl
G2X/Qug5jbmGfpHnv/Quhb1AxJ5tN2md9IS98jWJgKcgNawkZ1qw8Lo3mFucxDOimgDJhUiAkqIu
JZGUzmIc7sBmg1DrYD5Rxbjca+y6P3ibBS+WytKzO3OjXXWQFUo2NIR1+5UcyynshFgTqls66BCB
nhZSniMUtUOYAP9tqFN4msbqnFpWQ9OHciNG2YDy0AbrPx3W+Wo5qXnp5SluSrAzF9/5r7TLW7oy
4g2QCiPO+w2TeOMwqnmnFIxMQkXH24VNi2aXsWPKqI3q6FL3c53K2Mpddm0Hj9mYsE2rqMJloxG6
g1T9xuhqQNKSy8oEoDWhmFSGv4C9AbKMCOvASvTeYS+y2n8FDpk0Jwj/fuNSsY55I14Acsoa8ByQ
xsqSqyYizNO17ZNvcNz4MYhCGprE0OLYEmS5zzlLOuR9feuYwtCB2naYzlIN+Fto8kn3dIiOtSE1
RHa+SuOOuz2JTEhGMiiqGx0kbVSrKu7wU0BE/r9o6VFVzeh6tw9xSMIy8e0x+DTTFQLhQija2YrV
uNH4oPU5pbj1MpbyYg99I/6LN9qTbqi4EIXk3PZXg8kRXVokX/6f1St6SNAfNwz6AZVssROoif9b
gsjG1cDPYK3I0v3JfK2o3hK1rtIiT1HuZdq3yP7C5ZNhIZSmRUf9d9fJmgQT8HSCY6xOWdawyWFt
otJKu/+Q5iQTdGFZVEY+aeiQ2UKQXOEYvByds0CkwiTovKZJxWMu5oY7OHolYfKqH9pQwpEiAbN1
ML92nbPFHkgMVScDSCpSmtO0jwSUdfOgNs7t4JmCaEvuOftwDTkZXvF1yzNGeOtofZFG4Wemk654
xNl18ZHdkttpkkwCyKi0JimV1CN/Z05V5DDm5JzjgQ5C8ZOLDbksHRgo1ceu5Fl61b8YX+C1zi47
zJe8LaTBGysXGUfGGZ1keeuG226VO/J6XOsYcL8JPCw4k+T8zxSrJjuJoKkwzuGg0du/Or4zqgI8
B49uNltc6N3OVrKIzqkvhRkZ3ecIDVO7J60MzOQ7ZTrqslC/MqDU6D1GzKsrMdHG/lEIW1Pcvn5c
6YPUXb0trQG1aZ70ZaYTYH0AW2f/nnH0xSuZ2ACfY3L+HaSZg4jq0ekhgVl96LCSagll3Zc/VnQW
u2jkYwyLFdksWVcAjME/YHBApo89yE/KSIv9IGxE2WuWBWNR1yS6P3e8Lj4z/khLIqReWWEOuCqi
IptACvoq5kI2bchyZPypUaHS1g4d+HxZ5/OCSz+zELK8856YtFTK9Goy9JX3ev8QtU9n0EJKltOt
XPtth98+CNIt/oBeHiZ9IqxsWi1LOlgvrH1hiTKb9vEpI5BD9GEVfJu6wbBmO9uJgBRWXNXOB4sI
hynhBBCozaZlc/u7hLa4HmqMTWIaKHNPvWafFoHuEWC5s4jICscuPk4zJKvblJLmTDpL4bCH6aev
FxHSY+PzFSnYnp0F8hZjriHlpSAQuD3DkmA54ivQnNkCB9f0j6avClgzRV0xTCvXOQRXJms98eG4
Xqin1gVfM77vC80VicqBA0XfB6iC35NoWfi7jsthfXQhNfaBiL6uwSY5Qr1QGyP4WEEpDkIORNP7
nHRPfWh+DGw7BZ729uqQamEEmv4b+Kh7fL3n1kpCDnG5wHm8DJ6QqI5no/XCiMVr0dp5axO6WZWA
g6ZrN3w7Z85JM/ltfUzCF3VAjBGpIt/mB3qj4tI06QHG8wQu8mVxY8pLpXZdjss7Z1RSzovIDldz
fAwcvUwZOpRbb846xUljdBs+akpdHcrosfxsghEcMoBsdVM+x0M+D1xgFwRi+9AbZGO4Zw9eRr+/
20mHAQzSIhfloFL9N1ehohcCSpTDzEAMgU3dgytY7rtLE36CR4Ji4bygzB+YoEA/XrdIpvLDMcXM
jibJ4XGAoKZSMzDnWfj97rk4xR+17pX4XwCKoiSvXaXnIl56Vej//noHxJNZsZWaa7gQSgT7fOR7
HmytmszEfldUX9EQzBkzBLz9DvKfjf39TrL5vp6snNmponuKj549FSpm84QVDugZqaMm/u+6aHO+
XdphFz33y18ESd/X9c1P52WW9R59pXHAlrVpSyfh+BD5HvmpWv90pJ3ynUT3EHwTBoqhD3Q/bo0f
gZ8tpftAsCjJTZQWp+AbCTqk4ayiwwL3lDQt4OCebG5xGEBIpWiUQwgyIY+a9BA0UF8633WTeyij
MuRVdWJEZnXmOftvhfm1LgZ/AMtKLvRxQ7zvtw84op+9Cj2n5K4H9D3bahqnAb4PCVFkVolbH6Qv
vzJ8i12gW4C/lSvGiTkLpxzqMosjZZtELTfZyXAczY64nVt1+scPYdQEUuDPXAORdDKFAaL+8O77
J46b0c1l/6KHuceXBZN4iQrFLyly0FPess0tyP42+RWXhL6wXiTwXZeelikfojHMVyPqhZ5UpB4l
FW0epzIDVqtWjq91K1bZlnBVXUqLvQlPJj5+Oiy8ExPxere6kG3JCgQlwV8m1FFRpKaU6sUdtSHC
vk+8R+Yp0gHTpVSbyfpvx27d9wq2CgxRr9SCsMX/slhNv2ATT5cLjlUdg59K9WoPFIa6j5rhFx98
XvU9/yY8Sj8FcT+EE7opS4FfOdwAta4D08pVAOIT72HUqKR05O75D0xQSCznB38LT3L00O0Cn/KZ
nyzBTeMPbtfJiLVC3hDrN6UvX86YKNCFhlAlidO/QvgPCJzTnUvF7/5/oc20y6Iq1h0H6N3VdGBf
zbAvZRIIyJULj7n0YHEoDx5Yxgoox26rHf6H+sQrN0g+VEXIehM+CdTmwT8PN4kDl2wDwiEPprTO
HKd540StCVcdOEk2ZAGWmy5ZKZjSp2cM79YP5+Gre8/kRjALt8FwZr0Y1xKkZSlOmw593vABDXxw
34Pn/8KQLO6uF9S1fEh2q//OeGougkQzIDTXJhaRIFr9NFLp2MWyPokNTbQI2syp+n8UrCkvHOng
VHX9YN1u0jxcnPsi6S7uGjgYCszLtufe/QFny+I05Cf9n/dBaRybSAkKE+99ShtQS1MbDgmwbYB4
Wysgf5iB2P55LR6EHCXhp0drfqG6Wq+H92c7SGalV7Jei+LF+B7qlKwf2RD1fG4bphW2FSBNgZpK
DL9mPsYKe2hT2Tyts3GQ4ZQgUqOsXem9uZDFEa+pazHr6wDejkC6GGApB/XDoSs/PTSdUHKK50Yt
0m4C+XP3O/sIZbd2ficiu7UZ5lOZL/iyXQT7W/HImmYp9+5J5GnrpCIY1jY1K45Nu65gNRTfVhdh
HIFFEwN8aDYFZfq+ZApd58YPYrDSj2X+WMWZKaNyWLu3mczB5shPgP09hdRurgVQa3SEcwtEsHTM
T4fGq+ptp4cEms90PijH7MMBzc42AeVjgYz+pp+HvTx9Kag14Cih/W7pKDy619CTR84v8UNx6l9/
eD+JrqQlytenyLwCMXzGWhywI/LByqLyZ7TKsAtUhtS94ZZY9Sm+SDSMr4k9Smnzi9Y3O9I0VnJi
p+r8tq0vv0mmR9kFpv5tn4vtcB2nD3l3hw7IxUaknbWHnBwEOzvis5IhtWhD+EpGofWiyB/lEoEU
Hw52VS2tqh7VVBeRVgkSLHAGnLsX/ecYH+Ztt1HQCw/F9R76lZOAd0lw4KtqcU/Q3do4t48SZLbz
Or5DFZDZOmrBcSIcTjrS22sqsN2Ge2ioOJPUOZbhqtbK0KpjXPW3Hs4GQaECmS3TYa0AnGBpy9jM
6u1welhRdt4h3wQSMBrwC6MMArHEgf8WuOShbY53d2osTTO+Yqkn/yxgwCst5ZH5n4MqgLGz2GER
2iMIOQxTNlvZFgtSvCcpy/ljtE/E42VJ8ba2VFvWvA6TDRb0QdB1avhf3SgJa1dqSFWX/8bB4DrK
mB9TWFWbcf03Jhxr2V5eJKGr8gPvqVW9nrzqFmE0IFwYUumFnnF1PU71YH+lSkRc05cPtcsSgTWg
gPopvJlUP912qebGhN/Kpb1yNA16bx2YPSGjIVnLFiM3ruSCOsQWXkB9Oqj7DXGAOhMsiQ2oeDGN
br3oKsh1aUrI0N4keUiyibq8KmcVuei2cQDpM+Y2rmx1xqXppJ3Rgy3+Du6qwYIZA7d2oZnEGIbs
2J2m7jbhKevehVdPxn99InknggM6taf7UN0DGwHuQpr8t15VrqWNu8AncijASybLauF8gcpnR5vM
l7A6JHb7aApGTj3BoNiM+lABERTvgQEIU4BxKAeABd/9GRmUPkhoTJPhkaP2oMQXwDI/JLKJfyzd
0ZF4mBZbds+BG9YiXUwGIa1M14UB07VvCDmDUgHJJgXyqiyMDfLOPgloY/25Jwou1tjvmG/6WOcL
nKeMES4id35Q50nd5FdI5/vRqZrwhW771VRQX7++XGvW6Oio+hwQ3K9aq1R7doEV5hCQW3xi/Sxd
xLJwPlDyD782c4A9Yi3PYIZBCjXSovB4hf5YIxG4UqxJc2DK3PAX5K7pnRp2oMMv7T2HrR681SKd
lXyazPf07JIPMwHCgCutvCPXgSUGuV4o6qbunTY+GKwcxCkrKegm2E0yBc8pw0iR2YA2nvwgDApx
IANogbsVGS8xsAsQQr/29vPX5AMbs46Il5xHY57JWsIPT1xLDvCSeCURkYBvB0tLZTNHKL+U2l70
XuCsa0hgKSRQ/xhye9kQhyhMBK4cpeXI3F61UJTsyKYhLqlcQJJGvqjd1UoHDhWJDeKCQQsE8WT8
fVDuVuKX14ABlQBrvY6+w6Qque0EcHh6OFcZNL9PUCiJ6iuJzQ47VM1T0+xU6XCx/g0ThfIkCFZj
1NBdu3FgSWqN/j4yTDHRB/qilB1wM1vuAZJL9WE8ugFD039suBHrU9Wti4Lq/H3zwFn1nXRZeRTU
t3Q7r9N2ydGstfZkglsrnncyU5gMdOFAFMFvhb+MdyqsjdnXGGQKEgLBGRkqcmO3jbyybRlFLd2+
etjfHKEueruWOfwIPU22LefcLTReiA/V8IrF+n1IjJmFtqMloHfobqL6+KwgJcOhZ2y3g81onaWu
dfSuFWiVHLAHO6iW4fib2dsteZAbtRQz72Br98zS/eE0w8G7KEmaYUldVdXkeLNzygVPcenz5OUQ
RLzxrOdKvokOKcYizqVdldCp0PJzPLx5FxfGeyfECe/mFBvQMBkdb9DK7Vz0tSl9DQu9oPN14bZH
PfoXt8Qz+TM/zsmxjw/6kcwU16nZDFRzFuneT7IXmxtNwLxWvJPW2B8DqPd4z7D159fSpHvQPwKA
LRRvR1VCXtLe3hOsgebvQ64Iw3t6EmIbsUxn/ylXi4ipuqk2faZPdbOB13NhxUYsOoUVFdQ0lOLV
EJooTWdhdQhxinATbbaivO6E60wn1hJJaQ1aCkJcAdSA8XA+vsyqc6uoCryvGbtu70jK8h4o5lRi
8oyifix9Op8vAukcu9uq4FY2+Wx9uohAqFGuxfy/OFbXPSwmth9kC7NMHzu35zl2Q5sywb56ZmQz
M/eE4dGGTSQkBtWqejmDjjjqCtocJqMgz4P2UfI7C75ivo6jZX/u6wdJFvwqYY6yuBo4vwpDlX0Y
1SF+21mh3VUhRZwpMVWC3S/GzTSNAPw5h6h3qMHbzI0USvN3ebGoJc8fOro7XfY+oxAYDvyremrd
b1RPjx86E5EFyTh+Qf6uZWjWs30beXqpep8PbS6+L4erMKlqP2Njm+ezTWsG9yMurLKuBy+9v67n
sxHcBw9SpPjeq6jLwn4VoFgPEEovz/p1oUJK4venqZq0TtTJIJnlmospXT3u8K6XyoR5Vttlwn/8
saqBjVXZazNrQfh4+9qubvOS+j7/T5ne/GTe585vfMZwoX8fW8bBsu8d1uy9Zo9QjmpDljiHi2hr
pG5Q+2rWVdDguiMxxad+uEzl/hyHpaWxk3R7XrITHxQhl3mOauWuW5GO3Yj8jTwpxL/TFZLbpgDm
qXcA2/ZiqVK7muFc90Sh+YC56I63c3Kx7d8C8Jbnohm7ZrsZIojotimC/b3RpwTuoT8I/sgwNOsy
+vcNKEVHijuY39TlorL3a4nfzGrP7oHLNmeEPOfgeNCRDlk4qNH+NXKCYqdAc82kvnEjfi40EGXj
oZl7+IJlYj0MPlITUkUj5pcd+9Z+pvhwhbshPqh2CKiTc/+XfMnCeGWtc+yRt6yYI71nNj0KchE3
ZRV4Cf9eXyDmyz+iu3W7a4Lf6CQHL1SUF/FKXZC6z9DBz+/3ZD1HQ8/QLgMk8j5zHPj3+5bTlUkJ
XCMAvrjdrruCSght2PHDrvXjYyaa35ecw2N8ljytupsrrOheXSiVT555tjFhZFspKMOCJWHUdzFS
bDgpJP38xz7lFvCoCtHVMIO+LcHsttlPc+//xfJyOAzzekpd6Q3tkD74V+KKgV7Xb+OyNtp1sLGD
sARVks4YFlbl8kxZOivDgWoWY2qcYtY5BZ7kwiWhl+rxen+2QbB1AXj3W3dGxtktNN73CMkvCZGY
dJDFtRHifCP1w24FJgVr0Xsbn1rrvIfMnt1Hm74oZwPexXusyy1lBOVLqA/Wk7LDJ86Ap2yC+pv6
vEv4lVG5hoGaIuJOnUM0xZ1nddP2p3JCFN2ReevkUGYaSg0g4NiZHaNSA+n3Oz7XqURVAAmb/pkI
7K4ewSWRx3ZwgAfDcBcxwCc37lx9L2bRHyZ8YTxeRgrbcw2PEBgNxZ1OMb4Eszw5w68d0w2lk+Nt
iS5Ymv7yL86RMANHGGDazsigV2LCbAmlyreaxPPWU+6NzeUVkaptqYHRw/jHCeRAAsc5yQWvcGW8
P6LpoRZvKVNII68Y/+JqFU+Df1vDvKu/NWxNmZwtZmpP5dccmCZsVex3drag8AImKk4ZF0zPuYSj
hQsFpdnb/pwkyNtQCnJ7wcDIqLcdRxnYM9zUFGwzxwySmL3zX4CoSHs+hseVpcQL1tOIJpM4Vf92
OZ/MAM4zlv2LDkjXP7uC17odFlrbqOc0W4zpXQwU4nl7942nM/JaCjXIag7qJFXvP7xZLfFVUpHo
+XfB8Io1hPI7ydJf/EUOrqlTPxRH+6kXGKyUfaI3JIKsO/XKy0ut57Rfhg0M9E7ToNLYYThuaPe4
cIpqQJb7wAgM6OnzUvF7Xe2pxMRDMTFzxAwCEplFWhgerGiXQ3zzFPTXAhHbpJQ3hdkuWeyAjKff
+Wtl0iYmgdE6lxGBrJM+owxSN0Rm+fNMKeHu/PRnp6HwcMQ3B1gA3nf0cB9R1AjrJlpA+OonYtTh
/uNj+U0FXEDuRRMog1LdLlP+5k/HmR9ZXb4ZZGz0GR2cUXqKXm4UCUOGCzRUBhbUIb99BO8jZ+Ln
uG3FETkrlsZQlrkZy22gt7l/FYjIu1QYyMU5JFzdFAAo1VqAjXpIy9fmyD1fXUpChUUYsV6cle1n
xSU4nfh+1fDa59E/xqdbEL0BA/CVBK+qpUOaMKHI0fLznolTPwoSJyK/hfmh0BXncDVTEV5DcbdW
5m6QWJQwHKILv67p0fNoJKX/9xIBNtixAxOQKmNF0wqYS/ZTpNVJbmEMFRCW7keMVzqhZSVpe9L7
c5i7bjh8KgDp/Mazf5jD3rXMSqza9LLakmU3PNcjESnXPMEf7IRVKOceWK3XfazLp5yR2zLJ2Svg
bn/itDztAbdSmEl9fOZcjMJqGek3rxv6ZSqFcK+hD2gmtz8O+IE+UCkZ7qt9LmlhFqxxxmdDGurV
n68S6ow2FuVjJ6q02ai2IPHdeWn4TmRbceV0DQtqGvIImyJrEx2DMQlYJETB58oL2/N2I5SdJ5vw
TpyFfqU+lW3zQWHJXRGv1Vk+iuxG9rYw/Cf3oHb/G23s24cIvwPbQHJIQd2ayGmZwKLM+WsafyaS
RLDAPaYvzZS6mNUD4VjP/vIr917a1RL4JBd1L6zF69oTaHt0kMv7zweta6jBJcZ97GiresPoAtqQ
Ir931jQA7SFnmbDNl+3GIWlEGdGandQ/ypeSyuS0bCjHzwmG2Jo0sXWFIiHgFsYWJUWks7qbIxP7
d1LRMp+xqpi/cDom0OhKljoaodKTnO9AZIber1ly2jEYHEc9tdacnaiIJIuTOVi99yghAxuXfOGi
IYlekp6/poigw46L89cplv7jddSusC84/YTA4KLmeer62phzHGBZUfiYZcT4grjCUAiYWluo3mnS
KHqi6Xef6KODJQ4gAUjWvr66thgYQmXUZWnUwhnsZ461HrwDY/kHnsiz9V7nq0VAjKT6H8X9xcB0
6ETwGHVZA/FfnPye48aBx1UC8uCIvf+ktOQuTDSkIfxq9cHtmFGewf5FAvVRMnaKzY5dZZa2pi+t
EENtYgFLaXYd9Qai24zbj/YqxQrY3uUGXcs8zYuU5emAJd1C+4eQW5tCqQm/8jqiTh7mCQpK0tyF
8dRj3NSaYYdxOtCQsuruQ58/prg6ic/e2KoGaMnXB1MjFCD6GssanpFPEWR3dfVzP4/yNY5uDHTe
ctbk6n1kbIkjF4ZRB5qruRa+cfDXZktQCOEOK+NlT+iyFFCD+w1Xj6SGD56NFHyAFMavojC7dPn7
dPxcLV4DTYP9kN516TAMnDed7fIOdSKVEVlPRB5Lt+EbY9pn7ZhVqyBrDuaXrt2BMMsC0ZLnMTE4
6JEEFRWRcuSXSVfoT+QlYk1E2YG9D6QyHPjXgLFaSnV0EuXdMd6ypicFBHd3WrD2nbQAtrh79QPw
H/5CDfM+xpqgq8k2Zlq6IL4kIE081uKSbjD4gqZHoaMvzsdQlm55Eh1Olw6B5f1sM+tTSPyUrgJ6
LLmnGZ/iVkx9Jat9BMc2RUuydJNjjkWE907BkdjPhw3a5DvyldKl1lWv5W8uq4DhJWWeOtzfGkzg
YF6OGWw8PhQLMkSEREcc+/HwSjVgucdy5xqiv1lE6PggcFhdaj5l0ILWQOJRqlgsV2tziwGugEgD
yU50LdS4qRA6B93/wQajfWAg11JTrVuOf5+l7W6P87FcudnmMQ++srafp1G4hXYmGEWIT4xqMWpv
XfuriOLNXnFSptOC3uuSrnRNbK9TvinNdzQbAmYFchWywqU4LZzgWuY1sLitbvf64xMR3YbNOhWL
VjWNNDLvX8K76zLBMKp8RdQoJPQGfvVhntpDbnFwdmZXHHWFEwLdurLH4W8igGK+mkDWY1A/t4qA
KC/HT8xrjnGU6XK66gxVnh9VSob/LbRenCKBCjU0EnlxSiLvc7DO1hJKrSTeJ0GbzqcJBi7G8ZIl
W0/9vZ6ZWRP2bfPzuaqqNC4Rw/PX6Cu/ItmZdY0/PP6JYYGoa8cpSoyzONv9xrobYeMWIRTstf68
ejD45oc65WWj3q+Lmz1+o+jhzRYMAWlmXXlvyrLxNydySn5lkvpC1S7YZ0vLESwu+dLRw5o6mZ0C
Fgji6wpb/F3J7XW4QPZqix66qFfNYiTBBBQ/k4OOtlJj8THT0VqnDQ9y4axKT8crA3XBOV1ulsYZ
nt3dhJ/f1UmZRhp9VPNVYECaF1pLD1fnsq82pEYI/ccqcCJfQWkA5m1CQD7P7RVKkooA12Hw7p0F
Hx+PznKGzrZ6JTHYjr4MK1qQZ/FPp7Wf1YDzgCW4Ra0xZ/L/Z3ldmNUn2ubRGV16mQjI1wpKF1la
yc297OjsNR7MYXYC/2qaViWpdmE9xE2sW51uUpjjug1IS8ujHNDeW6Dkfkwn8xDiHYtubkJp56I3
+Fhj9vL9WhujRy4697upo3LZeCz6HJtAXYGu/Vn3gxUocRG0QQfqcSWfWtVczCke59AG3TiCk+pj
8dc/ITvjrnWxmOGsuYJnU/WcKcntrzLXqN0Z4Yw59becUeNZVmtnFA5XcvuQtRxJneO5roWIk9aS
Hl67u7cYiDIIC3iGfwVgxVbqyL9Xqms1BeDmr91eyPxcbG7SqYDQYOLr8OzucqvpKXMO2BiPMoVd
Ob5/LPLIl/gpNvt+dS6R2iUO6Ry2PZUJ1MiMYtSnT73payMKnlvl61YbwDdYjAIzDqLGWkLDu2DU
QTrqizu4NfuKqsbmX166sLBOEDmgnPmnROmuknWtS+bz7xDb8Tx3fcm8BxqIe9XKxHrCI55MQIVn
CVvb1eoBvWVpXvr2xKttPb/1zGXzfX1Owv32lL714ModZ9PgoBXVKZh2j6kvV0q5OxBLGOsRxbrE
+Q8AcFmWrUpJFNNqyrFr49KCtkBvTSZgP90ICVgA+vhQgnW0244O2xa+kznkiBuhMxBJg5t7W9e8
6qWGDHhSLol9FM/syoB3zjhxM3wWcCe0Rnwo9OHqAgdQKeAWo+UIXSB3c+q8eiMB3rtCDiLrC6XN
422YcHW03C+oVCua19sLE0rPRVkq9EDeuBNQAg+Npd7Nwqa4cFoPyJziT9Vba+AjeonRA9cdyb7g
BCngebM3BuygQPflTu9mxQML7TLQ8ky+HgKU6lwFu+E0VBMSJiy6Pr5sotR52JFdO7otkaVtmycD
rAtvznHYKa8+jRcnBPjmgcuQCI4qunubhSQ/xIEYsS90iBwcLnjZviz+jaBINhC0HqAOSgT7mrAb
dUSz2NIUDJ7fMkjQz4XuiduGj/tmEsIr5Eb8tbcnOlXfweqbvL488R9dHfHfBNBReoYZiVZvteZY
qKNx/oPvMW0scSXOhoInrcNl8amYZ00Krv+K0RVGGNcU1Ee5keYbrmQS2kCczFVGKcwmzRUZd+yk
KRdu150oTWT4P8hIS5/y7TrnRu2kLbHbYTFbrdbhYUt8RtmSEQ1BFXtvjIYUfLoRqchjdMCyw5Un
1sb0yXGNt8cvFUIoPMKcL55ceM0eoz6zP2A9k+gnFbGI7PKU1tKblH7Lg1yRdW4XAciH4Bx05c4E
y6nS9KMCQQNuyRUmcD8Lh2/XJgqFiQ8PRS17XrnTF+3bVKEkGbO1O026ME2n1w2C9O2YU4pn9URB
Jz0SALdgzlVdLYEcOGpaivEp7rHf78wDaTZaJjlyHLuWO9vvAjanMu9vlG/2FegKiSxTwjRdi+SD
VDJ5FOe458z0U9mSGQUVaFjzVflorW0GEQpwS7S9v17KQDYpeNN8YR3czQZV4swnvAZyVJ8LmW3C
X6xeao7rn+Urf5vQmhWuMxTdM4h5f/u+dz0Ltv/dYIf2ptsowVH/3T0TRKeGzZ5wtdnkbVcjwtct
n/AE530nxX1QgJwNb7XfVbuG1fwedcCB+D7fC/5PoNdANxeYvxP4YtbtC3Cxl2guD6u+pk4O68dL
qqQIQXNPkL4dFLi4C+r7tWbgLt2LSGF2+SKYS/xfi6uNzv0y0jV8O8JHagN19olLSuDzNVo7iK99
Q2DbTLtJhgYAl5SmJQ+ZNmtDdANW/IdwXvv6gMUzRzJW4ZFQqNEaaZs7/Qbsqmys3E3acF466GEq
2G23DxqyJXLJdcR1I6NpSbzuZxbUqrTBKVSqHlxyNAbkmCp+KEh/qx/HesyZOZAmv5xlLZJmnaqy
qR6fC5qsyZt8lhp2qzyq4lKZGODDZX5lSfTMRVN7nt304yNaV7mUarDy+c7vzer4WdHjl4COk9rm
eUppI7ENYuNu2CjI2zPOme4PoGk736a/85p0qUcVppVeLxF+sfzDjyFYoURyYqiRfAZdejSA91Xu
HU5jyK+d4K02St6rbwDOxCPKSMahxikdbx73RyoiQAVeU3rGVIj29bKqvXx6uxukS0U73cJzmeET
Xwm6ktaddUAvUIO4QdTMh+RqMfQZWpZZSPdoVQYEATP/ZqYNK3GrXpyJW3xVlNS5AW8Yi7D9LKNj
mn7WRw3FXj91dycwzO7QIG+8RwEj9iDBmCS74BcXhvyMfrhcLeuh8EJMjBo27xwGoNjQ11GNnsmV
YXPYwQHvsn7i5vO01DI6fEXR5izCNLV/2l3CNEIZTBPgkr1cxFEO63FJ+ip9wA/Wfd+ZI+2865Cf
baSVtharC0ANmHrTdphq/HCLVnWSNEA7EZFlE6DpIYvT+sJCnlMBjJUGnY3zghr0/YSkjQECmbNe
dBrWyqa8HLLnXIiFElfuzxLkkbYxbUAWOJSvdutr9oW4riADE758RYo8UfZ+Kh0XThP6ng6bVUDu
bsJnja4LVzz2pD/bNtVjxujWGXovPNQpLQ0d0PW3kha3bzGj6XkJkj/XINXxNVO9izFBoqkFyIGc
QYffGtWoPqPlDAlMkAgjdT4wkwf9wnRFnc9MPxJp6F59ZQPsPQ+qrYvKVK7SZwDIl/j9STkEVZv+
TsiUSDSYclbHYkxjNTFzZGWOrCZe0pPD57oHAvQrvFaF/8zxtwjc+FKLN4PEZEI+CG2q8w+QhO3Z
ufXljjeTWcRspBr8WTOBaQWZSintSSISNrqPJDID2KjBcniYcgfJVf58OohdnSliCMETotbgCkGg
0tuM+FelNVy6Y4BXGso41U5RyMpD27B7zKCA5vcUFMk3MjAiKsIu0C6i1o2FfJH6PD+bWRLiBzdh
Pn0sWtbmhEvnfVsyKgfxG1lowrC0HhijSXdd5aNaJbD0OlSPc0GGbkKCKugwNSJfvWinoOlN0SNc
LOAZbNeL6jqJsZ7drJqfYcZ5vvtpzpSnJBuzI5nohwM7hMQA6DzDngP1jTleUKASF8H7k0EAjTje
+dX+63nSEIYylFcYGh7CQVK9dbLug8ClWOWis9wsulFWOp0WyKav1dBOyqhFOGLFDMCyQa4ra+du
HKankYgCpGCLz+KRyisfH9f6TTNbVvPtQVZpqmR/F99Tjq1jqi9r8LNY4znmfeI/Zovj6eEX1km/
udUiNTujKl70PnxSfgNjZvRK7yqoiv/85aM57jnJXufCT/pv7NdXrdqzUTGvUytnR/Rt2TaRsTUw
1NWhcaLYGr/wpY+On02rW56/HXoGI+AzmFzgr/qgMAuX9rKFM1P5GrsjdbXaDBA/8ON1a68JNtVc
/CdmQ050aoXLQWiOnIgZ1FGP0KG7XCumWS1Ac3mp9EjYyWM6qraoDp/IzO7yFGSseO4WsxrrbyQH
/WI26Umfy/99R5O+ARyJUAMqbLTuEjNE18CwsxESZbso3sUOzE0pkLeFte6GQJQQvdncYqBWYq1L
yrgNJhdf8+kVXZXLqOETrZ6Oab4iNkL2R3TFV5jENCfXytpLLO1rUSxqAyOPo4cheFb88KMD+Obv
Y07WrkBf3p1LESc9gVLSe6MC5txQigxLgb0zAN8hnV0WFYnq0SMh8v9Cy3q3a49CeGxjzs7d1FgQ
RM7RXW3SQ/sBN0Qyff+GEhP5UCkz7en9j/Dhziv3q1F4lBKaQLGfTSRis2CHmRLCUpiOEw55YYEL
o+VNRepnjg6rGyLH9mBQ3taVZ2YU5dn2Zsz7zdWR1Vt6aqmcIiofhKAKTnHDfqVsUB2urX7L2AST
oSEfVWa+j9EOXV4736MMHz4T3qjq1LUlewJkWJgWD129UiG7hd7g3ITbAhd79MDjKYF2FOtisCGp
g3pQZDO05ebfFhARpU+B8Q67ADEH8ZS6/9BZSuGFHRVx0eoUh2nkF/jRT8m4+AMoxDcZuoOEHhcQ
b69Kp6slp/OH+NWVI0fpx8ZO3sTepXoCX8MZuIRvS4yQ+6PiwqAKFBur9oZfGx0cMhYCn517fAj9
xSpqvkhHcwFk53v3fuVcqWKoTSW68LZLm6XZvfAbJOjztuVepnQd49Tm8trzVUjPtVkgWHjY8mP+
yglTeyxLCXDmqFs93Yr0a4Kcw/BIAm3bFut1RpF3V3py0EQW17lqZJJaJM+i0x4AMysX0hWQQJUM
9S0ub9Tmhy+jlrZQ8PcoeAGHvBSlqahxyEzK77z2OcWRCabvetJqxtq6Vje66fNScdY+6Py8N48h
+ebZbDbsyF8ETQIM7VpJ8v8NjH9fVG9MD+lGdSSEU/Tdvd3uY+TjO0X6KV1Io7I0SdPy+Avqe4ib
eTO8KH1zOZc/WHyeeA534ezOxUF3OYeNkHXpYSX3F7RG/+fxU23cjUfOO0GDV9KnQRjxxyaK8kh4
zx9fIQEcW/FFK3ZR0as45yLoi0iMPlrgjinYgu82kDa6pfEp7l4DbcV2FFw00blkd/jsGEnM/oBd
Q+bKN+rs8+rJjrnYl+P7Nrs8woE0nsPLY0X4bXfF7LNtG4LYU6U/rQEPCnsp1oHCQLyqFXMfxkXh
njRO9QceKzp0UgmutoCGoXqj/sw7F+xGRwjgoOOXEKooCAYXRtkziHau+Ja5F2/ka72RgZAcGGTk
4l4UKFqGF+jiOdZchzQ+w7/jEbb7itcWZjEYFnOhe2CSkoqIPJpzjToTnyEcN7t+ZatBCkdzf3eW
p5kZzFlvE29IPn5Q8lrcVaoK9oqRjsn96y1emFOPR16F87mkmSZV0k1qGY8zjtNmjm6JP6OrJXfO
C9mdn4BrWp8LJCCcVUH5wHplJJRL84gB4A4Vpi8BFiYwIeDORSsNaGDpl0tZA9ROLPn9GH/V1xRL
h3ROThVEY/uYkamsnuIbQMr367DZL7i9Ibv9j60hPr5noPCT7SYb2tOy9ZLD0unuSQ90t7/yU/w9
oicOrbIWB5UA1vtCP7qbYOiaV09pmuQWIeD8niVQ5JVV/jx+FeBvdoi+zZBNFQrrEakjkktzLHtr
NcMNutYwyfJ0y1QvOb/HRUVPptjRKjY2VdbL8A1VbfyMjNCUi8qh29n73JTSgwjJw8dCP5rnPP6g
+rp2wngyxdgYzDGI4y+i8lx0zBsj1DiDuPyqSCCfcy3vHswvl0CbZh3oHk7I9Iq8T1/BT0VgJGO/
Rj/zfQN8j9LUGwSpP/RT8aAvRvAsQq8TfK/uxnQs3y4DoWxe89lclfjRvM9vd+8O0jG61jZOhQot
cT+WjYnKyU68BJ+dI3PgEDlVcnFVmza4saYvtr6EHCU5S4sZORx0Slni+R39yQfVJ4L3waFzHzB7
mEY0awD0Xv91VGuxN4xxASjoSmeK+xeR4Rf9DxTtJaEJ0iGr64GLb7aX+EekeIdaQ5TkUvoPBTqz
Mu1k3eIRQwLtn4ctNIwpjKwLu8RGN3Bp/g8/fzCa2GWjGmAAiD69fZq+Eq4RaohV4BNVtmw1KaSF
ObY5CkqxFQgZtSX+B6f9jnND06W6+6jx1Dn7XrDF6e/Ced4yn01GWNuQMa79MwQOKuGsataIVPFt
QWkBx1PsmI4SpY+uDN9VK1Y7v/Jd0aJRD2Z9Aa28T7HGCkiAH+aIZ3pZgiDPBiI5rVWQXFmZWG+2
q7//nsOAaHTgbOls/AQj1GNWlQdZYoZkrhHmvibHtwQd7XVhKY/QWz2PzTvouRXwGKaLdvWNHZba
PD75JMyK9CYYQLwnOsFJVQl/xM4spXkcoPp4tKMg3jbsiWEqWN8wVpPZmDXWq2QbykomyyvWNgRm
LJEd+X0OwClbELjMmCLqV25sYLQLI6/iiwbFIS6fWUBh4BjWjNtCTIbZYhzSH+zn8XF8EteIfTPS
qwaoIhvTOSoyNutvouhwPkDpC8lnRuFvAO3x56Q4VXPjHgWHMszSVqoC1PtDIhfrwPtuNEO+YyFf
7k4hsjR5bMJphk3CmpnmKwVYg+0IjccW87mXZIfmjHseWrQ2ZCusJjxQ0UDw3s3yolvB9fPTotgt
139/eDa/2QsVMhgG6hEVET6zGfC+OJpI679BeTjIUIVyHukYfn3DiIeHaCmSJSygQqDx9lU2UxpK
g4T1IDJJ6vwCWVpudAV1kmbNgkss323u2XA8Sp4NPCES2bRYhLS3Do6Kq8728olPJYDCICInLEY4
vv/idn1cm8jt0qlxRT94IydS1j20E8ELzUNGXVmO80xaYzPWC4lklDuEBQpjcE1qyvboBH6Y7M/m
5AFXbKg+EvJxcNQXhD6ZYaDl6eLfWrSa7OXHDOU+BjNyIpCkzi7lwVhSNcBn1nDxH0vYGmTLtiOH
a2BwAybxI0mlFXxbWknZewtSWjZ4p29kUQAAVUCE9krfznjrDIRlUAaTSy5YIWqQlXL2+ylB5yvW
m44TzdDR7yVumEbEXEDqWpuG1p7RqaU6YRXIRzsHZm4ymdSFANpTIAuzh+28UleX67nUP30Psdjo
oCVDNv31mkkdyroZAz0+Io4hNyIqhTRjctPjhtLk6Z1tYWRcS+mdaH4T1UykuCIQ3nEgTj6Tsx4d
mRrfnMBLlXnciJrcXyg/s5vT6vXOeCwuBVB9a3ecglWx37SIwUoOFvDJucjTKOUa++xh8nAoBRqS
HMfroFzMa100mtnIArr8latF0pOYGGztELRpkGJZxaguQpwRrSwPdUVlkKAC/5gJxsVHdq/WCaNn
a5DKZqdyHNej+ypCUgYlo1X41i7TQhrlOrr7LUpQJtNT1ZLgpj6PR4baNjogblsn/wkvLCfwDI2H
H2QmuCf+GoePqRar15knOxtXOTSe/3elPcx1vhtSWHn0oP0lN2ubOf1vgbYJ8oQYugAP76Pigwo7
1kww7b0kOKY5Kr9cTZj/39tmB7zBPV/n7yxa5ZgyEw/K1hxMPP3bnqc4QBQRzF86uhG1DSbDrqWH
RBD5Zfb4Lfl74PVlN64544jnPyccMX8N4b0490SZtmyqLkLnR8YixUntigsBIgOHL3DTGX3rL0AK
CAEzvh66rU3psfamWUwMniHt1fe8b+d1sL1P1yR4P6/K54tT7wc62yM+mqXbsvKkdsMMnnfYDtUt
SovPsbB5isEhREuqs7hcwuPjdq4JdNRvPoM6qjdSq0u39gSg9BVWEu1JQn6OBnCzXqUmy16tj+yq
BUKLzKvL6QSw0bY25n/VU7mMWRNpr3ZUjkP/uONelLv5HwMEQA76O+cVH1xJzUsCVp+ccqtUFCH7
XmWgAP37BpYq+Z4C/3aBGI+QOVr4sJOQNSUV8SuSe6TKXJ/6NxvEUXe587LYtoOADVAO/sS5tymq
OWWuUgeK5zik8kzm/oJuC77P3q0JBXj7TLRgadetLUMzsYP05mCcriqWhc1tymlCPw8g3o0Qtejl
wrg0SRtbAYugcTDm2mE8Z0fvDvkdhc9MwZ/v5ctVEIO3KZ5SeqNzED6+c8Acr3WR5b0aJ/B7YZkT
WoCQhV0ZhcLGVIRSJXl5cwfQp5kbJPODbxntjOBlhr7QHVv71VFfCTHPHZss4J9b16xTwlnsNp+/
cnfRdL7NEq6FPRB5vwUoz6+KC7GTbJ5opffEMkr2BxXCWPcLgFg+CQQEoBX04vw75qSblKUndpJi
wKbZyNx7TDsDUhl0+f4UE4363x+PIEXO4C+1G8Tw2GFZqVjJx77NPVEubs33H/9sai62/TVXx5dg
F3QSptzomiSQJ+PWePd6s3LFkGT7rQsU1p5V9ifdltYLhAGWSRJwPK5/057JmQV9cE1Rd/QLAydK
cwxAEvzvhYW5yJmuJ/JLCUwGNdlR1aTVgMh19rgHLnUinmoprrms/saQN30+ZHotaJ7EgfG5oo2K
KZK/uj5lO0HaB+jDCpWpQBF9i3VOrZCp3HtWtKNDefENS8ouV9vPO0siLwSOzrAVDaph3/r2ll+A
9tX7jpRCaJgKj5A1pgqE8N7SJuRTcB1TjlEq69wrMWqD6mLMHmvAgICUNYAD5+worQfNvLvY29uM
/lMXu7lmuBfqZtyMHyslnp3TjVGDnXL6NNR7OXjLn0BUJHICleFOArTJXwJCy/7KliUw7t2GFNit
kPOuIsUTMGulSpzx0Q/L0n+jvW+NRE/xwiw2ULDt50/u/ITGt46au9i74On1Q+QwoAAFqs/WXjNE
shVJnEbQxCmdRKQLm+ePzyXbqhYqOjWx9C5uot20XS848DuPFBa9ACy5axIzx8DqGRiYr86Vl0TR
a8HcBxth0QSSCQD6XTgZIp9irZSKpzrHJdY4j9u06pMmNcw09l23u/3vSNE28R4jmvdOYJUbjkjj
vEiurywW2QQT7aoLg8GQrKMFdIgy/0VDZ+yYXTPrVA4moVPnenSj9I67fGuGUCZsbQCpLeD5Ctb5
iX5bvIJMo+hwqtae0L9u3Ykb2rifuM/w4mMF42wXZJmEQzxDwaxZSQbdQ8bod8hHvirQZPzs+Fzl
6CotkJVGt/ajLLojEK8QZnw9NZ7c3xy0wVBMAKHInHfNaKScSk0IepImg0vr+TNEum1MmSxuPgNI
O2T/gSlSE6r56Ar8i59EmIaHVlYYTkXI19wTZ+hOfRyMOByCytiTz0UCk1cm5/ZjyEZ2kpGlWiwt
YIEZUBc2XUhn6NsCdWjn5d6CVsFemLNRFvB7FKf2zON2Kh6tLcXBVgahTidSfrCUsRMU/sADTEWU
4PRb+4nz+XWq1BEMhDRSvRAMitLGwm+R8dGDXSypNpTC/PDab/vZPMWsHvacxYgpt8z/x9uNEZQt
d/aHaKJu4RnAFF3MLyEFtIPUgDxuO8dQ0eEl8QHtWDavUfI7tBaIXFubRH9kSEfZqLIwS3DOaPZK
p5+yMRoAPGqWdt+UjMD7HOwxGqaFqjCe1S5daHtJZ4Zrn39I6YgAa31Fx95O3rgtTo++t0CyuY4X
Fb1icx/oYbdTW8NLW5ZQS0ffhc3+SHEHvSHw6uXjjEiQ3iJV6yMNGspIzHnTv+AOHX1qE/RP/vO6
gZAIg5VYstBvtZWPSH65zvw9+sk4BnhIs8pmmlXROO/wHmUFtqr8zKjMsmIsPvtI741Siew7z7Hu
V9T9s4UBWnn/snGzIgC7kCRl9bUAwSV7ffgp99FhdjlYSpX9qurnMSqEyyJDJl4B0aP1Zs0D1amO
O3DvxGfpiPNibdOX7yh4exWTdelmt8MbLv8Fa4YTLNv6qaCUiZ7JKQbctjXQv1K4BzCxwB0NG42i
PdLtRgc2XHMXLyrmHoW3muVai8pYa0GvRKTGJo4FrpdpsQ2BIrGkkTsOVf0VjgAOVkdFt6IoI+dO
K6RYB6F4fMaa4lFmhrw08ThkW2DdlsepGyhGT4m00ZF0LHMeHORqxFJMFypdvvD15CecEIQQXgE5
eJN/Oxr1iSaePwd9H/Ym2KAREZajvEnShbYR+zUQIo9YULC3J3GDeSTN7Tj0c0hDGh11bbHGnhv/
q9St+xS4GW9mRJKo/bGmkmLNFqpZVLOSTET00DV1URgMAYXAJLlieeviWbilb+Dx+r6EhIK4FmOx
nh6acAdtvdToGHHQgEN9eEoGgKqFBG+e3wAsoE1gY8D/qVmZijT6I27yCRkLr4XLNdvYLh0uN5gp
Nzh1F7ikbXA3A0dbBULoO+dwFF3wScFS6FiuqvxGUZGmJqLZ6LUuR/OKE+LgAspiNB0Mso8Xu56c
8+TovGDUCZPNUsmyXus2jL2gSOII+8ZZ5s7gqcCALxXgweZWLgXqOrHQmvdZBSocuk0/X8F3o01x
twyIBoC04maa0ACTgKQJbVwmpsVugW5+F+VvwhEES3n0GAmbR/Y/TIyVJuf+1YELmZWjrb1wXHo2
HKswqcIPFqUc6RNS5QpNPnbDLXiTzE6Kx9tfY57YYozXUaBRxE1hYZ9SARi1WYsi358RKy2FENaJ
jMJhKio2ViBpBANTwUsa4suwe+iTuN3TaY4en14wl6YYtDg3ESur9PJ47rO2Tf5ebU0PjabKBrM1
IrRCf4IsMWpIHkdJFP6gvnf4sgpcvBi1G6QvZItYptgMUZbF/Bs0loA8i+cbNjMW4AOtzC9CzEpB
EF+UqSqMTDX5utXsHK7N1fOSrVrzHZ7p0UUWwg4oA6qJG7OEf7ncn5cFN0lf+CetylqLEtliRqYL
2X16ZWpvLQdHr3O0QGJYsJ0VvMwkXypVwUfP5jX0cLnFjyjXmRuL02VurVENizdRR6Npse6gkR4W
Y4gqiOrRm9gg2HzCgwa3q4H8OCRL+HrSh0yXslbbeNMV4mL51FHZrRREVItCLyuwNzkgydpXqNpN
I5hO4wNvkG33DMFE8TGCTAoCbmHerVjH9E9JH53lspuAOPXnO1NgBTTCgpZxErDV0k0s2mThR4gA
DTVqe0x42Mu2/NPdVisYTQYpwaKop/oXwYV3viSsFglI26pvanSA9/tjlMWkvEy4e0tbjjycjZ11
do9kBJmFoiagSqrUbeWdsfmZXoSK/ZBjt2Xz/Ny1ndA0sHFZOqUySppfDhnWhQHyf7mnGs7Q5Dw8
TTFudFMN27/bLLfXRc1rBOyFznlx1Pht+H594KKnNlg/9/E6P0K+auwgLrh1fJnHuw6oraixHnzI
em2Th2d4p38hW3S3E4sPNJUO5jrTTQ03twVW9f1iKor+7XX7ckK7OVThqwKr97ITSyh7fwvN3ZZM
xj1MAXEW/pXhTp71Z3NDFFbL8JQzfCNPpJo64P8oWnfExzy1OLOjAJQZP4mqWuPyxDK2rdkslZnY
AMLmkH/FVLtAW5vIEWCy1LNXSu+f2nq1fQFXqS0m+z3YpTwcD974f4DPsh7+1iRNHv3Q/qd7K90T
l7TQATNjayUJmkHeP3U7CHnPYZz8vbA4KbbWWm2Sw4VjLGC/JoYP/uLfanZpJ8OqC+cW53zroC+d
FYPCk6fr/yVdapDMi8Kij8KfhjoQ9sn7CDsg+P6tbk7riDd2UkLOz5Unmjd0IdxXJBAr5oJq7R33
km0zPzvbOpbvxiMkl2KQ6esPGP05h1SuFTZNzk1XgUcYVuJrvYlT5ISNK/iuKKg8WTc+WdYkNOHO
gi9UNhU0QFC/U9Ao1W6JRcKKKJoJjdIZfengTbjjhrh26KE+tDIusjgbIO9mQsbW18igEJD/yJmd
qiUnZTrX5X0zuLjTMRf0xc66eGw9KmFtAG/5OMlPHZV2Pneh8edG+cyZSESfPMNsvvpL3uwiZWaX
cv1CDcVa2VY0Y8J30hiPpBK58M7IT4VjHZqK5qN3BBv79Z++vOhcVr2vSHc0WDaKCdOGWjMZ1JJz
053SkVR7XHKrITFBkZ4egfUjlbJbgrTiQf8avF1Xtc3a7o4NcMEdZWxgydPXUxPcYmhz4iV+CrOF
eFNIhhREVUmQxJZVJ/s846w8N3z2/XffW4cLpL0OsdWGHehJsmhqhm0rzoNckNiQ4xYvwOsk7V1Q
0QWN+xZOrHr+MNCsvMarDfU6KmwnYbEKmFH4g3hd6V9xinbGdi/nDy0IaAC1bF7DUvZPZDsfRTbE
aQpKNuaG1NdKSNz3ArutIVHArNwuWonMNNSLpFPbpy8Atyarq0Qyf6OZ69IU1yy4gATdH07PCF2D
J5Gqwh6NATQpQE0vSisbwtgghrvzwQR2+tk+qG5ImVaa0bycomOntutol11zFvX1V8cKj7e52H+o
60tw2B5OE22Lt3phvcF8mAUKwsPI9WGOsCLJPWn7J0I4duy8iCZTWsAhoIfG81HhdtGvjpr/unQI
NlcBd+GmUhlbD1Faaa0tA6O037yInQIWyjRGe5De/qSO7Bt/2Z0rTDdQMIYm+vjSSCCxa7qfCZLU
3xKwmZ2c/Xq4Ggy1GuA+z4zo7WoEKpXXlS+kwl/7dG4JX6xGg7XCEuLcK14oOeKV05J9hSBN7maB
g3JwF0aGjMg5LqGxYpzEOAm8lV0qPuOPxee6Lru07T+DbizVNwF69xsAmVOpEXjnfFnw7bIrNmUq
8hhoCpfizOCniznKAD8158h2K0R+K6mv2IzsmiSFN5Lh0l8ncwstrs+yu1XwXaAgnWjiUmczWFBa
hbdwtjSIa0BpYL4DcDKwPxnCcoZL2NEUMyJeUjrbHT2nvhBl8Yd2kRcoaeg0qQPwmYb43awMzR/u
cA3yFBk+Lf+EeQWQmxhYggLRteyU4oEtL6R3NyyshxW6qjX/y89qK8nxYv+JjUSiwgVaUDzYXDAq
MlyiamTf1lPSVL6oowULVNl0NYl67B42ZPZsMNE8CffRQZ7P8sG8gsSMMBg/daCTewRbuofuY5Yc
YauRdettsiyiijcvgvVqdDB+SzFUNe9USy8/s1YhVEmppMlho7CtReYJJdSDaXL4b8WZIjDypEji
zPhvr2R24JMzNjDw+NY7O+Sx8Zy/IGfQVooAVdpGwphJy/73KysjJvOhw2lgXu/sdeSMaCdgaP35
XkRXBVY6fiXeT/d5bxMPUV0GFC4MUxfhlpss0eswJkYljO/BrAL/pmyLvTHcCviIItN72a3P8C+3
ypPAgCaNoLTTy8wOQkkSRnCj7NFWVtaIEJ7Rsk45S+LGPHLEFVl8EwFNa6kHyAPOlYkpyYHiHafy
QzAqHNB9AEpBWwAyyT8QFgkZXMkzrStgfJOP5YZqWqC1xkQXlZdxwG3z4cmFDwP3nerQen2xB7tf
jK1RoyuJL2eIYwobreOUjUaUvs8CIC0NKFcWwm7g20tKSmntLTo2MyqbYqXVKxm/J2hut3Xxg0Tv
qdmsf+ucq5EY2bFB8O26229BLJT420a3IVHAiLrBeGVdfVpLnUXNVP18iN0yxXNvuFiP027XYrQM
q7t7lONrqC/jE4ZNMN2auPQMhGO6K7i4vjQsmL4BYd4M+8ozhRjZw9BJ38q+U4+HUpiZCOB4TTDp
kFB6oODZ17OCS36O4n3JBOIGUDY3l6cVtP4n2EN3Eq3R7Tbze9i7OnBkiAWbF5bsauAtrEt/njze
x1PiJUxkXMuzcAlgDRa7OdAl0SyC8gbF1b9Ta+no4pRxN1M2y3t2yOrwBi+mGPgaPl8Bo6+w3xUg
3iIKpxGCAOIHmtgg984dzqHGHDI66xAAhmVx+ETyNTaW/iboO/y0V2C3Yv7BkIk6dpscf//jjNC0
uNzt/zXR8woFVbG+sWIrhwKPMRPlKavpi8bGFZbRRZwtLbzfoW08vUiH4L2nbnFz+AghyXTB2CMg
2REEC4t7vshjgaVEx3yMWFf4cYzbd33HApuUYNRzrtxUp+wiDfCXwEOzlKFQ/mucT9nfU42ODvNx
vohB6hTp9xueqiqt3/AD83UD7Mn68jwn6D4mFTby9or3wwpFBwYd4C4ZbYW2DEmVyS1ip41GHKLS
Jg6XhId7fmPKZDUPLAWzANG7W/vbmTPIjZzg4UN1ndZ9OFdt/xpY+U/PPkwHtDpVQCj9BgRR4tJE
8oLbB1b6BUco0gqRu9I0FfGnq8kuiSRHIAUzCOpZNdMpDcgumYWmyGzyWekuo1cBphuBNqRd6n8s
YN/HeqA8yTLKxXhxzkagNR8pgrWMTTDyJxBBo/LDMhfOgUP0ZuVeLf8oqITvJfpfZfrReafsOQtN
XlVX5WlUvfi2wMkwuSPkQfk2xhT7PKUms5+x9P6Y8OM9tuiowLuNwCTkMB77DUFpRlWoyL/NPZKn
FVIkMLYlgVRvC8QJNgDXZ0DYVF62RyXFo1uk2JUgNZikw/hB/HDbPUx77/YIKCfn9grxg3W+93fe
BVZVhhgTV7N3YVh06m9uKaArLpog7R23hzDlHVnzP/wkvq07mIqDcKhVP6Z5SJoqJ1KSUbCbsGCT
mg9TNMNBiljvWC45GroE5dOGiOXkv6vNG8JaJPg+8vncZF+hO+kULmll3QUzZ8i2wx3ywn8N320a
9Gm9QUTkhYnKyDOnxA2fn5eirJ86LbbC9yWRUelBmzejBCsh8lUCVN8dSxHK7h4rSgCW+ji7hlgn
kzpgtHqTC2lP7MMHnkAZcOctQY75jXpSH0/bl0vwffMbKJB1Xz64P5l0v/HDX5D5kbvcgifJ95pD
AAK8nAPGqb9KvVkmWPqL5jA2LWsWV+lw7GgrHc1AJhntUGo0tBpRSqjuzYazM0Ml8jQQVWqkUCkG
v8b3GKGfgl2IdQIyVbGoGl4GduWkgR7CNENLn5Mztw+uGVpsMSq2O0Euq1++XGpIBdCvo1AB5NEN
uYYjtjh80aBSMJMF7tFMukLCn/GB+74lU1mGV36llktqsSIGoSOmSmlpmc+J4XsZAXIpDxHtSTlP
K8+RfMjxXwT7b1iKJ/bjvd13aC3lulQbAv+3iYH0dWxmMyBps9WQ7TXRLakkSJqsXMjiMXUQcg8o
w2KA3aOvxXNYPghmPS75Fj4UQGCVxjBf12ULzUc654PsA5bk68ey3XhjmO717rBaBV+EewlyrfwW
0i4x+h4qrJina48R9nCOLVy/J1zf2MIUInonGlPtJm2tevCgfoUT3WfnceVQFa8CH2boL48+/Xpi
QaEKM0StzZXSFP55CglI3nV0McRo93cSlA7exY89wuiaWQ3XnA+tVeIDB4m9vDJXKO/Mun2N5sun
A/xjLoOrJZNR+ajykKQQ+CEdExQtZKKuu//ur0ScNIymqXhNFWT5MAjdBTqW5CtpiVYQO+m/26t/
1EgEEbjeyFHMwcDs7h4WM89z8VBPxtQgJhZC76tBrf1Dxmu8thPkx3BCQ3eDEl0YHQYE20py2gs3
iJDBwmsyiPPVtEyInFgdfUOiLRj1rRmqtovYged6UkH+DujEBjyyhUIe38TzJXKzdR0ptsw7GiRE
W8kFsSTmSUPkOhR6FE/2/DYU5e97fJ8O5ak0akZKGuS80YRB6Wt6AjOnh45XbiIQw8bVlP/UfIe7
zJ5mpWqyBUwPgxsCzHBGfrZEgf0CCcPTfaSHuc/BQsl9V/+7fDTZWr3t/W7esAOSV8dWDYS5ZBe0
A9a6fFpw5SeOPqW+hwc/5QJ7fGLMmn1QaIFLCro9E4Mk+Mq+Du6KTuXc6MgKF5a0rpOKk/hJZ5yT
06h1+XTaSrgB55Jq9NBunQXPgY/nv+tHYNHOy2Y72JH5d/SqmUJ63l2haewKo/qAmZSgqEQAxDJW
ulRY9NZQ2ztf7A7TEtGcoWhFCKeBo8DsuXOWC1hbauT/EyVqMEKd5CgxJ+rhlWMxOCvXUaIe2158
EFYePhi19uAe7tVEe8oQ1eIOc0Az8YapMzpXBUHNVLMv2ca26FCpU9FxSGA1bTgJl9+WNilFZWjR
6/WblWgUa4SwjDvaCv8YxbxsTtxH11GmULIMWRrAbQfyAkTUgGWx1S1/02Q4ggH8DDMls0vDL6rL
IJ6nys8Jic42nj0caAzWrHkM2ruX1dX6BxZx66H/N1P4gEm79zqeIMX4GzzHGZUVHl3PLlJyJJwl
PdDAZAW4LF44OsGsrUqz0E6asn3tOHM8VWqFyRompkk3uLAPXjDbaBniwCSvK3rcqSCbEi2o0t0D
E6Y9hl06l+xS8RzaSOTWBdUuiPNOaVVlPnTJjpzRgdPlhQi8PXAGLniXTMglQHy93nVdAYC+pJFK
0loPoHwI4W7runn6yQs5k7YGajNhgn4QHr2EY5zUHdGVMW9bq4tRAJSlp3W+56gSWns6uTDXKho9
7PdHRdRwYhS8pl1o6LAghUGpPm/AGCzCVlCoZoKK/jMwP+OdQSftkMZ4v52W2zMujlrTY6fulIDE
OSTo0WLwuClFDtmoA5RgXjEbO51rftX4ZXmQrYrnS+0xe8svl7v26qFxepEKK1DTOxNFJLIlkAQr
Ya/ztLJFE4EjuhFZPMWo9daLiNbdd/K45SKHCEI2IzVvlxux6CYW6iwJ24zfpoWCaiKAeFPyJtGX
4fD1wR5dHlMbJDJU9QFie9wp2rKpymB1847SVkMBijI91nf6r5PzHcIf0L8mPazqnTTWfg+8yWAR
GchO0e0GTSrkcdb6/UpVMGwIt4BVJud6MWNNQ0tlemGZrAmUjecuS4hNJG8aMZDEhvQuJfs6U6to
2zeu+miaWRasN65cYE2hiXLrwizkaGUlc1gAFhi6ZC3JP55PiW6cVM4R23da6xUpDt8t3NjlyXR3
Jg9Y7+pOiUNL+lto+7snl2NdMS3p83+PoWZ5bwIxKhozjY+pzbMLOw7LGMVf6wrc5NXOhYCT7w/j
FPv3d/RtL/u0Np4e8f7jxsLlGwmL5+YPbUNuPkBpFa06FqcFuJ7NU7Wmfhbn/lKughInEKCtvj5P
3Iafv5dIX7JVZ+kyVo5I7uXr1JRzUX4QicimvGMDeH3q4ZaWzpFI/eN9pxv+wTjZgNaOUGPSsPDv
BR3Rq59MY4W5sM9LYnF9lJ477Mz7YOG8PvKZ/siC4NJB1MMIUaJ9C+2p4YFfjID16qBglJKA3zqA
K1vvMfYojQwt82U+romhpMICKzN4LKTiAHAI5oqXKUOvv/WLwjaxur3Yu1WPezst2YEmZx0xnf1r
t+EUgZN3B2HYDfWI3I4zABQoT08I8YRaldEdj97HkSndMapARNuJ2UeRYLdVDf75Q0oJQ9DQdArX
7XxnSLOL5+EtXv/R4CRXVQEgluyHDkkIbDsivF6ihVB0PAfvx7lxuLFNfde1AYG+6jhG6rgLrFzc
lEp1U5Si/AehqCTXw8xo1oZRY0Fur3kyjTKiamoZvfS1MvwiE7A3W7yqETxU6rhD9svFr3fQzlDU
2O6iXUoImJEKm5YCV6ekM2UJfaAFFQxmUPQ9kPmNU7SXq27K3tUm3xKZU6yNEupsLWPUzm6tDH0p
YUKhthj9s8l2cx4wCWGhwqBcdXEH45szfL+ZPV9c2GNJy71l+gqUgGyg4/aFYxykq4L2jZVAJCbm
k5SMg+MxH9TXOWG0BNIQiq8LtzFj7R0PuYGGEpzU0gOHH45L+kmBqyK84gGyn049xo9ayMsCAPBa
+78R1wp3H/2U+k/AC6lHC5ScrNDsRyfaqTizRySBFjIC9XP0zU7YZd+em9HN73fzjc74HADnXL3D
VZXwLD5AVAnh/GANB8XdNHM5jO0wER4j/4cGK/0HM78V9AXAVljI/34g+it+Ha2C+BUSXsrWas+3
JcBfwQk/inbTFg2JjOb/uG12kwE/LsyC+3dPaY2C1MW7AwTCu2dj7fbtkh6BhLUUxFvEfxGIXBMp
Tn3Hfn13XFiC43DcaIb+pRFJ29qx9JAqOKzXLGDc4r3/kNwo9LdSaBq9OnFryw10JhQCNykN69/N
+xe+MP9xjUoEu8d2apEiDbfLpFZomWw4I5UdlLvHuan4x1WnerTSZdTPvMI5onDvxbtZgKD7LPyG
1fk6AVAV6vS3gn8q9EbjQc/Fgzp0CD+/avDWZzlJSOEEUZ06o+iAO2YT9UcNTfX7ujEp0GzYRQXW
IXagS/lSxk1TLE0tHdyDJ/r/aCwnLjFNSu+hnvvLmlXMTyz1MuOsbBcJMvR/Z1YsitS2FlBMce/q
RLx/BU6+jlLYdcTjpSxmnkxH0VvstNFkoXmA1kc8WnIrAHvIvIAkT/qdyLLUBi7mG/Xm+/4fy/na
kg1o/idhzqywW4t5efncVpyR4JvGBcGlCUuXTexw0JiEeXGUqtRKDy1prdhj7xbwekxF+nzvccCL
DXwzLONcoQG9bITJb48h5T59lslsuOMSjP29kT+Nq2ymn14rDHT267xT8/tOhODqyngx+DQLzfik
SOlBcw0YIMApnbghllTP8zXxacWm7hc2KI6aSXr4aDJ/QDLiBuGvMfCKAoGcWZX0UBeqW4pGialZ
WjqOdy9q/kq+yzSNirPgUlENMYYQJgcMl+iO4wWnIcp/X9NXQYrW+9MVQT4bHN4JG/Nq/IkoQGrY
u/1iT6ttzqu9qTC+B035xNrGKhJ458CRbfg77C47AjFdMR1gKvBDDk5IJFGq9278GWKVMv8xUIAr
L8f56hFYgc56uZbedNCsvCbe7hBWpDVQ2vZz+BoU70vKFgZKqhJXxFdDMWKratuY12m/iOTsmAJD
VZkNwxkpthOHdm730P1iw3L786eyspAXslnBmt+TOEZ/gSkJoqkG9NNd5YWKzMVSY0CvCXfsM3yB
r0osQgJ6z6+PDL59oMVooPRbUqEfomzrJZDekDff5EOMWSYLL/u5R1Q2kRL6IA3LjnLtPfOD7qXx
MYYg2OEAErAX/ZKaVwQ6kPRvzzjJt0cqIejGx+obOUMkmiCYy+IajMkCggWXQW7hwo0XHlVRMNkl
ebcg1/hYtRE/Fhdxu7eU0CxZfOVEjOKBtYRIjjD93Yb5iO7T3HhQ+Biqww6VkCDW1xua7+jXIhF8
Nk3Gk/OcMTPTWIohu0yA3pPYITJ6pQc9vJXz9QmQ/1NYOYgLAELOFQFHQOe+snBziyRYRwfO/MrX
dDIhPd7KZAn2bdsxQWJPZ2EsD0f+fEyqu5lkiAxe7Fea7H8q8QSs/XNTvjhAi+nxgoda+srz/Oai
LsJEsglvGEfdtpNzL8S1EYe0ClxYJYM4+iXhzKElIWGR0o+fJFUUBwjKSPoeJXQdvIp/AG8A61Nh
Ars0UmwFSiosiqvqqIT8/HGKnIN9p0JER/3lXJYd9qF2+1rGAmhlgNsBUMQmaG8UFZXHFUqh1Mxj
nYEGNutPcWiqkv+ir90rKb+GA2yoawa9wKE/RuY+E0+jXBPinGcl7q4zX4rf2DYBRlDFhcxgnNPz
e0MEdhcrBAQT9hVXAyp9NMmfIl5Q5JNTnZ6uSH9c1Cv4lADEeVv/YOk8MhgSHMoCaJwqxnoGi7yQ
rwehm1GXrT/7wFQ7qiVRMzI2q1SncT8lIJROF4VWVB4LqqKVh7j9RTbKgv7AgIuZS9CFOk2O8193
K/c/r2I5OkdhPw8uu+8fEdCcRTbEby2ApnZPoyEump3RekFpPXXQqen2G1mnlr8ryJGtXaqu+Lim
9lJqImNDiR/g4PCtAihLuUdsk1Zi5+1dWjpISKiiB215F+ADNItskgLdrv8o4rggJxCIXVS0qmTd
ol9n0YOihXEj1widG+qs416eR08Q++A/CpArPUr5n/ADbOUX8Wg3OxUjD7114oRVDCPUaVxwsWha
hkNS89tDkmsObgiO4LFV3FaxxbarZ9TARmCfWutuZB33Xp8ubqxBZoLnJ9Sg2rq3gXLscn7YuSpU
3Cyh/6P68/++AVPbrmnWH+YKhaPEgseAgu4w8nLgCL/jedpvkLsknV74ZW6F35U7E7NnQwaEOiB1
Z8/gwryGU3xgKPGJOBukKD7JAJU+gYb7QUpibc5MyZhBIqFrdM3zCqyKz9yXdGR7VeD3Xn4Dvnvh
005n9dQsEghvBC/91LVmfCpC74pIPq75gw9dLKaSCHjSk8S7xQ7f3958kgj8PUua5FiPhW8auaVW
1+e4+jpOatCOojIyZWdiw8FJue4pJxtiDdwE1cvUEJDHo/Gj7QTTTeGXNvnCLuj8wm7C/9gUGGKc
mHyTz6tOFmm52hV0P5vdIAPCCgtMFCeLoQ3v2x+A8h/l/VijhvBCFe5mHIO7pXO1ChwfpdBf07n5
y1ocdLo+xSMkcDyUqYIuwILnEyt9u+K95o9rwckRorKkQ4Rfn+ANW9JM56M5D5MtxtfNpOG6q/QW
wfPNvVLJaqgWnwCHG8skMYepAUZty7qTED69rFEqJrqdPAvGNTFiSFzPeYi+6T5SCmgvG3yy0ZcM
zOWG+7yFTQ/TutFjFhGDMS5wyF8vshyqfZfuNM8BJv3Z5yXeY88JE+/ekO+7oOcZ98ZXbhhKwXKL
ZkiJ81GYm4g2QDF8eqOvgkagu0Z+wchsfy35rYE9M/GKqlXWPz1xvQT2MOIUNyeb55ep89LDEfZE
APUq+BlTdAcoVClbC2ZHPauKXaFpsquTF49GZfHYMTIO6cBPuEq9Ppy7nkLMvv0o/MG7E4CZKih4
Ou2uNCMeFZTB0mOwLSrS+cLNhggsG7nTuk6CILtvGY9YGMd5VjpQEJG1YhsBHy0v6j7Z6Ae6bUqF
PfDPAkZig2OQcK3GSrVmq8Dcr/m+RRykZ9LFQbtSqcGdv2D+4sBjUWYyhGi3eBiAdTtrN3eEFJUt
WTKEHHSzAMh2EqRavRHcTAfp672V8b0zH6592h/YtOfxRgLmSm4ANHDYGEGEO03s5LKTPNyLGEaq
+O+BaocUQs9uoZzpf4It/BFl8Z6X6sdmDEkPz9a0N6KMPrZDxnY6IxRHJq7BXMrZDOrCODP72U3q
XRiX9Kc3y0+t64IjiTN2Tfy5AXPiTcVTweVGxEbIj5R+irigTfMmeQdrturtBnKLhCauCfzlOBq9
G9sAJ7wQ10TYIxjZeyOgFlnehMOjxxIrs0IGw5nKsQQiyL1+cA0HDsnQdfrNddX6rGkXdG5yxhzm
YDf6mrAUp1zxJ6uDFb+QE7bK4yu3ZdiRGDxOqSraPKgZyjC7D9VPjNl8lIvcoNUy5Gl++M/ezgDV
3BtUo4OnkV1Xi41i2VlVpmhohD/5IUErZ0e3bt7RYoxmLzgjBa3b1bD10pjDkC9M8h/Nj05vmsTA
37h7s3JSiwdwc2E0tHzxa3Sn9NOK4lx6TJelJJVsdd6r7dbOGsvCFmsy5DCK2ev04e0ihqQDMAuI
lOor0BcOTvdPbtLGO+gJ1piyk06zK0MmkBI0MYz2kmA8MdTSdsPwwcz8Enm1DPYLbtrxnMdCrbRb
ZsGuPNk647PtEPh/ROTtT/Rn83mPWg50udLvcQDJLDhsAosaFS6cfocKensRvKcBRMLv+dvWIZty
EoXKTfpDvWiT0dI1/dkpxH8KrxzrZbi3zOv2gueD8rhf3q8uTFENh1m9NFik8GSP/hkGajCsgp/V
hiagVOmovrWsmwhp5/xxSb3jwaXbgefwj3mAzJd+rUDMw66XbSot96cmSxz9UJQlXClOhG5ucKdU
4jgAChyyNncBnMvheKjsezGgiAkfY0ecLxCJdA1BpY6K/AuHDH1PDMTS999DrC3V7C+XsyipE14Y
GEMpUD0Hr8at6O+GYyMON9HwRV1KO9PgOasblli1RhSy9D7iWwq0tSoM0fVUREKTUXhA4XFh95lJ
kjRkAvgJ4E7/FnbLmReWVcIh7ZNqiUbFXVQ0IwzU4VT37hwCozYshACbQTKv6dT9gCgAzcj4M9Ns
2hUs2kkMBMdbDpuoEZ1uHBarmhGNGrxhPwziADumLR6xhdT9GC+uW/nFc35Q+U9M5ds/11I/g7pP
2TGAIu2OOoXH5ug9IW9O6c7NOkGbgYbC8B6gIaKZ1acFO+bYw8FjMH64OmMMYedq+VZip2BtpiCs
rJkrXiKBx/FaT/iMRC7kuy2TvRHIxGmPOL/BoUpxwOLBdPmLXp1dR8MolM3D2w/g3brwxlUZLD4/
MiHaJvy+FI7Asl4R96GksML3n123N0FxMRD6nZAp7vKEtQPKxnWVNhpkWHvaG1uFccc+Pu2LULRl
fZ6qr3Lr0eHa6ecZaYkmCyZN+A6wSdMdXVrnEESiEr/hiVjB5A62HNSeQTI9TjCn4pVJXcU0TY9s
HzrC1e0sbhHJ0N4wXxCLjijy6Lr5eVxrN95mZOYpZhFLz6ryGdlukS5w+AZZUf02JB2x34kPsJ1N
55ykvZZFsufc4sohvl4rgABZwPEDh21fwXInoQz/ZmB16LiLIHbg6VTyVWNv6yfRzCo09POmjWEc
WSSbJG5ULwxBC0CI8ZQ90dIzGY1iB2uI25AxSz/3VrtlP6bl9zJPptmVbQ8895SlZpN+pmlVkTs0
VixYFVfpUY8e9nOnyxTsRLQi644SR7w6uzhX/qWgIGhTHn1+oL20PUYajLzVOhl8i/i3sQNBYNZj
F5g31Ie4wcWcO7BdpJb/WVguv6i3ev1Cc9R6++jZUZMRs1aeIlShqMghxFQ43N++x2bQjRtnXm0T
JDgZ/38h1NZd77LBa5NoEAg8rjJgsO1jZIHqnbM4OmMDT5UUttjP4qiGaxHapGiI0M4eh4ENzLG7
GTJSOqEF1+6y7Nfpx9Zm8CWWECu3ip1EXAsrzKf/9+YvkrF4npP1SxmMMT4bGBLqLlB/FkDXASZu
IwmJXGzEL9XAST698PD0Qni267oD/7fPCMN+MWkOtTXBRvEA49ml8T5YomQtuDFEL+n8+LchgPmU
Mxx9w1ZzsraZhA/pa/gzAB11RgYVw7u8WT2iMuzCt4B7Amh62S64k15xVYVCz8RkdO2sSM4Bie8i
YKYC/WXW2D89W4RFQ6On8bkyOWPYv/PjbEgJctLMBk9KW4G9nKpYT4ORinhUIwwdudSvWyiHkMaT
iZvcSZqRJQEJhblQuN+VVOrDJ9klMR9kh414xIpfr5XpR09wb/ZVCLy3zzF4oyAHXyXS0SGlx6fM
O6vGaQSz+cOgqSNrOrvOz/VE0YrwF+8Fh1GQtmiYkdWJHNdRDxxk240qFe/ltbo2+nUKCF9a8+Kg
+8KGA769RlhcRuYJyqHfa1UGJ+lyHdNx54jHOYwQiJuUf6M1pYWahwgBjRCv7ymzrUTb4eG86MlV
VtCCOMpFtCrl93IIgSAynBxJcHUmu37GlIpZM/GqRzZNO3D7NbWl16iph5GUzeMG9+0DgsMFWA1B
vlKCknt5KSHVtYnS+ioG4FmizRqHo9LLKuCBjJF34cgRIq5Hc7mfrSZBr0t5F0tfo8sigy6Xqf9W
alhHQ6ihJD/Dg1NgV2g5CX689Q7G1CqcQykMn9VSjgn5Lp1jrdn2Jk0mfsW6QyMCfXbOuGW/XoAb
OLGvYVjZ/3i8ffzzwCShHQeZtaCJuu7PfIV1DwqFg3udIgSx/prIDN7enJr+t5OrmT94fSdVBgcp
thdfRBD+qo0UFTn0iglVb/6gMNW3qzm4Pon+tyPKIbJt6CsDQNqwUX12Edb8x/m8xVNxVzVts6mE
FriZ0+EuStsXIxOD5h+T4AwJZfTDFkDZ8ApvhAsfx8L0Pq8R0UkzQPy5q2UuQR8QV44wFCVEttZ8
RWkv968MJgYo1d8jhr/+jz5HNyOWdoxZEYK+dVvburLhy07b+qz9PQWw9FeVenI4wDb3l1ShjrFP
xihH8oMrDxf+HSdKusyy4a+xdAqV6PFicz5ypDgD4lwuEhIc4L/IPBHQzlIGMI83HYp68Mnb8RDi
ajpF9Jo6fjB1Bzt25bEdANqlFAjKFQ1/Xr5+5z/kg7uo4W2K1TeDIZD7MIuACy1PqriGilU075ab
97/hVOaT/Fy+tVJRLx919MLXU1WGKVlVIMKCpgMlcnfqTs2bbdsGPuHPYX1fYYDLLDNNE19DqQ9g
Yd1fgewGNXTAsXmcn6UPmAX+6QiQXYCTkmmoPP1H5ijNmZ/CwlFhjgaI0Hk+uClBpIdY4k6nN7Uj
q3xfnTuiYqA+BlFw6T2B9gqWQwPGQPnCEFo7538Ljkfhl7UwSO1f5Rsdv17gc9Gp9E9d0Z9BmcHV
GD6ovnJRTm0dI0EbSYJi7YGUfcftOseXIP4ZRYtODLEKq0MQz3H23hliJu4a2Iqld+I6UKOX7siZ
MI/8IxvNh7Bf+RLEBxFZATd1FfpI6A3a57xRQH0gvvBPd3ezvmmAoScO/ZQ60gSYFay32a2Wi5bM
bCow5FCVIj9POC+S/eINfdfFDAfkUCpHd22Ke4aCdJ/EdHL0hUqAUsDnjXkuPWqBWMrtGB/jobSE
47TffnIPRv8tyEvq3qO+Wbme4xhr8H3ZCjIJlzrE44EdxTHBnBkZEhYvd9si7EWKlvvxGUxIiW4U
ESM6/HNGfb8xPxyWNQd6jK3Cm0iA/Mn9vSVn9fy+T2GpBpv7HmNAkKoTACjGcDjvv+BndPPY8z8H
UrRTEXZ3n6CwI+NnwCrcA8WJ/XTpiPsQy6ccRBm5sHpfAfw+s/OPCf/WWVGIzQEKRSNhhuaHGxtd
yMMbYsziNhwyZDclncS79U8S1celWx2NDojtxs9ZCix+TQJ9eoMJ1aPAmjt4MfnK39Va7ABWz1cI
HB8e1RGIKc1QLrkuJaVqvtmdIWGC48bcsXq2GcXFl2aPLGIBQLdjUZdz9EPUEf68xqCk64yLGMKY
X/NoIe7R6CAicvLfAiSdoXL+h9BBbTTXEE2NTcCTfnx8/sXwpzHRFSwsP46zz50Ras7Ny1GzLevI
+vdyYZyBT+cSLlMwCatZb49mJpnEIrE/WXtajexWo5A+qq/j9/EiuqHAv61ayUBOWRE1s/qoXqYC
Sd7kppMfJu/DfjoGT5tQUCr6qnIk9WjOSI4+djwaAytAtw1Fuf7p5gsssVRxMsQbe08+gbkvHhLm
WXQd+ab3jjroF1kZoZ3hMrZaPy/Zadij+omeDhT4/BISxVvx/EM181eX8JAiG9CfJxPYDkJ85H8q
xE6aWm8+lMV+BaXzOpQlX+3HDJqAfzvhBc2570HmWzzA1ZaCpSGiagRQVTxGIHFG6xxhpYs4ndlC
cYR/IMD1WIzcGA0yHwY6ZwE8q3OeLfG78Yrek/u6lucbSMc3/MRdrdXcxz1S+uXvNh78uTO0kDKd
heeJLzBgQJWxnyuKHCCswpVhkcI/9wN/ZVcnM7lK4sWS0kLc/veMyZuS8fwIm/Xmv4RpEeZUabG1
oRone2C15wQItyBOy9YXbfvXdQtBp0ZC0YWI2IAdmaIVH15VbOMT46Soqvwp19BKO2eDBZEyvfs3
RkQ+awUNpKxoRxQ5goMfK/2mWrBnLNBizfaEOpp3a1G42Pu2RE0cqDPrLibVfG7yK5KQW2XSadFB
3rp8UJYTEjyhzONuQveekpLW3TbWkhlHdJY+FAAtywRmS68iQsiwTC5fYGIltiw4RWyCNI+KKUOo
RKGU5ik0DVI7PoxeRtfEh3RrWA1i6ZuLd0xXSzjdJo3Ivx5KDKLPUNYsuWCyWFmdvY6JoiofycF3
BzuCZLvAIhxQ0Drf0mBWtCDbip+dX0EXbJpedbFHgQpqTBFiPLgTWKipuvuGPr9PLRoU4EngDmTc
zDjtUSOHd3173widyv3YnPOoxu6pAI/Ton4z4XvwD7x9oTgfiRbQ+9k51kaRSBlT1gqg3Gd2klfZ
mbb8GVmtuB8fu3HpRYbIwqUdsH3p6sOSjU7vA5XQgGJzpNkSoyOoxA7q91QX8OeEgj3h7xfBbvM5
OXxhGQRb+mCJyZgPRp5C7NbgLDR6a8yyvrpObusjdrzVhP2vZ/0IaGdM6ZgVbsRYoDWjoi7jts0Q
AqKnzxTHcLEUTfYQ6mdOztea4Tcpu0Y3Ve8TOEvrdpzJjjlP0yRQSUijjlLBXHyZ/kxuoAQWcibc
TA9o8jrFm2QiM43Eluu3/X6XsXYjaf+qbUBHnFNwGHwW20uusu8+qXhjRN1q/M6rkY/l0Hm++Ygu
iCE6Y291C/fMdZmeWcUx1ThHwNy2w0ID3BwSoaD7Fx9irrn0SNt8R2K+Ila1lAfqZJkAYHjHuMSR
UC+j0+/DJhy8l8PPX1AGvlolQHmDxS7uUWqr/hJTnTuP7L3a8PN/6JphH01u5UNvCi3y+gieDMi5
Z7t2RIWzjGjIdo6CcdJd4lHg88V8KCFMbq9mbVeY40kTGXDDhRYbWedYHqMzukMQs4PmK7tLrTs+
XMC0G3EwPpyWCfrO5RDoeYy/I9QEeNFWE+jxF6riqT/A0d9h2XU4pCgJIRe5VBm31ALR8RfkEegW
ykbjL4DEj6Gbs7dpy9jqSFar8erkipL3HmHVHdgPeeDu70VYjTP82yaoxDO2uCKsLqCg/012ZOQE
dnB8mj9Dmk4Rnti4K+qhYEhB5a2S6IeGaE4WanMNEcZz+N/x9ODcPkeTBM6N2mXrWOFfpLwspDNx
HQJkTHQNMI8Q1b3MylryBq8PFY4+SBcCSadxUWtd8f3ZDXZR53s9RGA16s3f6RpT5CxGMIHcIQZp
CJFfxDw37hqv0DCaBD6YEuZijIE2XtwJT+7RRcCClcJ0LBcbGwhD0FbT3mwTKn+5fgPWyEMY7hfv
COr6RwQpYNPE+zW7XfrlPb2vFPyISKw/QdUPYyfGFdkxXbMpuglzPhRlwYE7/ggKMBR6bg59p9pe
4FEJEjjJRXcY2Oh1jehE1WUah3IuaHdS47HzUPGtE4B5AlNlM2EntwWqcokNFYqnrFbcsSrPyOYf
SliX24zmqEIT9Y6XrUlcjBlPLlOMMbMYHqaneyOSYqaccImxLB5cKehozWRQiglE0fsiOlD3Dj3Z
Mb0r9wznvXzta7e7lKA1Fck9tGEbKqRRxJpT6Hp0BJ9Qrkw9/WRnPU8/Sdh2LZOsPdq5+kK3FvRo
jQ1j0GklUtL3lv0Cc1IgMi24mpG0UuvFgp1TW6vHWkTQkgRSVqZjc8ppCQbBIqCTuKWgc0+8KWzf
SODN7s7MoYz4VN3FD2GvriBDsLwz1iD+PlKzmXfRBdvvoATTq6Ej2qMH0/B8eMJYrtASscBcMY3w
9UHRHjaA/khbOlxpcXhjjYPT1qdoJnGFQPSTuyQf99OrrFaZpf+aj4QTASffiN7Nh0C5zoiwk/G+
7ExbFPFZq2QTKLfm1b835WWMnuOHcQEVtj3lh4bqX3GhZpMw5gnz91t3qGMoKCZdH15b8M1Kl846
dTGNbYuerNsh2iZ21UIXTEcfRVMS7rJJexpa/GEMtR3qBrZw9PkWuehEec7lJOg1OT7K8M/Yu/4P
Ci+/reAxhyriRehPuKn0+6PrirwvBO1X2W/hcIJj5w1BcLrOfVNAfa6pHz7V5MjQn4qPYXGXO0Z9
poU2ZCLL1njPl7cvnUm/WKkfg8xBSd1SzUkpImQjwF7W3WXOTP+pL/ULWLO/bi5romioBEyZSUAV
rLYoTsugBumV0w1qBea/Wryui0eLKfmqJxJx6qDK2PcvqAKov4q7I8gLxKPUhb6V7eL1ljcEpuOe
ZdU5dM6oezrJXkI48Q5KTazha8yfJa0BEJLF2RBK/CBvy3Oqeih80R1c7A/WOdIJo7IoMahC7gN2
NLry8LKCvqkmJ/l1zSu96ggZkuBKqvCe0lQOzDCpmxYWs67mv7jzNHcNokXlIoE0QyWceS+p8/aO
UkuQIYQQoZcN3xCw6TGMc0Ra7Phos86HPBreXO4CTuI/FheMhsBQrbJ5CYW+BvawyfX+U28LBpDa
6h79w44Ab8P34cCPMd8xXkGHOuCrN6I2e444++kCrQZW1elblyI3CVxBByUDpOJLRZK2gZ5BvjNc
vDnZ3X1Msv5ELUgtFaGY5frLOi+VheadgPLU8h/JYKB4IgDm5DZsR3Tlm+9PXKIlDF0/d9sBpxSR
wvweKjYJm3uUKD3hFE31HmnvnUGxxOb+RQA79tncaspsWoPjLXMfgbLT5Zfkny5iCxYWUl0FZxVt
pTHC5NHud6Qil13DLzMcA8pDv9JivlV9Vlvbj8/IauhN7kvU1I4nVCDM+fK+edMPNyJMtEpe2dse
r9v+2f43RYtsZfPF++yuvNK/K+V7IyXoj6fdh3rGQfou7Yhu6sIV1FXNKNw5q95E12aMaCiGnjP/
bo+Gf+/ExBzj4PLGJqiOnViIuh0HPBZG++q14xSEes1KsWVqQOlr34SW43sy7fm6H6J1srFsXjtJ
/W9JIEVXLp23xbkl4HV0pkDRBr4ERCs3z0aYJdEq5wm44fCCphd6PTk5OM3aLXC7xVzlqIbxAFWc
WOlSxrwzoqVPO9WOb4MGe6dPUJPpI4IcaDG4+yKmOMPdH8kwcB3vOv6uMgH2HXkQDtZJaeIoKFXF
+ipSSm3o/4QlOz9otFdF+nFBxfgejGIN9FnKR9sPlguQ4V4UqI3ERu5XZ5/0wR7EGRM27+nEgkZH
YNxnQW1BPqlGmc2tVKD8YSPwL3g/8/pfB0ffhilXFq59TTwc5ltiow9/SGv9N17DcjMW+tNKD49q
EBi0KxJUDiC5zKzOIKKkY3s859v3O5F2TCQ164KGeFPZOXVGg7oEVIQS1As1wXYgGpUVFgsLLTnh
mBsN6Orw1T8bFXA1w7VzmQCN6MLnG40EPljAFO9E96G1BV0oOQ/ZbF3eSFisDEeS1S5OqpDRqsDE
WJo8ElcYcTB3T3fxtuYZm+xUAyDeHgy2IEbuvC7p7wCnOv97JqzIYzV0nsxy/lS6pEiPAUYD7O/X
F8RDPrqgloBrBCaFY35YWVc2gPoPwLE7USYABYNOqbWktmHZ2r/bWW5hofTqvurKrWRRfQqAxUeb
pV5t5CF7508K2Rq2qL7FbdtaTZtiT/Qdm3m/GOvIG7/KP5nc9zri4b71d4mQRoroicVd3hQqnJ0b
W7UGXIWiGGZMDK8qN/KcgcjPPAlOTkFbsAZLiLXrJGteF9oORT3Lihjt8AuaZYVh+mmxH7MBSSqp
5Q6ppykaUs0ukC2KjCZnTxqTdcAJPkru/5FErhGpVzlFxxXy/lcNycBOTVlcqBsDFFB6ZFa382ff
p+gDgV0DRbGdh+Zenz2e0u+xBg7AnyMHouFo97UyCqoCEtcogv24cdHWsPE5GGn+0Y8pIjTGS8LO
VQRPlzEeBtpw1LGp2GGsgvnqjDvjBKFQx/GB8tkpqqEbCYFzPW/8goFK8PwrW49yuf1RXhVu+jFI
GKCDQDhZwGWe1rRq/8JpQ6fMM96Vn8AS4m8hkmEc3yg3RlQn1bySDb4Zz1gltdZZ9khD7Vc64L5e
pxh3kBVwUzi2R1IplnI1gWhKex89/NhzLg4CqIva6na+FIzYphXi6Jl4zbSjiFfcEdjExtXoCfHH
JrjWPloLL2TTNaSsatvdvUlt6T7A0OkXZSvo5kqTjWm62ZFs21vEHfMv2PWFk3GxlhfTp6pqR8+W
ieQjBWrnfzmkHLc3gQqUwtn/++IZ65n8v5NmJ+Fbz98z0AYAI/ojg1w5vPuP1ABzPbH7EGyOILV1
tuxPKApOy+b12w7Zgcmqncf6Bs/Gi6WlrP5rTq9qwf4geexdiZXloE97vab8PiFvFfwHuNBb//k7
a74Kck31yF9KoWzUGqHXxJQv8OTkoukntgHvxVU50n4BKYy6DGgcE3kaaJaarfJaNNX4FavJ+nJA
mo1E9hl6zBDUflhotdfNo56NNdS6T/JOSIpf7OvdPPvpI3KMpwUPY10Ap0PYJ4mLQtQziFbnu6ES
EAqljmol0IICRNI3/ci+veH67+xFFVibYmoc0bKM0mq1MODKpOh5gMtVusOr308AtHtYtEskhXsT
4E8ehK2Hm3gbpGLkgea4h1PBEBeId/1fFzvpRi9Y6acoPQxTZ3iVpmL1SLaIULrW2t1WPU/ATSqZ
TOvfOWg03hnFR2nJQMxos/hhWBlUv+tRafTKIgRAxKwvCCdN2Xb3+3wcFEDnJuWGdKWUIhjRDmfr
/WtzCFA1BdIPdA4JWYbs84o853GON2sWx7+ozaVPD7HNqTJf4QfjtAstLosjxtMuWWcPogcOBx8x
2eeGBUTMOU9ONLBkTBENQ11MnkoPDLPeO4cqFjaJGiO0HTm9p/qr5vqdtugOGsb2M9sw8T4Tromk
4ya84rkDFa++k0DzyZGDXHDURqqg9BZOgZSw5vjKbJQa6w9YPjKhLnMya+3MbrYe1R4G5TtINytE
YKftHSx2tL/4VQSYKnMNSG6nfhMFxsx3KEGpD+wXJFQSIZLRo94PSzARS5IViHyewDpXFolgQKcC
PfT061QJ170G4zMjDMtYts+fLE1ZrnfqL6XZLRPNUr+LYK0BjEVIvEqgFWmx9drG1cifanTM5Fk8
GjPIsZNZeUSVSz8X4q3KEVE5ID8pd1ue+GzRCeHq7XDY68vmMEJu1bgn0MYMSxlw5BdkU1sl+4r8
+riPE0kj89clIceiMr9kl1+dJC4KdPOBMAeR9WN3Y5EFIED9BcaSU5kyZGjDQwhbZOTIWmxAxgGi
SvPcl65px2s0syNWVLIzGrRXj77b0gNlbxlV0oO0+ngvXb9nXb7HpTyrWGQfCJGCM9cQvdrMrQOL
qIvvV3/lBDsUzlUJlUIbW/TkE1GZethfSGYwNyHwFVqDg5zvQ/5hEBugrU/2+AsxUAP4/mDrlx6y
UsvoHspzU2+DgGp2GdeuSkMQv4zi6d2KGpTz32RNXyCbGP4U+gsC2qemwBcKkvW7yE/BGqN6ekH7
/O369ag+RFvH9iK5omE94GbAJaDGkG/Gxce6+TOBl3hncsyQ8IHk40K60mJPEmp1PW6IIHTrQoon
Z8xlxtbhxS/fwnoL5OmKlhYckRFntxkyZKU9mdUqwmtUWhWNZZDQQ9AFZTmjiyL22S7Wk69FOx7r
qDRuctRoJP6mKKDfkVeftqZthfLIPvg2q7sXlVS1J5ImfQPJp/jlVRIhvRadGRN8CtD8bDii/BH6
RAZdddxoLI39tGC7Jg9vsyoNXrcd3wA+r05d8QY+RKZXtCG7SP7DR/6PH5iGGDcl66fcTkw/jw2h
2dvAJRfCD9iWFa2F5aRs4XK9caBK3bAzf/ERTmWxw7zzSo2jMOngiO2M8PefdiUp372TWx7treNJ
EsYgYRdGmhfiiQEoFFc1F6PE2CSauMcuc4O7kaNfIsJRGriQM0+x7fiBbIZRQRSbTTyJL1XMMjDC
4zmOiTvFLXy2QERMgXxH2GPEuExfvjs7Wth4rrRa6F9eABh8R0oweJ53zIZ3/6kDM5D1vYBDMQPS
8eFXi5eyu1fhEtA9D3Exflay9ikNqyJhV6ytWQf/4hbcE7lfo+XZk4Qi0XI5doW0iczQiDRi0+N8
LjYfeGcySgWp8hsJzaKjy2rrLsmuku66fPZgp8cl7Gm2N67cydMDRtxnJ+FYTNTOp9ftU4xxwhUJ
ofpViaWHEImnwB2Z9yvW7jMMLbZldeRsOBQzKcurkHE2hrja3CTc7KW/7YzdWl8lTRSnuAOvqULJ
oTFQggMiXKuJkdcdanhBWrYmixszUTA8JtvrXdVPER3LIFJntS3C/TKe12ZdRJ5A1/zLJJNwK5fm
YWp+8JqaJq0X72P1Ns7nIX59ay8BTxBSeROUhVYg5A8ZiBzWipNLeSG9LliPJWPG08Y6Vr9TAI+F
Hz2fF6sPz+XMFsS0YABGeZlwl+hRjqwnSQWkzDKRP9go/1H1eJ3NEGp5NYVJ2NXoJA5L/G4aylaJ
EaweL3RA0tqcmIQQp7arv5NxVi7DFzHh8nYYa+4kPbikXwEjtLFguHlZohUQwC6r2VyfC9v4bMnH
dCSp4tOmARLsZ4UfaEeFUvYWZYhWtnCc+SiXz3V8FyYp3UdcTvwyR7Z4dHLhgLLPvdpFs9xIQmNw
NXKgx4DLhXvw8tx/HH0gnolq9buvFbmmC4hUIjtky1uVfzCfKj5KVlMwbc+iZYskOq+1ettoMnNK
DaTRtGWXViWMY7fZikUQeefhZjHUywET8KDaCuWzrP8X9zM+CkIZWxoAvyVorC2UwxosrZ+qJzzU
GZKgfiRcHbFt66/j/gCDzOSC8FE2JCGm4JXnfoKwpxPqqd/EMoo7OoOlH4m4VZfkhFdu7g/DOEki
72I5g5bx1AlQbMN/gjWuJE5THqOCBSAhYkYL5Sg73B4wEKclvuaJ1Hn3WsnNGIdHtRB5flLrvhkE
Rc765zL3JsKNnXcCbvjR3yf/IJtSf+8aMbJv8B7hEGe59O+X5sJf3Pp06Rq1Qe4CqcoyVRoOLsmF
Xzg9sCWLWtDWSReQA8W9ixoVv2/0WfHpPL6hwuaXj5mAJaq9qF/GKQTAcNUQgj2Z+xWyKfTfBWyh
F6K6o8VZLtXUzNmT5syiHKsHuX3bHYm/wqZ88OUVsG2HdAxt7uLV/JxeWvU7wSayAMoLwjqkw9AP
3yrthlg5cAXu9nkahLkGEBLRaDf3pMAq3N8jJsrCwjzd/jIlRMPa3/1p135ovJMWa2TKebs7S6wM
lRpuFV41wRJbR2q4mxQOWJfgZWZ7a3q/TjYNpoltER6P/WCAUd5TT4Y7QUHCGf9gqJS/6AFqkKO7
c7WhexfJ8vLTts5diZ43nPozErJKwxOjPRWDiA9xc5Uy3wNoo+elP9okfFEjOEkjSuxEFx/2clmN
Y3638ShLLGnQSIc2M7bFWB3gDbD0OeVGlpN+VyfblsgozbqbkHUqzzmQZjMKl1ce8jnmL0zzw0F6
tIUdva1wvXjRMsQL8vhMZAW4Jidzh3RS/DU1warMqa27rD0uGUeAGRGpEcCW8bdoXSOLaTmZdx8n
RTTY3581E88cXSt/51bouXzJvB562fZbpv7+vTHzGx8KQI1Z9INddRQHNfwCAu8fJiyPRijTvoum
8w3Yqz88Fhme/e+UQIu+zFUlh8pdWbl8ZpcMdJB9pwUBkQCI7KAqUji94aqHhDVFS+AvfbjBQlnQ
sZwk/BfkMo3ZnEtiZE3psXkBmJBm1Uy03KNaLe3+MYK9uBprycmda5ehPuzEWL6wUNS1deedqTEz
fM4wknUZ5GHOOBPD9Sa/1FObsu/lZvOF43UIAj+4DZJPBuKRtIA9k5ftqvD9I7eZYqqpWR0ezdoK
hBbepyfg0pWZ5OPRw0rEbQr/k5WEI99PNMt4i7Fmr144hzT9/PTqPxTzxl4IyGnR2WejHtAr8Xp9
6HkHXjQE4Qs07cpwf2+UYwMlQ2kNiB2BCuZ7u0y8k1D+t2HdTf6kcuiSLCifnPB7r8fA80vamfKB
7NS+2R2Iwv1WEhzMKoVFJ36hHY8KdSToXJ68WqsjsSbU+sFLCdCmqZ9ox7SK6fWAMmXnpwSkk47/
USkoW48ntSa+lG8gRnYBiz6NJk72bCUctvV22cC0WxuZXXDxT+eOxGEmkm99hRqm2G0lxjZv9Lsx
7ZxZZjvw1egiJEIfW57CoauNmZX304S4oJ+Uyl5hs6+sXLTEiV+jxUu2iluj13DXwi/854JUuMxG
pzgWP8rhcM8auu0fKeonC2QYYT6IBorEO8WCcWrG8iDNoCVXdDSzvZzmYq1F/FLnBChD8XjG0IPq
btReytxt60vaHYz0HCXpoLtctSHc86dB5/lQQhh7udtIV7whLHXqYPDHSQLHVTofJKtvl6TFVz7s
68PDlDC9haPMTbbbTnM1AiVlM/ucXC5ZcCLjnXDkVWkymy5yICk0pa3IAXKT1v2PIxnkGxPqPwJI
6TvBDxcZdvq3IHkEoOkjpnL000RGgzjZiErDQ7Eaf/4iQR/R9t+DFZ4xaoWXyRwDNgVYBzWtGzQu
NR8O15v7qGJPy4wQ/Udd0jKowpmAspT3AHaCw1oiK9BLElAb/eG6QRYXC4q2O+QnT6mO/Tq+ATBi
UZgMgaAY/YdwPq1+3z5T6do3ZDaZJmD9uqFpMR0TkZduZggFRtJWX3f6rRpoTrO4rtIGVbRVuIz0
nhcoK3z2I5x/P8KIymjqSgEaYBSqqp96AfGTvbWtYYnL0d62u4NJ9/5UtdqcEZb8L+UTaHfn71vh
EorbYSKEKKiM396DgtC2AlZt+m/Z+VbWXZs9RQmv9Ct94fWxAU/FJhqx+QuD+F2/LKRHH38YYoE2
u4igFeQSWJ2XdNLbMHO61l556M5QNQehq7YUomHyO1MhtyTYvYrQtCEUl6xhL9mcQ7plEgL5sdvr
czs1VPR2YHAhu+5yhta2shKq5c5cS+EOtCIXfaM5aHSCulWcDMjmc3WhW1lrmiLRSTpGfFGervfa
SE7Mow2J0b/917jUtVrAlmCv1hy5vqsl1/MhTWWhhDLdBkKSVpApvWOT7aTCdAn5sPzlgKROmpuL
18tJUQP+fbU/5Jz+54hyyE6ZPfTZdFkYBc10467ywtcQkUo9WPGkGveVXnUefr/v1nseaJVzIbWu
h3mjUweHZcy/hmDDsGHCJ+ijVK2G+fyGanZfJ7fQ8veWwiD3AewywGKs0hYI4ypIn6Q3RyJLIj/r
zUXVcfj7Ak7ATGMHTjq6Xb1uA0wxFEPT47LyT1CWlxPtvo0YQjGZHyy26nlxSPW5lx/hL7L3V4Zn
UziM8Qp1VREKqF9LU1VddXjAzkcvm08geB05JcDrVK/zYFHSC5gCbIB15f18WSS765oJS7r3/JPF
eEFowgtcFTA/QBeB8GgpiP+tRr7intfVeriNlQAgc715fH1f1HkG09UQ96n//mNBBquECLT5+GMo
54ZH58/uPTAh9Mbe9NqrjhZs6gDdAf/D6Qepa6iMfhiyWpefKCRPfJpjaeaklVVAOP7IqjmxHzne
SIlTknKtGrE23y0iMYyO2fZHl5MSbWHpBiSuAYvEqXAzUu1KVsfqKAxTcfEF9Nuw1ceAEgqfWAxg
lA14TGXEtaD1SN2DFfZ6xtMfeVaq2VBsNAdHOK7TWTWxkK3ZbGmbiJBGfdw2jTplWNfYA7MiSVDO
nTJECSKzNOgx47Wr9CC6PVZWjVHpxMv14spthXLD3oScD+4tBEQHYukPKkmKzbSOUJrpfe0MRCv4
OqXO9yfCxjiEwGGhfFhXLsR2HXLeXsvLxUZZIr3IM6ZpVheWfCzJSpdtq4NN5Z35dzriyZQCuqcn
QVrW6NznvPw9xATTGa3k+NUm6wDgw/jaDPb291Oans3KnQXttZb4SHt7yn5AFrXfq6Zxj/+d8X6V
QS2jvxTD52uBI2zuSwcQAw7erDnmWrwelfGw5pXc821qd1WCTBZ0vp4IEI5L6t/XmYyQRm/kSerg
b0WSaJiSy7ri1aHipe7gwu3lAlAIbp6nvO7ywc2DujmW5ZTIkWsY7BEPcj3PBhlEVHX3EaWJODH3
byqXk8b0NjDEFc6kluO1oBV94F/M7JiISM/qh8n+3x2Cyq3etQRvuSqAHcqUoiwJbCadaXWwZlKd
gJmDtq4uyPDDYZKc5LfSGerzQSCElIIuIvSxZ7C8NBgXmi+IrzeiqMe7j3GKFbuJhgHm+DhgB8Z+
MFaGACCVAPAqO4fHBISMc4gPDej2kZwdOosAiSTNIiRGicdgHoDDdOjJsSgXjMiKfEg6Eqn0BKpF
f6gdwA52dtYq6jtwByKfA12ZB2FAc+TIgXkOVxyMNlE16JODxs39AWtH6R5yqo4eYwhm6Ezx17+i
wsybxEvrmMY8gjysfE+dhdAM1NDsS86MpVnC4qqE1MMh9afF7vMrL/OdGcjRcwoFLGfSzZ6pwo7y
YFZ15ad1FE/CslcXKGlcapqD6OjKVBCS6irEjpqlQpQ6nvsvlgw4C8/q3vokNc3itDQ7ozJ36oG9
7+N7r49096u2TJOED0HIVsuPOX/LmS1L4f7f6mkhKACQZ/JuO+53ZZDndExikznglAuVt2yMrMSh
bMJrTO42RLCoHLVYwSjlpLq8lLZCmRRaaMkILzwNaEqZnLsRFuoNWWYrngn9roen9/tP/Us8K40f
a+91jm2ZwJG4WuZW0Cr1EteaHVCvt/F99si9tQIN/wk5/e3RuDIi7wLDtTKUlmCeYmtXRtl6McQV
EpqL4DeyYYcbWGJ4s7nAwJsauzVJHJBPEjSHq8LNWbBPelyCxPxtKpcdrLtxwQ0O6bVGIxTabF/N
5eyBGryreARsecMbqq9DObikDawZIf04GlaB/50zvx8fXmYbDjrUspTK8FiLAkiBoBZvn4BToPhx
oHwq3XqODQYMo5QMHK+VgzcYduM9XvUp9YWuoYo42TLWazDXsHkOfa847dwXxuQ//gSSEohLZ06C
Q1J3DdMhw5CELyiveqxGENUdrMAfVW74aB3NBfeZ5SYxkCVPUFJd63VzMRBRR/30v8MG3RyFA1G1
l7ek/NhKKtCw7fhhJfVN+cdwOXASTKAdpsbbh4eaJmZvoEcLD6uAD9kO3rFhpFXQ19mMSKNhPEg6
+rRYCIRq3b23QuYXUCys1rLlbHADcoZGKW0bcftQ8W47v9/0Q7hSuxxi2TVLpFlrKJtpt9K1C2Hi
YCvP04KG7nbtK9kkgmFyt3bbMr8a6cdeVDqYCdQTfIeXqwhdDBXGp8Ogiv0Yaqp0u7hfukwdb8oz
JVYdSBTi83vJCwOM4446F2CSvDLvs6gVQApHB2KJNp0cSWgh9EjBoNU1LMNBcYBR5j2vQTL7eESY
u87YCBVjEEDFWn4UPk7La/1LDKWJJ4duSHAW+A1/YunO0DdjVLvwjX8bqbq1L57xp4BlhOV54I+d
/AH0pst2LS7BCz31zejEKFiWHa0wfFwYsx6PCGdTeZ12RrA/gI9/kFQkYXd2QcyHOYoatSP3jQc9
PTeQVQ64uTNRnME/P9QXNo6pUR7nzfmK2SUg9dAy/yKr/vaLVupTfVlt8PkFyoEfpaOetvNo7t0o
Z+VJu7awuJcQ0Ckw9kQNRZ586iZ+E7p7MVdcSloF3OIwAtozN27odjdQTphI86b0WnNuwGvaQhjL
bj+LbWYxZP7wUmofekwOKJI1SlmUZgczOD5jhNV3YXkQDZjIsWJ+jEoBs9Sjf6OM6wLt88bBC7Eq
WhskbbUOdJn7DzPq5XTOU1X9bVL2ZCS1DASIp9VPdT0kT4TjucVi+wpPMDj2WsUCarPYCBFhl8Q4
laqRcR6a9z6+PH+xZc95GFxuKcYQZEx/aSGu2HTP02JWLdTNnSudJcdw41z44YxAoK0XyAWzBJ19
tAkaMx/s5YezlYsPJnjncpgRCXA7JR36/q5jXWxDrm8Y0T69L/TaiA7OGVdwnklvOvrKUFrh3Sfu
a0rHaiSs/x6gGpnFg14tAMbMoU3f/72CO/IB3YtKxFIy/Q+9RkJRr9/8WxEHfuVcd6gglxSsEvqF
HV03FY0Zxky0ykkXC24oMPXk8nR+vfTSCJb9L9Shw/Y90nTKhQDtw5wfv9dsgQVo3N21ke6s+5zo
mfxDn0IW3rVZnMiEFCpUdUyFPYA+ycrgm634BEB0ALpQu705MatOLqEhSMHVoBuRp2An0cG5pDAG
NZcW9IfI5QqHh91C+HyisOu7mi8Vt3Kl1dzxKnf5N4LCd/awGBKGqtxcZKQwWIWkuHQ1EGg6rDpm
0hEhFRQiaZ7okgLvHcHizDv7VAXwP0/TbN1oFrhU6Zu+EAf9bupkjV43amiC3wldpNHlL6V6iu14
qYFkCdGprEmFaeqvAWMu3MBFhnQKg3JQWoFzARQrw8dwkgRH7ZpRhinPNYRsRechXjo63R3FSlhH
o/EPXygsO7ggjPq/TkddrUQ0AxYsC+xs985a7FfcsFVTbTRgGi46eFz8aKSZcwlwFEVW+kXYFjxm
PWRCzoCs1QRRvYv7CeV78pFUhw49ISFtmFKUtSYmwRIhXNyKjoJrrMKcYV631lSPqCjdidMX+TMg
Db6XL/EpPsc2lhL0UL89r0ja30tRZN5VgdrKIaQzN8VqAzBXamJTqocL51b056v9pVNpuLJHkUIO
G5q6iB8w6qVg7W1MxmX3YA4FdT0zbQsiH4D079Md/lVAEC81ztguDXShb4HUIiM9WF3B+Jks0QSA
F4kI4fJ5214px7xvkNMga6KXZyyE4FzDkUpgR/wzdxufYL5JtZ3rqc2kNzqV5IAb/KrAy19R7J38
dER10hsJb/l0kx7sPAO6HdZO2OM6I28hYTb76xfXoLxXTfoasH0F0qPQk62lYpEq2chuMHzQ4HU3
AthnZk0rigyi+u+2TUdjcuFAWRQBLXnGW0D9UjBWtGL0TBD6E4swwgUuz3/5jWc+4IBuovO4VNZb
C2vyZq/9UJz7ZsFxowCH2cm5aCZFDmcZZZ93UKfEDBZjHdxlLCD3FoEMSkBEYFaFqKXRTMvvIkkJ
sB3JAL82Du5IeUhHHOAS3wLVJGonZ0DDp6JozKCp9EVvncXnV+5wt0q0lvzhyv4A9LgXu7AS8sAR
El+Sx42gMj72JQ4DIHxne5phIx7/vmhsoTJwFjW8ahEG+u+S+FV8FN08AzT1ApDdOBBt0J38Ri7R
9Lswdxvcpsg+Kcj1jmNGsbLmkNPcBsE6n1MPtb8qkHqmAPfxFQlbepKmGUJ/OSkFmyiIHqy7+TjR
eE5J0HnxAMHFQlSgp7GM57Mw3OVEc+15WM+pCt+vEYIGIE59tO3PEifYUSgZsbuvVJhk9FMnW0H5
6V5WuCzosJyPvVuGzFLl8AkRLlTXis5MyFVFycWprChGUCnh/8VBhBQcxxOcUNX82G8LPligQre0
nn7F484YTLOMWHNOneMFW1VZRFYxSD4aex3ZTnz7RF3fgqB6uUiC4i6LJx7mBbTvtdqxJAdNX0cd
4ssph4QDvnDoMytFWGPdlAnFB2b8SAinBQmVfluYjmgMwSyUBOvCI69Db75OVwIrXyARIRoBqkIv
H8jia/80MR1Ixny6kw6CJmf6svc6QJ/Gjjtg2eD3bF/a6nSid6gg5vRxAGOOgDV2DMyG+vafQmhy
qbeuneviif7893JbKWJTpl3C09WuPGHCJdVcCQ5fQH+DcvpxecgJUpGSS/n2nWfm8Yvg+ka5yVED
lWuP5nBAKX/FQSmukMaq1merBJcjWFOOTsJHnEOug70cl/Q+dDF7r0n94s1htc+aek7eo4OveD9w
r6OZJfUf4vS57Ip4MZ83Xk695f9z+y8jHk1p5lHkSahamG9YDo7ZSG/WVOnfykdFyjXjH2fVK2r8
QKJRpZFaQYlLgR3jpp7wv1R6kEPtLSjFUfEPae3H2z9/MrV+EWEMCHL9ElRDGJmz49NNnbLtxZ1K
/WB+gWY/nYd3Z0THJaKFgp2VRJx7sicqn24EwanNpwMKmWhZq0cGwJFyolclsNIK8bRoL4FjUZ+E
jR65ce5pY76HOVCkC12FD+Ss6g4PxsmTZHN+I9nA4+CNzENBbavfOKhRchKuiNK8b1ycARQv1KjL
vfyZAFSaSCrzSr1TXZECXq8zZs98CPzlRIs/vqMrjmDR8vM6E0U7HxbGqsPQA+mz8xxim92d7oSB
Y68Nk6a/C6zxvxBkWOHCHXxDxdIgL95GSsbkiE+Lw8TsvVpTrW06KQ9B7NmEEoAFJ8lJbNAD3dpL
ZYfi3igrJyHCDYb4XqXN2MCxbJiKKk56YZWGd/KXVUiuaktW022oPUlBUSDIBJOGWRzWS/i5vLqb
Kp/fmcQ1UVY21mNM0FrQqFjZFq9qZaUXcr3B4VBNCqi7wJpMq+G8DJXWSSZ0iZhLbbH2/olz7QU3
KChbyM1wHbYL9Z0LXUm3xAjzBbE5Ml7Mi7Ca5UDc12m6JD7Y4P6mn7TVPwS6gVCkfMaSuO3u6L+8
VKoZJfe7HcYIZwEo82EQxpyeDZyTzrfZBSkUjqITBCGPwN3jzlFd4K1NzNeii+VNTZlBLQxLWTS6
iH28fMnaQ8dwtDZQsEc6P6VL1pFjBiVwkez6sMDWuXySMI4G27EGig7SJNWTsjyOA6atknf64JeF
pTIe4+oTLzWzSYYPfVwGyDzjh09acSFfpc3RQbotwMV48jqKMZueJ8LBg6TgD9HI2wypS/RhL5jB
SOhn2Xn8AqVZok8tn1SbuFSZj1uL0Z/i6yg+INFvERF5k8u84l0nEl2xFmGfPHT07Ye8JDUAMLzs
XpYjMb4lkxFlQHjRbteDGlBcAmurIuggoiTPwkhkSeoWlTm/Bs/aXTrZE6y9sW+j3APzMlFuNn2x
ETXyqywzGeW1vQ0PUfuLVwiFtLctk7sYh8V0qwNH+pa/XpRHuiWHk2PJ8qwmDC3bSqGudV4SrDiP
I0DptQwrrX3y4TwCof/1DWaDAsa6hCoq0lq0TcDBAoIGiQgus5+ysmZ92K3p6bPAVDw0nTtVlDJY
JojV903usFDDtw+JgRiywhy4XUHMjkgzOW9ZDUy/Od3FD0fVPe6Jwqp83ruBxc3rI/+ElGSMKSSY
PK6ZsPVLhYUsMVgQHqFpMoCwvwQOu1MMyqgjvlxn5ekiQKyvPyZk6mwztLHQ11TXMmYCb0IxrDAl
IJyC54DGvqoRtoen1Vn8UQcAQbvCg9R4Pui1sGoSc17Eu1LkTe9UsoXeYCFgTeNBuOozp0BxxY+E
G8tlKM9QNo6+nTwPisgVbxRIb5JEauWztAeijwHyLycxfBXNM6tVW4sxX/mmDI0+UscWulWR75YH
8/i/tIphXLuFiyVvKSAJqpo/tHVKZJVhA+rEr45d2REmfQfTPC+/ljVNNM8+uJ1ci8afrJCbMoI4
idqRXoIsumxla7UVNam/CUALZafm5gnRSaBwXriE6EHjO0NpI05UwTfj4bF4eSVPz4gjL/J8lN+R
dXm2ZtXOXR/hIEPx81I2U24pH3rF5kb960HXdDOaWhv0kcJuGY8JeISgSiT3KyA4p/sAd5Exuiwf
A8DNNk0gqtslPGol31EGpozX9bL+RPSi+hwX1CMCSC6kzDSN7HMeeCyW/rKZOQcMgsEzinsuFQa/
FPpN3L/tEKLUdLduoX6JSHKg1BYP1gxlChowNGuP8+Tc6d0pao9RMTnqB/L3oyQMkRS5fJUcilRU
ExJ7Y6wR+I7IUYcdTQsTOADhhhakrGRAepAOys2WClQjms/MWNHZ+LPdg56Gi9DXOcurRqIPBaJj
P/WKbpHtTnsN1n0oepOpB5ae/mPPjKn2cQPgPSP7ZQ37dWfWYg1qrs3j0wJOTD5sx0Pzx4WeBU0S
AT/MPKo5ScdmxanDEPf3yVD2cnk6j0D78xImtMLZ/UOrz5JHD4PgoFEiQJpnjQUTvI2Aw/UqZFLa
+6gbKnNNiS8VcXo7GUslR8SGkkzUlkA2beLl7SGQzOEXwi1pJ2Y30Pg02/yMR/YNBaAph2HX+FLJ
+x2t6WaNvhKqIvFjeLAZ5fS9q1fgRUHNRhigCZFVmk4GHiVmXurCk226grTvsCzaymF7ADsoCTG/
BlaoO97nzXHXpzSvx++gP82D5AHEeKyBKOivJ4u9BWjDPNw2T4X1YDyRCQS6GBiBGEhbnH2am5Oa
YCCZbcPgUvUVYsuEZdxh7RO/aNDhNAHCDox5BXY0kJRWEZPNCHCGLoD0pVnqzUmR0oOYsX/+M9kc
0+We/7LKAqqqfzvMCt4d4kwsEb6T783AtezZBF1rf3vWDD9wPE+xMvhlEfHSSnK8kd5ibVtZ5itg
/uqGLYTqHTI3fbhrd8LAnlD0aWmVZIc7C9nUN1K8J65IBEDhSc1fzgTkKhEI9qWA+CEIaLjykGVH
12kkKTldKK2VmucwfJ0oKf/WPjObttEgDnCWifobYXUQ0bGrc+UWS1v01T4ybJ+NJDf7goP0ZLYY
wuJyoRPVeI1bc3z/dpFrn/o2yWuvMuc280rg5rVMWI4psiIvGB3BiFhunL9lQ8lp82f2IbXyojcM
fGs7Ord+6jxymKPzHT7Sk5tMcVj0gcxHW9zyAC+Rtk2DASphyc2kZc1avGb7oA4QK+efzOaMnEU5
qwzbeudG7W2lr1LQQFYOSwKHlLMkEmOPjgwA1RBnJdMs6UuzFyiNWD5f3j9dRXkbezmUF8LAptsj
oSKoFm8OB3NnJV8p08TNt7XIMfQ3IIEX1IimqLoNaYz/0yZw0tnU8mdZh1+N7e42mWHfgW2Ofk1O
xcHOKd+6nq529Mz6OHQOn0nBVDxNe4tzO8mngeKmkp9I6ivXu5tst4/dgPcR8g78yMxqVr/vd4I7
TPdTZiB1nWRymSB/MX0z2s06bk4Qx7p0nPD1jqDMQ9La/hosY88mniiAxrIjm4z4VTdNY4fYsWTL
s0rq+FxuNxMAWcAaeK+Re6GDJJBiTYaVVKKWAbEY0L+u8OhB6LCHxYexSi+zxYIeHNOM9xkEpzzY
DzBwXlCpB28YvwzSfhxpKfFWDftUX7UqX/+nRREL8LV5WxO0JX2J1BzVV5aR+n7JCClzNAdgSnQH
+2zNRzrdOOAIBA5+Nsnn3AIMaRxNozP9aD4wZ8EimRqyvxfvEHa8+Jif52+tg46wnTfIxdy9ztsj
JFGrEr+uQb6IRQjLeD7i3x9iksr7XwIxm7soAVJW4wmmj+y6F85Ux/6xxRCNEtcjbiIAwVVmoIkI
oinPFH2uUvyUKYcKhgPGE67e+wKSkccctn6usOJBeyZEUfwfOGlXNEz/ROmkBqlzo8X7z2+AEO/n
XSGJ7aAMVj79XdMkGbT0JwV7289d9ND1L+hSpzMju7zwnI6F1UqzVHeaVwo54jk7eyk8pDatCSF2
6AdWuBEqL3q0jQNDYy+T01xLg9PvEseTSKHL5RDSBMzb5BbJq440lf0zJuS3/3q4q6Dr96IQ0NBk
HvESdQ10O1DPx/BJpw9y4sD43Kcqn+/c9Sb7458EMbuqSzdiacjxP1kSGVlVwlLwun4U8s0hSLR4
3AzMbIKIgzcELb/j+i0UAPtiokv4DECdUjAD73URK39iw2Agigf7VnJRI0r6kswnQCoZtCWwwq8J
wsvKgCPO+YtYqzvppxUBBEnOP4xvLV9x1Ty8fP270LimC/bQ3wq7VCBZhWFaExipV3ZChxqv2yx0
z/bJ4tzlnujt3MINBiD0pTB5GlZlrCTmCanmYtaiVir3575L7Pi6rGRDFC9c1/XpOa0ErA6PSyka
Rrbv8lkzEG9RoSt6vyP8v5jSs5oC+YSX0hRQk3oLZIvVF5yX5snJQ13cWV394fPU2saV91qQ9dIC
SJeUSQ9OGzM0moma+e/LuG825tD10jwY7/G/dc9o9XNqW/4CIxz/axN09OpZMJ491Xb0h9pw/DHj
pnxn0ZVOP2jih7x4hGImAVorfUtcetPvzNRjkVZwoL7GdefNau+lwO4uzNZfDqFDmi/06qqLQwvE
8/FnNrKA/AgRY7955dbOhGwNTuWcRhI1W4Y9gfu5cMHCctmfO3GNePgpVPb3s70QpcsHloBYBqEL
+MQnZ2ALztQy396MTgzgxST7AGj82qj/vnZDFIe0UblPJuIl9f/xBBxZPe4BF6VWl9XBdYvzSO7I
s92EdByIsrshYhakHXaykVwlY4aYHPsBlA+Tw5BeLpAB2VccJGGTHEYPU0PSe3LamexTYlljRNtZ
vl2Xr4RULLc0+8M33uYx5UAw1MV/HkkHheDcWYEMpaF/DkpoLDRWy/CVee1qjZ/bSw2d08XxCSFD
dMNImNKgwMbHsI+DCnkzPQWUELtXMTRVx7J5OUFT+PCsdsPwXp2gDxPhsKRBIaJro6SRMq4Xp4bd
yRGqys93f1BQNaFLLpqfY6CxzXQl1JLt1cG1UjJ0fVsNqPRvK4uZ2K1K5hz5cQN0k7QS5PDuDdE0
yqKFcy2QteNtcPFh7P8lc2tRtJ1VBH3Ep4PCwg3I3mpnYEE1zWNXRLaEuzqrmLkAR/ZYDnyF3oV1
wy4Qdk0GfIvxyCVICONW4GfcY7e5LuC5gOysHxkPpIkx4Ydu24tV+A5RbCmH4opXR//OgwKjqFHW
kJxlYh3b+G04t8BOiMhFYX3YQEaGPQDCWgjN5KZVhWnD7LpZDKsba+/GxZxzLZBoPrLR8ExUfPJo
NESLxYVwIL1inSoi4Kdvrull3RTTH8S2ZWrUbAakVsbDupI/ZUmJxRB6hZFK5qwd8uktZLaBpVky
3PfnoVK2Gwap7ntZ4O9VyuXQ2+F0j++YyiDBB3PKIBg/LgTIhcWI/lgJUUpIK2eFF8P6b+6AJsfX
BNn10qG6Lm/LuEgoEjGer7lbx9gBL7x8vy4sUMcw2v2vBf0dEJkAaUg/8FkanvEpJXGQah1pRuMD
ZcS7ZvvpM2QngdOyM8GUB5gTuHE7Rnn5phc2H6oWPXfBhXCRrtfBpEBqJBfSU8h5wAcaWeR15T90
41wqd4uEkXEXrwFtjEgrZEfpsdMnUffa5yLjLgP62Fq7zbb6OYosW5yHM2MGBGp4uU9RRx0J7oqz
g5/gonAYgCt4KnOINXuD/oGNcQgFQgcns85/UpF/dh0yXRPqOXOHG88vZDj5paC5aEIlghxHfLRf
OKO9Pa4rZNEoLzYYndmT5PcvVIsWr7x/buCFB3V3c6+B4t7IPO+Ojd2LDUAfL1jY+1GzzWZwluQP
t5O7cGPYFW566e9XHZra+yM8qD7cKKqmIW56bT1160quv23ELnOxCPMG22i9sJGQHOVxQyhFASHa
15BrbxwDH7IMsUPkOXVA1xj5x6JrVMgUpY266/ZiDc48Yi0ronbiG5lMUTK0WWo1fPw8EmlOJhM3
N+duWR+qasIbdbScLWsmH4OfEe8GzHX2n9BPaAIWxTR/3PE0e5MjsnGpsJRFBtvCGlmtU98VRwwl
IA/rQu72g3ewwrur1SwL6KFhCZhgYccHLHgdfmBpU6HS1nE9QdlMnHjbdiFdaFpbqaCfxMyqN8sj
rjMELB3pzGLQYA5MmF140pcQMqRe2ruC7CO+dcyo4X0iGGn4Ia+gAw8zhItTyTTMjopvsyjvQy5H
neHZpL+Wls1MZgrWfRSmUg4Qnkm7ADlMuGRtLLTAvD0icZzrh4kN5BpFjr8/c9FuzCeGBfJ6RjeK
Oe5G4Af8HnCfAXUEBfwwMipeUQaZrtC8xGg6s+PTQR+Eovd+Vdrrh7okgCkCuSse2jm6HKZ+vq+j
KeDnLydzWjvk9dL0To9kxapVj5eSC9Z4M4Kctg0bOFUwj0ChyHwkcz95ud8SjXED7JErmm8OqMRN
mYVY8+UQt675L8L1P6/77efnFXK/T2W2hlo+5QTsjZg3BZqv2h2FkEC+aCppCBJgdzHAbR49QgMR
uxxBBuhBeVY8YWQYScMxTwuhW+ySluHeFwtgZiFsjJ9LAXetWGlJz/DqE0RrgRzwZccVg40w4nAV
CzFfxjcA4hhgjeVW7RGYxhY1cN64cUzsUjJVoSAl8uNEu2sXb8cbCgEM/9sNCT/Qswlv5OYmwFG9
m1/G4qkHiak+JM4bcq2aUM24CJutaLVWd51myFnLvTdfUYooQ+bmbdL8FB+r92Ed2zqnAgyieQZQ
OVOeO632r40iPuwURdNHzOK5rKwFBATXz4SUYG+My02fiWsdZsvMt68j0QhsofujX4c7hNoRW1xr
25D70hV/7hSLHnSEuzt7tlyEHuT10wZ561SvJj3seQ8phppQIRUijoERbxBwcKm7muVieVFWxuER
hAmEKcy8dVE/uJvy3CuZM6PWzD06KSTe/SN+lBAO/M8QIxn0L3ojvAREtgbInGscCEL4oPMf+ZqL
MWeaxgl+ymnYt+I2Oe/L4MujFCAvPnrlFDLLQsxp8c8u59RT1YGfeGj+wgIiVKyQMmg8IDeDsg9v
K7i+WH+zTo7PPi4Kn5gq/ruZFc3cEevpTmF69Xpuh5A0ejSupbJCxahY5fhFax78xYfz7UDot75X
UG1a1xXUlhQWDFGP6cvYxPi6wzJcBi3Bey4XrwJSb0m3/EvBheP7POsP8jJ+Wy/FmFZ1BZzQGENj
1+Sl9dkPaENqSnm9mjsb/t7uWooTYhoJ2B67Is3PNkReUADXcB5YaYtcuLJWphrggc64lr59s03K
wbtXtoUYESLzLK1lHEMc1UuDxVpqIvHE8hM72PzbZMgqIqha4XVwNulnyj1gJ4TtU4i4I2IYfQXi
yh+MrITTOQJWCShxj4Ut0t1cxL4pSoBAUp/ELJ6lk1aDq3f4oCnTfAkjmJ953w17PqAVKC/mfHum
HzcCmM7SC6oPZ0ZebR3YVsrpJpatMnIvNm55sI5cey3VTS2+BAGdOfA18lED7n8cKivliEgMDEfS
EOwEyDY4yvYxQRSClDzbVs4fQdeNPKyhe14vM85rB59GIPzbcpbezy1aelMFGodkA/ZQrhSBxTWv
xJuy11IQDcOzCTzdEaXKaMAjpqkY2+iknjWoGvuZcT3kKlsFHeVPdhn/NFI2/bDXppew0lmZ8ZrP
tBjRKE+J2iYKNJBl8/wIvXu8UOqDFO9BXuoACO7qAjVZsB1LpRXI8Ma5XGFl9OGUn8inifiPiP5D
H8uPw7EC1kNvh/3Ovdssdzh9d0+6Hj5FTXZiVKI0SCxsYfnUoHbAO9GSwVy1dNeuzezz4bzaTa6z
Py5cOPu0hgHHW9JGiYW0QscKO7E13NCHcnPl+ko0J8d87ysk2o5SkjJA6MR15Fx7HO9fhypYGc1u
woJAv8qs0aNlI7ZUslIEiicrF2fTvMByOy9Dpzo9mlORcdqJRH2EIp0dvDVHY80P1y4P+loCqq7J
kJALiK0ymNPcjBFNe6jsMIvD4BqnYiBJwqj5PIlFeXZZ9SFidsSUlM2U4oIc06FyH1ljx5qnTRgj
OYg/wxszNgE6bwmjF5joP3jWxATNQu/wefmP86C4ifHeh9EXDlKLec6Oc5+RhkY2vQ/rPaus6/Uy
al4SQ1a5xYL/mGm2eOQArWoD8v7OzWBCu2nJYChQDEuZTXY+pOjHhYh65DfKOCX39XiGRtuAZoOc
mJl+AORZvbzNaayhJ25pZ7/HtVfN/bYrSZXFvoreodm6EVwhRLB6m1Sm2a1/2djWfNmaQuOCwb92
GZGqM6a/81qnLOsr8QXITHMuS3/brhP9Z2pE1XMK4P8C1LhDAA4J5np+IeXRheiaBybfEj1iZoGu
FM/vG1CXCtPrDh8thRVGNkJMcKbuYwCSTTcmyTS9vDNJV1gp/kWdXK9YSs+n5ArfjapouBstcBCx
FhcmInFlfF+svuAtygbCIypanCOzGBAyFcX/Z/UjWaSuxd9dpxjtMMXD+nzJi3QExBHxHy6vzkY1
7sG7DRsLQeMqebACMUkR8GjgI7JN+aAMkRXGp8YgbztYMZ8KgalNsTAgB4tsE4VcFmQTrEjslms+
50r6NUSdzgdbkUS44LgIpoE0O2arhpC3xiLixtzMKeJlS8H360I+tRSMpthZnNyIZ8PcU4jpfk3p
5GvcSoAHDxHyEmURBdW78buSiWgDj7QKapusWlOGkcLnEA2czhUreRjn7wrRh5aUaFrLEbDnTXy1
uKH2MfGySyG8U+aqzXWuEiFplIpMe0IBDzCnwedWa/nE+L1K9dx8Nu+cjB/1Zd7U7FxYCbXCejqZ
qBKSXadEgQgzW4lMOjizA/YFnPeRhdgZmdDmW7I1cDxRyuyPplwgVXDkh1I46Na+iaFWoF3fjdbb
cizmoLVhHaFU4nT91X1QG8yYDzjqYUzlRWmfM6CagAllnywDO/JAG03KJMlGG9V5DZVbvH5CqJp8
9OBc4PyoX78YU8NQNw4j7y6X9tThiz4SlOPDBmXcrS+0aLRkHbsfBt2+fHgo+tJ8ggeyTN9lwngk
2Nx65nXuq/PPdNoGZND//4plScworrrE4Efww6uubaEwpl5JZvEbAEGG0AScCxYNJf79jw+Y1SZM
M4yaRzevhgHvlsSjZFIRXQrwf5EtUHM5bBFs78slhGctyZQ8rqFrWnidpeoKfLmMXoUU0La0jcT5
oDXUXJcazlyuFfX+lnZb4kmeh5V0AkxrAHyGig1IrjTsMM1Ze30NZPACOCyYpmbN3jaacu5X37Js
VLGrsPssiMRoj7jThU0GJYekChq6ZIgjOZ8uNqho01eV4ykBN8KA1iEaid3Hnwq2EkCXYH34hN1k
gbBJ/m/B/lSTt0bgq5xiOrBhPXJOlHID/mJUuzWV/aEnIpf4LVcV1/E/hZ91wtzWSAxePRAJNFwm
gkLqQ7rlB75ax1z9AoRQcE+8d093K+N2rMWLmXME/K+Ah5TC78JpdTtyNkRbnOcXMNkcd37FS03q
4bB2kIezrRiGsEZCIuCmUmbg3eTn20yqV37ZmsGWLvsOEaxVHmAJz3VOyVJ4y4F3EaXPzQVnYEat
8CIG4JPr9FrT2FKHsjFjLcWPXzQdKe1Xm0haQCKZ4B4Kuux1uWw1RaiPtZntPnp7TqPHImSb2MLh
KULcNAVqiSiG4m1ucjGeGordaYx9gNxJjize/pllNWvy+bPOpV8VBz+Naw5BBaz0Rijetd4Svnkc
uhEKHZk82w+tabVsRxlhn33TF2GFDKMWvlQh+38k5Lv0DH426cRlxhOeKKeoLk9TfnonPzcFMCmm
ZVwQ/7gfFTkdgZ3arx9GUhyCOKxjjKCQ8eiZ1yqKjcraxw4keexcUx24/NiZzoQ7TV4AoB87BIvZ
B4/n+lPlaF+th6FRgqeCQC7VdmamuIxoA8tVvjrfb2Q2zUkQWxZRKZ3AKO8TWiqFv9jYjsoHuUDD
NnlY8xclEz8/TiQp+Evcl4W54b8VRDLZ8KdJKJNzKAU/mI3J2dzl4/MQNdZLGmkS22Omz2is/h8F
GPf69E4aiNt8w4VZZ5CS9MYxofjX9VoG2YodCdE9ED/0/iU11RSMKx9FhCMUifAVARBIdmCs2Ovz
5UI3bn8MZ/VNcv3YE8r5XCUD6Ti6GZSlSBpw+TMF5sv9pn7CBBTCkOpiFF6rYNQvAEYIvq6HbgMV
Ckymr4I7fWE1N4taj0CNeN0GKL03FSdr16ajodKIT7fR9x5+DoUZi1DCSEJlOCOfhDnmrrkBxvJs
9rVaZpkD6d659tzSQqOaVlle3G8zNnLKBdhbFOVYJckbQZeY07S4l04AmSul8IY7DczLepIPbHzj
/Lj4HHIRiIAxaHbNIdrJAFsRJdmlgtdaLZMRnXtYV728vqctdBikur3VFfj//r4oMZWjyDXal4F6
KKB3BLXTgYJVp6tGXWJMLIunqpsG6toNcptPbqlnUILkff5ICnsAkXD58iLNQyQxNTqGGwGvkPac
H6MpIwrVWC95Q5UeZURgF/Bpf5Gc3J6p7AMuFH5RR4hfPld6LltS0KgmUSavRfSTr8+h/a7udCB9
Z+5Fbv1ro6BriX4ucf9qhPFQ9N5QFF6fhGHnh8CMOn5HfSgAPLgRxm0YuX6ZLsChl1smvhM+vXFC
DgyZZA+qNxi08yxIx/rI157vUV7ZW4GEfg9MdtE5RUyKznQbH9j2ygbHTqCo4iy2IzYZNh2BTc7C
2iOhSn2kfAI5knHMNafjsuJcJowaHgN0vRclphGeILJOjkbXD1F0Y+eisRMMx2clGvmb8TPgKRcg
2rHhi2v6VD8vZcH4Q8S46W3YaYtoORDmAeeOSP1tlSAseX+GfmC8N1nb1UkiNtyhoMUpYJU3VrMe
eYVuhH7rmNVeTxhOKgCKDF9A7TvGlP2yQw4RW5SBOXa5V820Uo4Mm99ll9lSdNtOiNtweAyLV/3p
tjYKVmCaTUo0A80Bz9k9M1LleZ7lKFz2VHbUFwlV/8zI8/GGjO2AJ8uJ2h0TrcMPAC0VJngS+SwE
YOR+Bpl+RvvqbuuJJvJtGWOaB1Bx1Fx+ppHeW6oIP9Ra0nHjeZe3cLsjyzgRx3gJydANVnIxDQ2c
dM67BbUPEW6UVc7rLMvtJn/UeUr/zetufWq7n8SUJxNYDKg3oIhIxZYJG+YPDzHjFxEJF2G+oedp
wBBc8uWDnbepTc4YypH/lH6MuryItijfEN2zbVTmJDOVrGb1YsAu0xwYw4gzwqo+DWGURSUEHvvY
OpgkLtI+YlNnhpKIHcftj+bgAdknyRMtDbDfRbm7wFi9KBG5J8I4PrbEe9z2NciHjMKVyDd9pFmE
UiIfBzFUec5HJWvfPc0Xws1ZGK05P/y8rqfQb9cfOEdT7wQJCbsR03rnFTSaiELpXcbyjMMjGGM2
ZcE32W06Lcnhyzg0wA8zZVoJkuQyrliRXVs4UfYnY2zXxYT0x2Bi3i3so/jYyQu7L5lxqkI9gXjS
D7/EdvK/7cwylLnYJ7E62+GMk1tMhxUhqCRuK+WDSsTgrZm/oQqMuUh2Sduo5DfYZj3sKPo4/Gnj
IAaDziV55ILdvbftPGURi9KqtSL4/u9vvcNy1lkyR4n04amFxRQ3KoV2TviI7wqFR+LU7OG0Voka
2uiFc4YlT5UUEWQokH8f7wyYCGR3dYuo9exZ9kQi+Yobbk4FXZnu0y/VXXrpP+ZTVpURZNscNLAT
iHI87fHyTU1b5Bfjhq5YvGXD7RZ841TY9JgmMnz0T/S5c2od8YiSb8LnVmTaiuYmk+PPLciHw7Qg
PJwNKcYTEgZBwD282OwUNoKk8FsDxMNWyeh8a1nxHfLY7bjFbfRqVjfshg0eN3NETbcwDS/bdOda
2JV5FaU1zKQIf8XwmqVTrLUwB6KVSPvaohpmSC2Dk4YycAhnjEjduTcBeqRPVF6NFHGwgJ2GtkQw
S/Bl1P01Fj/rhDKgoNa14T2NMpDpNmJ6/QFECczDRoVusgzEqMXvlEFWjh8S2waAs17KrkCgQ/vx
sHnZMAPKC7/xENcA105nZT1CP5DLSi3nyKQCPa1Oz2IZqP/b6rh+me5PCtirD+sdg9LWh3EgZZ/2
kts73IrlwPWnW+taSr8Kl1wO5oRGeh0ItUmkC5JnbSx0Zd4ocs8KjEeYgTsYcPHff8yg4ZFLVu61
FFLxaII0PZIPpUxCvZdhHlqhGNQu5e+z3RxYt2XvLinJLHHUrVExpn9uK++XKHkG4pV9UNTkqLbX
a+3rgdYzyArA6ViWNNIaKU/+rYB8nIPamq4p5EybpweTBOjjWOoYoVdVcPshya4C5v+UTkzS6EQY
hp3FOAuhVpYpIFedJqGr/imldFWk5cpCyu9mv4HupDbUjYJarbTj+Aee5HePbP6N1O6n1kr47Dj1
sDD8CXRficpnxMcch/DC9XMxYfuKfd2PnGmjEcCul3235s+V5KkJvUDPjJYpykuv7IIqm0Agxcqx
MeuUtVBQ38pmzG8XpY+K8eGQz3RHkPhUrMewpDNvZ4F/03Uc/9i4RewSxAknoq0dH+isO3fFwV8T
7WxA4Str7443gr/nVuzj1bE8h6JRxbv0jbuXOdfQG/QG8J/O7dvYKITlhkftNIjCpTEmGRcprZMp
ceELCCFVLHv4oiX1IiysdbdKaXjnqJy80Kn4ieTpoi55Et1DM+oSo8IzYj+KspMW3GQviXd5SsGI
/q6Kq5mOrofiHV+x7cOxD158wsTSqnUtEFyGvvsbaTUuMNJ/VNrLyGnLmXeYQkzop447ofPkLaUC
yEWnGIlqDvBjEpAl2phLNufsjC0e4WoGLrAPKUsxgEH2i5j45m9km1brBTEjli3BuoDkoaU8T6/m
oFWXVStTENrjyqEipEZg4ggte3m2NUPQw0ryMJRzY7OUBHSeEOKdhqGIfQQ61uy/rbnNzGVmgzpc
I7D1nXAN8WNKZuoxIJXv6r00RFGiKvzCWTneFUX0kDrsWirlXWnieZ1YzWCq5C2SE5DtcftsMjow
pub1pu4rQaZAKkLNN4LxyVtsxWRwL1xvnPhqFZWZ1JQaT3Sfv4SRJAbL0FxgK22zda2m47GX7suv
AxLTVOg9tUr2/J0Acz6uNY633bMbBzll6TlvvZsbloGE5wHAZJTjUwyZR13sHOFl0GjkzNpAkmHD
gCeNGO2PFAlf255H1F7z5XU1kc5vNhlJhE+BhNPxLr10SPV9Rxg5g264JPxJFMHSQ9N1b2ojusQ1
V01kxY+lA06K04Ew+J15iyWxidVJLEMT21mPID7xGw9WirUjiHBAoUB+t5hvzu5UZPXHEzL9U0Y9
9Ah+bBxXwwYsRwXhxjtdrV+NApR0Bntzs1pYOPbOUZuYOkM950Z5MB6YUPVC9R5bpINHnxLQDIYF
IuG2dZ/RXhyTl8vQcfthftjaRytiUZaxWKny/X1+fKCWcbc0ctKvhD4FrOMZYjkHEfZLaij3aBNf
NDITTT3AawdIfd9pCtbdbV6V7e+Vcacf3Sw6eIU2QIr6VQ97tuKeXy9WG9Q8VrNgfTvX+voMpNG+
gTYnevcwz/gSVV8/3B41JaZGvuyGuLcuzTFLZWzt3ulVy2qDT87/3WVlbRsSo45hblqSojJmHmJV
qd4uvgMRO/Zgw9yS9sJKf6+8m+vqv57EMeVZ1nXD1SqRXUfBzEUCZG5Q6AkmYV3qKGDUZwI3fcJe
8aNl1MKMeHXswBZ8MzDLoap9NUDlTZVukkvraT0Lpnvy3M1cuUZHfmp38+PptAsl2UyslzymdNj2
zNOWmCIAZ2j2/+6gNBgrWSaDCiNdMs3GS1weLr8M5oHILaqX01cYVddJy09Fk7k9tGNBX4QpdnEG
dPco7LjfL4gwGLSojY4WdDJ8ACUZAGBaj4XLufsOy8rOejtp15x54m1I6pCA+G3chxRGDDcbMHau
fSoNeayLa7GydXrEGvFx8Ij2VyB5WVBiK0LRsLIphYEkd58rM6x4OHtCccTL52llgoQKCJVodKn4
H7mQZziUn9MUuBQZ8aDlSgODHrkS0Dl5iR4OPPJgmCEpD8j2lmXUXzHCZRzf7367E3gp+nrdaPPd
rQkaCXInf9Z/GapPk4whOU8lA/NBM5EloDQT4ZKxwOlOcCjWxwzF9nTifOviBCYySn4hCD84RLgS
GgxLo1C/ASuv9fjRjAWNe+m9mGNKS+vVXxdPZGebmmCFUFnAoaDsW5+WYJzjIkMKlBnOLIsjVs4u
xkx2xfblJ1tXtVb0LPrM41Gsruj5Xyo/WaoLUJDX9q6K0DnIxE8u/xnkHcl95WaH8ldBVG6Iz033
Ue1RW84jQ99bxvJ1CAGbdK8U4Vkxz9tlZAEsKH2NEzfvxlVT7QNgvsbWzaTv1qMgCXMeRqaBPi23
bnVi0dL+k0MdyXh8DCHL8FwpYh1GQnBbxhasQ3xj0ubIj6KaTX/OcfLwy5uSzFaJ05ulHIWpCHmc
Y7w7zKz9LVuRR9t6xDWepBreqkAGNfF8x6ov291q9tX26/rC/IWBvhscRa2UBWExkvqhEc/ZvqAt
YOWzwSuncGxNXSLEdWZr92rnEyE+vNyCnnXpwGmSMyAIg633ztm03HLv7DjYMdHInSwxG0XXJAkM
RKEaTo8K/QQxrBMpibA1SRKdF+P+4oNVyva9nuyMmOaC7twiyzT7kIUzpJ6iTMB3gEdXKEPyfR9j
4OUnF7YWhevjmlN4u4+isDwtLXYCS6mMmyo9Fh5suJvzbQNq+0kZrQNskSouBBJ4mcarUUb7oqOG
YMPxzn0ZtWyj719vBKmuYSeRwXwmdSxDZBfEcXr8trw4znMBZdRNDQ9+nSFPChCDszQwSFyo1lsz
MEgk9PfhK9Jh2Ezbuzr2HOx78IVtM3HRC6hSh0M6qjueG4Y/zwwF59vAJAS/StI99zWMorVTIBOv
PogODSfCNuGWb6NKSMfZcznwZgK5q7MVCxDYJnDHkpd8iKcDLi8n9JYz3PbgXhzITr37miBj56ux
C2b8bppe8kALfEliLRmyqUUwlm38fG34aRLL5QPP4JkbJnbd+45DIk5AtCAxXXv+vQeeZnPIwA4l
Ga2j5RoAOX7tZ353OiYDKmred0ZFRyMffsjN/hGSbORPrDa/uWhkDjwYL6C/45pj5wjxJlwYE8jz
J5I9XM32bmw5o2oJOYE1QQc7thBWXGNWSwFLuSCeeBrPqwuMzLZ1bv6c0MPrLV9Y4sMV0Zqv5bOV
IbI5CAq4v59Wc+bwIbEJesAcpTl7KvC0D7LBitQWy8LltQe5OWtPTZf3Ne4gchA/JRFFn7veCLyQ
3Gk4XbC1UZVnOxcmH6Nn9dubocKtJioKTmWO6LRFahjDODfqszmfktE3JRnwInMB7YgZJsleRfD4
U9XD4IeIZKvCA2BW5W22rG0wgpAx1plbWzKnvYl4IC6m40ojXsFGTH3eBS/aQqaT7s8sh4Fa/UYl
mydhBRzNXToSf03WMvZHOU2Bh3UDR2iivphVxfKP8GzGfurTDWpEgkpBaB0xbStgjZf4N4qRgBNc
k58CTvHk4BpPbw/ZB/yw3wSPpTO9hM9o2MYhclg9PCq2N8W/oqOM81/J7w7QmcoU3byFZ/pHSUdE
qOdK9xcOowksSuzzYqurKsv3Ax/xfgWIN+yno450BAlSWw7HKGNxnsraSIU0GouHdO5nRVIPajFO
HF0GlJnKr1ZKFj2V/Utg3SGyeD/+A+jtEiLEjQqAHiwF5qFRKR3N+qY1Que/4ule3Ren7fc2BPq8
nr3RTO0stHIFpriVZpH54SPaBWF50guOnEPBYF+Wg53sMkJjJx6VHWuXnDskFpWOSQ4tmdzjEztz
AcxA6TU/I/I+/huktTsrNos7fV2KrPgojy2j3D5RTq5uulpC/RqggRevW7tH2qI6RX4IKpKigfQX
esjthLrrufTrLPsoLM68HvsdR2WDgJnY2X74VgLRYU3aClGgOgaW8f1207b/3ZIKhtUGvUpZq73i
iN84RSRVGUtQVPxyBk2d7vBZInxI1vfrZv9tNPiOc0F8WWDiQagzo9EgJ8jN2svBpjirUDtsqNIG
95hLf64r/tsjtu5JolWOpC4FHcgzufxX875i3PNBUcz3OBR0ecbNdVgcXUw4GLTaZNSmhjORcmhK
lTSTZwwtssWjS7WUKoZtBFg2IdoGMwc/g2ftyAK2CsVx7tLFeatmurzwbYbePc1HpoFjek+fZo/q
7NeSPiG62fsh357tdu6OFMQt1t4KVrFRDJ6ENpDa+wyl6DkVxCG4xuDGUosphH9Bj37ZT3q6n4hk
yKoffk/+LkEcINo6YvF/bRrC1EexWwQ6Qu9zpBThPi4UouVygGjkN2vfCkydjqg/JOqH4d7BZB7m
DDPwvhymp8PXzHSqQmI6jg0YPMN7MqmHNE5uxmeI9kAeK5nmKuoNed1Qx/l70rJPNyf6NB0DhrQb
vxYYbJV1ZYohySPF6DPfUI3aV437l4G3pLw+F3OmDwRSPhiVijdhy2aQyjoWPvwAw3GoMgENhNea
aVa8xMrlUeoXF9RtQ2DgXwMGYBXpdQup1QgF0DiSr9zbNCWoI1eNV+GHmkJK90wWrW+IB/k3d6KP
exLVKhcjjNzgHa1NqO/UNboWnAk5748gVj0RQzbUtlz9f2SzjCueCedrPBSyw7Hnu3lvf3wAbiEM
h4qW6EQRgoB/mORynncq9G+ZlQ1KAWcmz+Xl11Gl64TY5caJ26BU/AZERIHY5z42SQGCrFX18qTG
1LK/SbNhDF5wNONoJjY7K3JnO9OYwSyQEYB/8cEU92W+MNGxduuv4CfWQrDpQQsdZY8c31jF1ogR
FoTVYdho3SjL2B6LufWmrtnqWxNbEYAp+9+Exxwapop1DwgItDrI3K83SE1c3FjagX5DfemHdPH9
tBRoriqMzzNzkFmviOFCMFDAS+ReW0d6b/qSDf2oHNbXelagD6T1YMLkHy0diQfIvEeqW31/yIj6
O6LYRyVRqhZpfdxExx7Ovb9r+7pHKkRh7+OAG8MHVWvTt+nbr6ZnQQ+SPMOpJVwSfccI1A5ZXzOx
d3ZrqmIpE8PeBe9kg8x5Stn18gm+ZroMagcf7M9zBFsIQDqOk5G2zn/qKfFe92b4jugEt2YORUlb
hbasKtGR2QguARtRPniyZF81YHE7uUXNjNg8JucrmM9zDZBrJ4Gpke+Fpl7Av+hqw5cUfkabxzwj
QmPbMgVTl3ZS6HS2TA7LSSpxiJvd0hGdd4D61jMJ4ttbpPdqlErJ12MeVhHJanphHBFmJDj2GDr1
JySZhI238HXrClOCCXyWyJL7spLO0qKT3dMsA+xf0t/EOdvPpNZKU1apxJa/T5faf/dgnxvMQbBx
bWFjfZXra1Wk4E1aeZY9DHLipIPtEMV1SwHTRcU7AVH887uJwJzHpJ6oPm6i5v40BrbkKAJ6JTeN
hVgbz2QgwMcrnmrJ5PjIcMRVSOy3UpCMmf/MpUzUZlZKkVJH/5rlnOvXfO376JnzCmvlDCioFhGB
jme+LAR7xS+wwec/cCR6L4thn3IM+tTdqiNlv6mtBbB7FQ98efPsbjti3U00hCuMpYIwqgHSiPEN
ULjGvCpksNI/pECqO085Vx6mDuXp9n5OyVaNYj+I48QtFtnovjZ6BgBJA068XxnAZC1CF3yZPKN9
jKexsbqP3/DfNdxnT0DHgAMUTzV1fdd7pfIK0CSTS6Wfl28FKLaLNs751ZinTbXdJH6iYgCgmK/S
dGkEcoiKaXNq4drzJjCuEVWRPna+TqntqOwg0nyAzfJfN66UXAOHLZi0LyIQDokSs70vXf9b3Q7L
UB0CCSrDmjIIFB7fRI1MMjmSvQB76fVbJqwkfO+2KsXxSJaaWVfy2c6cd12UQyK6/ZED3PG1Ocbf
KocURsr5Hc9zliJW8GspsZnJ0MtYeJKJksJfQlxt+bDkNrTmXxAz8UlLFanmodT7ViOgLnmKxkHP
6um/1uwRrA7Y8mLc+I+3+rt3Q8ooJEOE+waf2PTDsWaOeGxpPYLTL2H8+x5c5imld+b4JEEVZtcH
5pfBbRDjpp7VOwCpDSHWeHtCqYFBJJ62cGoQorWy9yroIjMZeDMVzWvu9oPNn1SrpzIG/Hrpj2pp
uUGU5qk+qywBDoBqv4Muad0MU9ut10FjDr8n2btzV4WU4KIuqcAx6noUPN3cCXWMWtTc61JXdEbr
vB09kJTsggdB9MiFTVFfm2Mi0J+HKS+FciFDvWifxoPIwbWjAICChIbLMsQh7ValbGyd3IicnbEG
m7H63ulILnSGfeV/lLUM5V9c2AK0HY4hQG3bjTq7atyohju6OKISCVbDCaUCGGnsZOR3rxbZpAYo
0YBGGBj7ai27QA/F0UAtOG+g30r0mPMJCwMQkVV/YhNXzZ8yFEIeWbmD37dPYwjo7/npkTlUe83f
bHsqJidPOxUee+RA4rn7f/tEIxdZpo4o1bYY/4So6S8bSyuFO8Sw5+23V9KP11s4nPMpcc+6db4m
2cmhXH9oSpSF5gXVAOsZnVLQvWXN4f3XhNrOmg2tJ9Ws7o2md7sdvxh86wVssttnM0l1ZOnm5xMZ
hQPBt1/zlNlRP3iPjFQ4r9AwuQg5S/PwBuDHz4e3RG9yYV5RxdpqLc4hxu5vSw/Ie7ira7jQZK/T
mz2URyDf0FCmNX3Ihi/Q+9v4ERXKl67jJDjD2o3t9WNsIv8KGBwjmhP+DWXfjogj1Qm5DBS19Nic
HFw7dB2cOO26+zn6NcOt6raP/rqsXLahGFQBKgkFdQ4fBi4joatTrjQRaJD7dDgRgYJEy5WX8EpV
ovKMIucR5jR9tmUfan0m3EJ+roD+SGj/Ye3n4E76bDR6R+yEiOKQrhxufX3FJmbmzqxPMciaz/Hz
Tq2PGJRaxbkCxAC33WQeFxNnYfjGMexQQR5upc2mpKXR2GYwL/mKzXXzumVF5PrIukr9t2lOmpfP
Q4WrUCk7R0ZUKiXHCwYIFvaJBLp4nkVcdsgNbW19gtuPWPk+dHb+g2hqs3mwRPv7+ugra09VAuGN
YQk1eu8lXGQt/MWxVZbV+N8nBlxCpsXomSEf6cX2vdamXY7MpFIlm3VYCkvQ21DF1M1VIkK5DTYx
bDaBqCqSIbYlgofxcOU4kEeIJzT+AVNzmvgqU8eUD6zFaIiyun+JX4rgicygH9jDqLwoy28aLJNK
9bhVZqqvV6pc3pTK6QGfnPxFohIGs6uWWHCOcAM6ZaxoXu8Af9ymcIn6SiHbm03VlXvwwHkYnz8q
BxGnrGgDIR8oOZTyuLpv+sVeSUognnUKSjcr53T3Rw377KtNiRsuNiV0K+veC1DVj8zwrjWM78q5
GNhqRnBdrfZ+ebE3N3oJ6guSLj752wiPvJvHm9l2JLVGPWy+dVgdBv0C3jrkSjwBzlbznQGa7R0X
YCfsIqwC1JUEvrZn+0Nr7p4adA80yAkBuTXulmWycdKWlbDRS1TVbqq7fzV8ygUMgs6HGuPHm7qh
xqJTYBCHGgzgaH98XDeyk6qOHvIExBt2MoMc8W7otwnDSjsTuTv4eUxGERnfRdQwjA8FAzrlahm6
vAYoTy0zW5glAIIBVeVX7BJDqCGfe7VjNB5MThNC1LkXJlxuK23np5h3LmcdKhz4+mkS6JVNyTWt
oZFqIYsbSHuUqgjyR99D4qSeYBQrigX8Is7Nz+CEGCgX7Y5wV/0heLpLqwwwWWmazhzBgoDQk3E+
YxGBe+XHRgMXqhXCJjCyUVCcU5aFQSiCRazuGePxtEkLe8lfStrh0GZO3ghhURo7wXnmh3279dYD
DbykkuMa9x8J0ST9TWvHp0UlVXDe7mBfegDsIif7bQlYZMe6rdlpiAeAUX4jOmbkYw1NwZ03bsU3
A8y8UCq0ArXaNJGog/2pIB+P9Vh30QXUFebTWyRZH2FV/OXvrhcd10Bif2dWtCx2UkwArEDYjfbc
ilTIJ9g5j4JHJs5P7C6cq5G5EpgOYs/uXn4ewV/9IDvEPSEY2qlpx7LJbSWqvxo5S1S/36+snJXR
ne4H7DlUxClDqwksq57nAIMV0SmjLWAYo1TOEd4nfVp0TGK8xi0LVXuGp43ol2Sg/w8N28YT9l1w
Bprdmw4bpyWy9JfPg5FIMoRgscEE+j0atFM4ArnDHOUq2Cs8pEjpLO8S3WXEVG+/4x133khEhFvV
0P6r+9lz25HNfTs5r2SUZFmmoNjuHVoon5i0Ya12D76nfqz0idyiTz6B/ac8J7xoWj1CNIE/Rrd2
BVptTW5/1T4sd/P1SSRnfnh2aDN5KnKOSLZmXRVjKnHYE1qoreg+QYTJkK47DYD3CxC6AqivuWnd
qoa1FTo4ymiCIE+KrtPF8tjN9iAF4mlemit3g26LEaFE3qVMVbozB1zojTpiw+546A+C8czCSpk3
Y+7V8ftvTjR78JBz9ZVUU2WlhET0+Eqs39y4khRcRTZtymLH+V7MqYSBL/y4obX/t9dWSF8/HHFW
VGbMPw1tniC8Hl1HvypBVAT6e7/BepX7G5xarPmbpdURlSQWziXD9kAa2FFuDLLbLqMmR+PsNI73
/DBVy96LrqBPsiBpL+sO+kTXHi5NBckXcVRF0DxV2FiE+2w8U/gRaOTY8c1Iibx8srB/xuqORDo/
7qKrE/fnLWvMJ42A1bb8Fq968/ipA2OHnbTODKL0KGMdNmZDiXGxLx4p8URwy1BUrS8Rt68+oeRo
qfSVFcs8i7Ows8UzFS1U6VsQQt6zS2CEislB3i1TQXiiXTdX02nQYwGRvIFoILnbiKtioeUyc0t2
mvYowoSrUnG57uukM5fPallnsOuZyTGfhBIuo+DeXFG+tbDUZSHvJBFB2mpQLc49m1+QyCMpN1s3
tbVmX4g6pGXsClr4O9chljGFHGm2JKpjzFn7QCCZy69Wz3EU2U1pzvtu6hmn4CPbfFJ+RBhKG81F
w8QljK8qMFpw95SIAIUmkuAgfMq7LZ//KUlkSGuWsc/XhuF/M6JKRuqRq9sxu/Hbva6uPTgx5eCE
3ET2YfNGHVysWSWGrJXMMB+h/G+StPoy7XS0hRNWSSjxOU2FPRPU6xOFcj9ARgsutuf8yQGjcTIt
AENQsI2995593rFKPUSH9t8OVQuGw/+kzRlYUV3Qe1rKx1q5fb3pRAtm8lIMCx943g2p/IOaky3K
nX5WR62xGu6zSYocYSjKPwaC1fO541AvdouH4OilA0dtCJZAWexWlVNes4I5YCrAzEUJhym8ngbE
wqEpA1BJUvwOcfBG9JzDznW9btcVOewvm3fprjgB5LyQFQYnfHqqmzWbBAwa0OCc5+2307zCDMze
8wm7ROgX7S9HJCWKjWRvJ4KsVrg9hhHfr8PuHHIlcWfTIAcMykuqFqPDNEvXplhSxVC0D7mZSLsQ
QQVXw98lGfz0/MMLr3zLbig8bUGVCuIt9/xxYnbMQHxi+m/EggIjbnJv72S/zoV7rloIiF6LHZGA
mJEkNpoQA/8Ynzd49iw8tAXQwUMzaiFcCJCs9lZL24ZBRXjp8I0EKzIozqjy6D7JrNxrtGuIB//T
SNbo9o2CaSRvVeDdOVm09TzMxRyTc56DK0kxvCmrkRLAv/AprGh/dsgM7xz6nyZd8ZlmScMjoPH6
xcWx2Wm7Otpyx0211yFCh/BlFcF07BOC2taynzFK8QJshqlnenFLR0vQAGHHYrn2UH1rQ67zsC2I
OlxuC/w91H6cgRiC9PnROOMzsykTlZH3E0olrukQyqek9qIEksn/DIerqEXd1utimW0xErjZRsIE
GCqQoUm4v0zSkLFgwsJJlQpGNiLWIITWF8geMn15/1LKOFunnipTwWdBHbb9CLhT3nlPIOsHUiJ2
Z6p6koyb/BnD1Nk7uOm2LV1fc/ANtpoqcRX8ye/9B5SFgCq3ORjC6zoF2Nyj0bDL81n61WrZdKJK
jmEa6hhQgQ1ir0+ObhzbhT3c11K/a/Zwhd1G8oFj5+1rsKX10O26qhp/ItE93SRnlhXYYPzYQN9F
6XswH4jTy6fPKjFEwobTQXvYoZGY5UURPMJ5X/i+DLuiCsp/eICgJfmUk6PDbt8DPk0f6ImFmy8K
Xz0MZPc2YfjJNYvigE3NvZ+UPiR8cLwx/H2QK3JgDo11EHHr2DaVfFKcEi4k1RlXsqllwEqnan3k
8fJPbKXe9UT6DVPKWLETCm59aC2EsG4G/5Fju1Nv3zpnafTaxdCj6Zo2zV3i+HV5y7X2g7u4Wow9
WFYo2qeoSPm0xfCSutYWchh1GZwq5l3XahsAF6qhfLx+IlWjhs6v+Ud1Dc/F7Yy3y8lO85+NmR+x
cyu/fByHEOmKrcSyZWxCDW1g8CyDDErUn2UMR4EcPF79nOz8I8Id6uNUM+Vb4ZUVkSG5z10BIvzf
cfsynkkwf4X0669gO5wTvdfGYs0jN+iPNWAyDZzF/a2FaNQBRYBrsIfvOQGNIxVkmsMtjJ7C9tBR
mCtWvXQFnFjjbJZRlcQoBGszI5c6MFYtlGFBYqWaKZLhnaWdRBurNGGajZuH2YT0ua+vbIMrIHIj
rq/wsHS3OOo6b2jeDkwTyX57Ug0JPn/oA1xpiwKgJ8Ty/VuGeD6R4eQaVmFa+rrlq11tXBsqaOb2
U0GWJzGD1X+cTh6L3DiKdjW4U/sdpgKjE5hkNdRwHlvevbP4W32blxpHdfmLJX4+MkthWAaJq+Ol
b+gOzJTfwsJYRQAjz36rnGyP/kKwa+MEhn9N+g61ZvoBDnfOGS4x4PpD9jmm8BduC1of/smpruxA
oEejz900uI1eV6cjBkYgPhyWoAMXsdPZrHltpORABdhDDUgGrEKL6VrfmOlPDdyxrule6oZd8MD5
PwKdcDtfpkmL8H8EhrAwYv4WA3F3r7v/AP27eruhV+xzalOwEcXATAA4+KxddvAvuRvhhWT5eBS7
Yld2p4kyfpqmdOynAaV+y0lr4m/QM6HvaZA9ViP7HxDfAGw8d2jJVgeRI8dGNBTv8sMI0+NWAAg9
uDL1Ulf6zw30N6hPzXnl5cZYFZ8Sh7s3g29RC0oyUzqkLlFPcBTJx8liZeOPhGzIRNt649w2rMlY
9z10gBxLTx0jcQQq0EqEMldkWaSyKAoJ4mut5SYRuEaP21vbPxFlvHx1H1jK40J4t3QInvycncKq
90c/YYYOJOqCUIshAwDBMiGwJpsg60ALA9tX1tYSFEe+fGfnYTPg3BgI3t5UIt0Lshw8DS+DseuU
tQyH1bVS1L3rTupIx3/uHOXcW12sOla+qYzRFhXJxUTIxlpxgP6EbqIAQTpfyg+Ph5M8wXmfgTkW
M/DxF+pBBmc/4GPH3aLew9BfxHzTQDdxwr0Z3IQqHwPUeEPtks000ADpSqlbwrN+8FjqslS4Pf5r
id4/ULXrMuCrZ/uE3IVU6hs9ha/2MqrlWFdn0AwUF1/y05o/VFUdQqW1vmL5Gv9NPgbSy+5bdJ+A
IM21Xr6RcreOoNV2g5BTsAOYGibQHlOzyQ+oDiDFwhNEAq7lJTa+2scvfa4g1DAhSuPcPvrVf1TS
01dk6njIK2f+NSZRrZVMqYyviqT1cdIAeCt5QbcnWdjZkpIQdY28xV4mWfs5LeeippIhmOyRRkdu
fl4NedqFvRyjLXAFVtdCF5ZWzBtD98Dv/uxv9L4UDdp2loKjcsUQXw1SBVQXEbbbtrzs7ZS1e4dv
qdRwYBpzAak/tkVb39H/b1PcmpF3KUwip0JQwg5vNNxyOuzVBLqZPFpX7ccdtALGX+KIdb1QrwRL
GwekEwXkhJv0etefvfcBbLA3RYqGLGQLp2VRL3PofxTZufjMalg8s57AQhQlNT9w+kaTeSNSZFf7
K8yOuRaljKjSzbtNbzrUuv7wcrilt+BQZc3nC4PS0QqNjCDcucyUYFJPbFGeTU/Ffk4+lMK31ycl
KU+e1zG1gRhJy9abbq7jf9zS0C2QnDrwCWiP18VVA/ninOiItbu/YjkFzRiPz+R9lbS8kWauFv1o
pkGDLhws/L79MHT/BIkitDy74GogUZ3d7EH0+3QukSvSF9rFJwegkoGGAx62kY4mpm2/ikshPZP4
MCfWxqplCQ4MFKOpThpTQlCMRTyVy2uKNL7c+mvzftbNZ4+UcK089JnwtmUEO+l7XwlgHO/LW+ms
543yA4Syg39Qw5PzINi04RZZgK0NDxOm0PxXKMJt1QlmJJ+xq2Sa1fmJJ7kvoLBNV0LzvoHcmmwV
fpw/4oCCPIKRO4f/C7dR5yuCu0oenFvhPpRqdQQGwCbYqPRhHHZfr4c9B6xbpIPCRQ00Tlcmektj
C/bSnb2m8lbm0ILR7OfuhaGlo+6KSjeNJY53SCisSWunUp5CZoryOKS+LWu47ushVbwdYKkQjhoG
wgm8LnrA56kZ24mgQt2HPLsSOlynEHE2xhMfhBeXBf3+uW5dymoeaaIrkqxOnqrvRfWhDfYXTx7q
3/hmOtrU3CztqYhtSlicOQbof//eJm+SWkYW0B9BQMYNvt6f953aGNETsrlV5G6V9j1357jBa+Jg
kXDFk0lGLbrC75/NTUEO98GlRneQl/iKalrz+BrB6mD9a0akoqBNWDzJK+4gS3MPF30jvnQITOdk
TXfuhig1aFN1PoEwENHmwrzC5oJ3e7jo/6mBcuI+0wiGWMrLvKAiRIsWJ2EFqCA0vREuwuqfmnPm
k73yQYLJGHd7hdZVvqZ8kXy1a2i+g/KfO4bAlbhOpvW217SwFMJ3GaiGYl+c8g8e6YwQatdAMasB
eB61GJL+7tTqr8D+JB87pZI/AdGuoplW7xHP3PS2ZyEBvIzPug+tgpGm3/conCy28rK4WkzqhyrB
KmAUcKVXiEbx4aHA78UqlJVn5gE6q9h5LAqAcBLLc5IUuSEP8OiCMmHuVr+usQunNDkIR51Plbdj
B6lzAsB9mqpOnmUx3Qdb1u+aw7Tsi1LgrPpp4FNzaYXNT2Y5Y/XubmuDXpJOQxb96wkAZvfo8nQo
OMEBITcG25Guaj1dlaHYkIZ2+YXp/4947pNUKuFNazKk/3CRARJn1e7KIaZkUjg0wUbhOaUV7krT
1//WJ9eNJy6BnjND09/LGOoLL+74BLpTC5yFl3Clxv2RflsVef8Qj0/WfMSg2vGxccYVAHisIN0O
cdzs0kYj+tgOB89fE5E/sT6JiPxMfChiVBaisberZyaC0TNtF/0LORS+qvyh0HMNa2ykMtWieBLI
ZNcp5+/JITZ3g8DJdZxz1lrBbvmVZSyTrl3BcjMRRB4jXMkcah326CAMKrO9XclVXniFKTWJUuu3
NeQWDG73eThJqWl7+PJhb2+HoS4/u5i/SuR0WmPltXIAUUiQg7dAYGNIqcjUPY83kIGyw+nJFErt
cuBx7lScRRBQ0hutiLFfiz0m0AV1faBbwhWu4BxKqaDgSqINrPQVNZVnyX/5IB/MmGBg9SPfg8GF
G1TU1DtNHUej4Z/o8pDHgk6SDM2ICplDVVulnl6vycfhZE5hPMhaMcTUQpFLfcgdojFDXRezdLkO
IF6Y4H+tfcToBPZBnhgSCTP3geFqaoxxBs7izAwjmfUy3i3cJc66Vl0xT0AwBJf+rcC9RzgaTpAc
SPV7mJrr69cp4jkhYI0pd7eQzY1GAus/D+tsXAyh0sFen5dpLp9CRn69uMBZqmDgiyAL4lNGvfdv
puRMlHMlAuzo42YHF6QDjhdP1405V/s3p3Af/F6DqGW6Pu4+aMT48f5/kSfJj43UhbWgNojQFAx1
QO+zze2MjeQApZ+7q8OvEhp1VdCuV2lYUQ6YOZoiXKd0JdYuid4hw2Y/V9SpodLCPanyWZsbPTS3
koT3rHAgUjByycTnuwad9o+J3v1LLh/5vYXlzQZwbNCYJZSXrK/7wApDxszBgk8oFfXcU3tXUy4p
bfKaQ2KHjBIXyI4RUx93LbX20dXsO31inn2fQQhd7j54XEZyOh3D1rSyhTHA95lcHXQA4lckkyjg
peWQe+WnW80Jwypf+3bB/kFwmf0rowMOYKFbmhF9YchCLVvozKyGM5CzXjn84w4rGxhoFBgNZwZN
dUpStU/6Etj8h94bw2OZXNOVexFZzI3jaAE8zAhX68NsELEEy+eET/ToZY0X24HMaWPfa3Gnz1jp
0FBgI6rd97gdOAvnGKbxyY4TAp6tawWMF7+QRKmIt+THrHgVC3SVtcUxWaaO/cBAQ9mpfiN6eNGX
e8PZ6w8uE3vrpRnqIHZnD+0qag4HS6iZy7HBhC3GDPPEMm8raFOkYJFMij3Q/thrp1rnBlNF8lj/
1u0LWgjFaRz6XZAkQ4FftMUzjTmX8C2sxlGVUkqA1Ni+poodHieNkqrFyrrogw6UqTeYpWCP0+eU
cP1wE47mUwbujjSPDpaZkmmmcRUcCfAVI5L9MCk3i/nOLRnQgoX0A7NoeyEWujrQUfpkhn/MC9F8
AmRtebEBz6r3m1Aw82Swja79zLDeH8FA4zk2OChdKPJCbhy0SZ2WAPoDQbfR6uW4Xt0CUu3vaT2m
djUxfaPyQmvHMrUbwudvC4ktNWKkfdZ5sLVcJAEMHeF0XI88zR/Kn+TTPYGLcNdOcudHpkcYQHkT
nbepxEsh9bsAvx1o71ZNSyHvY+Vg8PVfmbl/Nq5RZQu8xbw4ZGpQX/t9beSooSypgTTVMy54N7fK
i1sIJ8obZ4kaWAjYGzpMubJQNOPFF4ucomoXskMabtPURbhv5amX5R80kDkIobrdvwQp9mEPeMxT
ODetSQ4hJfRBOOPw7QCg6WaHsETN3oWm1ZzRG8mPtL9JKqwsZCsQvXh2330MOFIChBYdFgKh6W3P
Zs18gc7x+x7K3MvkIy7LeBFy9Pq7RNtx2wFLA8P0c0Mvq8UeCnmQMNcatATHZ3pz67QajD+I0rEF
zzzXWKEtAq+q+r7I2mBAl6w/rPNOMulYIV3PyiOZQT5Uo1zSqqp6P7gaeCjs7dgKBzE1XqbXkiUU
qfCJIL/T8gjud+8tbSNDhMwYOi5jg54VQou5ygC+6wyyTbfOpYJ7cbawvQeTWsGap1JVqyk8Zc2q
bqGu+Wjp33Sw0Eu44vljZjsqxvo1QquALjaV/x2ELDi4qMyT04FWFihgpbIMkRcdwoMaRoa1taH9
MSYvf0O3vZN1MRaiNcu7qoqW35/TBtLaltS3C36umARDZdoRvlsJVzydOnnCFh0mhnylFM/UUZRc
bqnm0XVyL2BvaX+kV5PA9+A/TW+P3dWBSodnX1EVCtBs2omKTqlRuNT8kIFvHwjijzaxBq8/eVMw
bCBz7cIS0geQPE964KWFa9vpvEjGdgYz4xEkfHHgyNhqeQ+V1aVYWdnKHRPS1RC3madIEtCsMInL
3VT7Vaywq0kpMbjd1LrxVcHFrL03CbeFGigIwUshTtJxfgA7I7uZUp/J3anUOzLcKBCoGp2IVw30
KWRIhxwiBtrIXOZrRXuBI44CN9MsuRpikTBG23k5f/oNFCvCVtvOft/A5bXJn+nRbgW/aCw3HB3I
ionhdxocOajOS7a0VrSXakPNSpAiQsQUWjecxtA2VnNWtJWHo5yb++QhBskTHHEowLxqI7zn1vIl
MxX+Gy2dX8JoV1ICUfPnstjh4UURR6n0s97o1/YkhtB0/OWcTYS4I253spKsiF1wOQHWbsZjTol/
WyX5H5YQtW71C/L6bCxrG3OkmDHqCp/XjuDyN6CRyq4nUnMqDlKR0fSXH79KCLFrAjTnh53Agcqt
A+mPWtzpUVICS8t5n1auzJO3xUD8pbhQr6AP/fwGbRVHEXgplnucWxK/LnmM/Gl7MBdNh2JhGW3j
0AhuQuAfs+GbLbqmuKarwCoJaQauQLWR5tZuEyz6dGMWlXlAfPLahdq+6nPn00IJkqkZL3E5eQtP
mpL48zN2q6SBjVei/+SgQg5BOgtbS328t23j/u3bUAXykvrsWhfi8M7lES7D02NLlErAS/0djMwh
iev+gUgcxlX6g4hSoytmxioeY6Sx9MrkJoZ5OG+IKkRa32+zhyZFWzXGcin2CPTGSTZsTZE98zdq
pktaTL7i964JWKp+sPwSVyU5fxPlbTdJo5UfHRvEs2+226ImacbeH/AiJ8rkNT0vHaaqqaw0JyrH
YcyCiCXJiqcoZDjASNJc9sw5o0lKgDChIeNL2ecASRCo2xVkDhOAh0v0+3K6Vqwm/p3InWhuNCFw
z9VdkLkrEcMqueCjJNJRLw4WfF4HtoVOzeP4I9dBu+KqOC14D2IOP2bGHEeqIfM83UM2ChMYm8JA
tBNMr5QOtXnr52eEhjw6pBs3RJcA55N9LCfFEAegRA8yH2ZvO/czDhNRM7tTwsAnhw13cZG2LvoV
t3wHv/pV+aLFulWhxl2iXmucontIMtJXKigPcrUAqSPoD7+tl4C4O/t4+1r3v/rEWy7Zpq54rGWa
inL+SuKEYVYGGk1q3EgAWSN6Woi+wm4M+ghJF5WCjFGzE30tVGDpOdabf2aJBMc5IAt8YozpSXg0
Ueye+/UNWw5WFMBfIKBv3BnTGF/ezLOTrpZCqIui+s51XwqxfE/h61pAjyBYqcUQu722N3IfhUKw
xv/KWQPlK0emWdw9SQm+BPGuivD4jbwgbsUyd/rCENFFuuqnNwPyh5LzVn9wMVGgLEJwPzg5MXih
in+OXkXUCPMEFeiSJTcv3aposEtL5+5VWglZusqm4kBQlmPK03W6bdLtzysOzXgOzn3iOTNf3hFf
eWw4NECKqyZbI3TpUBO0bzENFs7yUyFIudIF1btS+fPVq9WURYi4OAsBnO2RVY4rc/R8qlaPMvyc
nx0OUzJeHVMGGOTwydGMLE7WnUEfTlal4CgNL5xyeuk466HmN+f7jhxX7gJYDFdzEISoVj+JUbhy
0V5RdQHgS1PHv6vkrZ6H0cLIWmXT/Jtp86MeWOQNIbHMI9v3ffRaleKtN4m/5ohLomUv040ETtej
puqkN0QYA0MUb0mwgXK33db4QyI+5TOnQh+JWGrjH4YNSLubhMOXwrpml1fTpdwTopl1GJIyko3I
exv6jDri0c1IyxbQprvuFyERZsXTn4nVLEneh9GbJk4Ezi1YtH0ynDw/E2Qtjh82nPuED+b+WKL7
DIajCqbWy38h922YBrxJtx25g2kCuuWWFCHGjn0ZM3pl9XUEDywQ0i4mpcmlYLkfcvqdvGFPTMSN
71A36oS7OcOnRCTXffRQm3tKcTK+8Ck3CKgUyAGmKDa2ptQC0JGOAzjQJlCImo0Tgqg/MY3iuD6m
EMAf4U7r4V0fzmSXRTj/O0+nCufeQ6KXifI9QGOCciPWeXWpy38Pii4faLcazSk086S0irv2PwM+
GP/FAlM4waUpV2VBpc/snHt15JXnFCWNdEBf7P9+rGhw7l3XOgxKLoeTfHzdMTGnrsqnINlUmsWR
opQrXssJ1Ny3qVOO1yDsaYJMPZJL5lF8STbh3d+/Vn1PK6P5Rkt4C953jZu15ClJB+45dJ4kH7Jo
FOdW+oDynocC3Ut6zI+guAlXLadgdT0Z+s21FtCsiXxPnkR7wyCu+itJBIx6T7kAYJirHAiJLWMF
OAsaAyP8r4iMHIjLJhtylWNdSxUAZTh+PCD9+Eg6xaczbkiQ7XFWFZB7hiNwEFLd6Efxf636mCA5
PrG3KYCJpJc8+ccmICX7N3+9bkjo8+qMTGkiSyoMbpZALjvUM8XJZ1Dc0EEL5+b891WRsn0iDgLi
6J5g56Se2gadQF1tz68JuO/CLxgFr8DTAyGHtTx+PoLdQNlu058DJCA9o6SpKd3eaqcgkacGpIfK
bm+R2waR9BR6z7f2m8rT04KuB7oUZmC88jvsL3mOlX5qjzs3jNDyZPbS3qgZnPyH4iJYvYq3QgHi
D0OiBpWozyVYwy3MS06R09cqK73o5zr5xkBofXy7vNzSEpdBBUMgSM1V+/yXuUag3VUYL11LyI5+
n2+x4xUdWh4DotdE5eJ2CTFR4sZP9h8IaHA/dQ4cMdThtQ/4UXvSMSyMy9rbG4th7lDzBeEOcEIY
B1BfuffAmKXNqC5n6Cx/P8Mm3FoNb0g++HHiCICpe/HPnbNay4NhZ+rLxzpxPVSVmdW4J6KnokIg
P/SyufI8JRyOSqm2DppoeKl1cPaAlNZyBNxDI9DwCmnCGHzVS7L5VtGkqgrQWZbr+MDFFaKMxIOM
aQD5FIBFaMmFrBzHr6H3ZfTPaxdIqvgI6H/oL7ORRMTjfvOqWR6tHJgqoYJ5z6xZLYfLIIafeU0d
cvqWedFJIkh1dDSn7YItkJ38yr623/nNefDXOkzgw+Kakd2ch3cDyvIqoegQYrletKCfCdqlUmrg
/UrfG0DLbre8F17UI0iP/9fJiP2CDmP0cFPaM0ASFSce1dGdYU4kN2T3Qyj7Y9wKdEvPzYqMfSAL
45RGzLBGnBJGpa9RgdeEp7cp5ViMJ0vrKyG5Enkx9B8GqQiFRsfPw8qqmGMrNNadNqRx4aKPxBQ8
waJqx23IO60TLVDSrLJvLtT0z8EUjGqBRovuEzROApgMeffDNrVUqnyNVcQiT+f8EkpMoU1sDdKm
cdjyFUpemtTZJ+2xrkigkRTWbuFlQhQ3uvvlye4QCoSw44qFomEwNRgOjF4VRgl+3kULkP7+pHyl
YwBL/w4lE5ddwpr0123ZgQWjE6jJGmKSbyRB4X9x8ir0dbPXu87LdpjYuT6SdPLeafYxBwZAR8BQ
BkWlpyVTWQbNdWTbfFUmC2On864pknO/3ZmGtGU+70WTe3GU8hv1gTmpp4F5NCp8WQMpWzOGdZtZ
HcipcxXyOC46ho9rpT2UMKLfTTjjiGnBBYCZo8Hv23gcC0Q3cudbRR/1BnRzctJXcJQZ2tQAGji4
TIN1d64zpmKZE9zjY6LcH8XMVmpe9gKvSjeZyuKDhnTIe8OHItI+rX91/1gK6DSa5UPezr7AB/gm
LgSEhA0EV++OLwRl0dFlr5d+n7qPlJsNXAMhVqTYLM66+UAnrfejtjIFTxJ47jQD9K+LFUcsuH/b
obD8VMfmLWc7o2ckT3IKu86Fc7bOVbCbVZ8FlE/TGMQowoerx2FoQyQaeIMjNTNn739w/m/bjRGx
27FzkuAW4WtuJD42dKhTsdpk/TNYaAZHWgdric5UZmo44Y6GquZflcsiSylrJ12+SR0JBxlMcj8s
6zLbnLHblyDREEI5txtCYHJiA2a6fqqhunLL0zfAuzNyvyRg8rkYHWiLL/HCjp0WCQHRMdo9o7Pq
rnvvtKTuQssxtTr2WcoepN00D5vMJ47XxNWOIuNbObUtkTpraX93OfA0mcd1vaKfIqyBjPfUfNln
660ZJBgfvi2IRYXckQx6B2MRWP2Kq3YyiwXHPuCFKL8ny2/rHEpoBSqsO8w4cfGY2Ob67+qC9QNy
BzfWIf4zoo5fy1LwgdR3tTFMgb4cvl0LLB0NYcLuWYVV4Uza6AUPOA31VZDD1IK9qAFYqKCLmxFf
2Ka+IZCEeAjnFsibuqzm0PahoJDLJ4bE8azw4jbLnwKGUhcS/lXRhMedTID8mtoKlL/u1ULZE1h8
gTAiyvfvFVvmoFkpxMiM3O5yKBp0GbVMB6qfOf74dn2mwUcOd927bgZe0QIRF0wwCjsnuVCXwEUJ
P5HTbnsi1vTBW/0ZwmhaTBzacqTRVkn2FmC+SplOYyqy/BTIovGAsuNQFKRGbzyFTHVqP0dd+T8J
bAm2S7NrfbU9EjV6Zg8kH7x/N5L4NbxfU3zZKggxOB2mew3TfWph2RHPqAAkQ6gqgBJ8DNLbqEhx
RbaT5iMn5AxtN0L8lww8VHDVKdZqqquK3hGu4u/dcJN/HrVv0cRMnofV8WNXLIYEcbOidFHqplZi
SU+zNDHVqehgQKyZaoNtdZu87YiO/oC5gS83gVYJb3fgX6eeWUwrHIkDF5e5/UUNftvnkCtIBG7W
LdsT0v7Z2aClGqzV50Ri7thn3NdTOKk4QF5qma5SBfwV/XbIAywwiK/qY72SDDjLFPIl9N52PPYF
UGCuEkSjPYbRSPNQ64Us4Qwtl5xxJl/cS6qFdMDanC8mx4CyqNxB0l9DKWybIkjIfY1hjMd0nqbm
b8gClRrRzEEolI48Xfebf6adGhA/U1y2Y+XBXo+ajYxC0SXFLFQ0jz71EAp6PEbkbjc0U/+bf4nv
8jBNO4y0iM6bTwNkCwCqU4a1DTQM+AeQNrZqMsAkXGyRGknTDisraT3x8cViJzkSnn+ZweYWiYCB
ykZbel17ZyLvNRg6tDdVjjwpHxaW1J7KERUHS/jpTcsCS/rlJCDR45Ni0J1o0RowqixpBz3Ksqiq
C2t6T9AL4LE3yNKWkXKsQ9cn6EfwIgzIy6LYH8MUGdOrdpJI7PiAqX2Sj4InN0Ks+TfN5/jd29f2
Yi3gjn99MhDPZy7GYTd49z2CA2v+g4JuWABiMIWzQduOp2TpNU6Q/BSwEPL6WB2gp8A0s/YY7Ebp
3rdiSbLbeQxJfwK6Akznip+vUD08xUq8F6NnuSIywlH7XX00HCdcwA1nUuxn2O9RZ8828JGoUNF6
+H1tr8bts5tkbxSxHWiU1zpZeGrOfyq1ceysancjao5dTMIaKmknaOqlRV6i4KUsfhcB2NREJmEx
rHnaIlm5vFmKNDW+DcTx9zkL4MYVTF3T/wirtY1edprRC/MX82hFOmDySM4T0tpXzbqYVS8DeQm8
bVS7p8fRrxzeVXL8CbFRVQwU8XugRieUUuaP2W2fYZbjOLXgcbtcE0E0bbLV9OCq/SEG1HmYzFMh
GGeIwG3hrzUc+jc8w3+yHl9g4oDHUWRVrCd5kJJyh0NmexLYBMM4/Pq6TUwj912HFIwSb/Y+QzaX
2NhPHE18cDCMWeDcxGOq/nO2j9CIm3g1cgtPOOHkc0nDB/SBxlaUrr5GDLLhCqr027TCU1PPhs7G
uIxRwVmoP8vipk8C4KN2n9+fhIBcuS8SEmhmaPUbJlXEJkhCmG88+scCxG6kV64NhiwGPEq+khNT
r/91YHosDH/79ItFYqgkOVgeqnwcibwzAUBEovs+k3wlml3qJs7ICIRGqpJa7b8meZQG621hDvLA
IJZytDHoW4y6HLszPzeyiIrzxjAItcWXHmn7AJoDtCKqAkd55cUfKIs7RzKNb3Do3U+76Udd+clx
Cl3dS0buDR4JF3M1Ie0zHr1M1opKw6Gb4dWGZ2giT7Xn2U/T2aOoqhJUEcgrhkdkq7tuiOmdd8Pk
FQqHuhAq6Z7/kcRGdXxcHmh70Asvof1RYlWqWLMSbYI8pMGj0auWW/yjYhRIvpKriHVSd+9fjsuf
FhAu6z8TsZ1ZSq9ja8lBSahlm+WrY4WvK5Vc8Oi6q+E7vx9+c986kABeiJKQHGKnh1y+JmhFdwj4
f7Lbmasf+Jfcx4qUfqa7xJ1EhbnRO5rGVe+ozbuYVVNQdWH5ZnToik53nwsA6h6SoDCK1F6OIfUg
AmCfF+QWo13tV6Bu+fB096JoMh8/oRTC3Msi2AfeY3nN9JGJKqPQ+4HSx9e5UyQ31F8x9B3sVejy
Hzbb8qDS0q1s8VGkXufDpqhF8c5W9K2kZxVvE7a0U4FqgnNa1765UZQL0vO+NhTLp4a5i3IP1/kP
e4PnQNEQ3pWqj0dOOuZVOlYOf7+qXS+saTBjAxrtMIdXIg4PEq8WPdA8P43Qqq+EtaG69L9iWybo
7Gw3TxoCAOSNcshOdmfNiZ1wyRyd3LzQAl/3vI3Gai7PD75Mcokh970yTVZEH+Nvv1Ph1kJHe7Ly
V7umoJfR9TRZMkP1hGt6EZlKViP3+tc8HFl2EXocgBd6tGseEaaSRM67JfPI90qAFz+0nKZuqjAc
6Tl63f26hkIMQLAYiPcpPUACRi8Iz1yLWpgXL5NMbZoT9gPVT+ZB6U/A9ciwYxbm7tBRnGJFs9I/
om1iw9lgTBpLn4p2mWOoxL8WWhqNEDsEmbDMgPgkQWBWHix/8ZApyfPOcKd30kyEt7l9+q6tq1TO
QFdghi/NPB0Pbz6UtIXbbGsR6pWB7PWYMu74+iD3mThDytSVPkK/Xe0rRJx3edn8aGIbjYBK2r8v
0Fsb3pxKqdDwkLVJhhIql1+TfGioPAx5fk9P/aUqcUpkD27WldN9alvwgaiOE3MFSuYBB0F6qUT8
cDITI82oPD9lvvU4ZivL0zAK8JSJh9KkdKC3Q++WCF83Rv7MNO7z5/DTSYigJcHYZTEomLmQqaPG
5Ju28r5o9QN6KHKCKu0pthNPVJTYEyND4t3n8pgUyblWQVA8PLd6XVLVptRN8A2m9oclfs7fiYNE
+91Khra/Jf+Gr1SqDDtXLxtiFWoTwYq0950K8A7x0m3MEAZ9mUBSI0b54A64KgIYN4MNlKw7HkzV
58evK1Y4g3ew7Q202CxRvAD9jrRz8pQx0hW89Cj/r69tQQmkepdM83P0eCg3qRmldYRQ7eJpPHYP
7pdtDQGcaki0Hc1ai4SaCVPBYhMdADCd0sgTP6rlnjf5quKGlaXbh6UnqSCiXcE8Lq+Fue/9WxMk
BjdTT5sfVWLR0IBzJhqF0XfmjMy8WXGQimpe4fQhE8F0kcFZ+zsvFgNCLzBKftJMUnbBgNr5s6Jy
DXCAOyhXNnYD3STLXescnjq8QZdUcakSWExYftNHBz8CAz5LSBTo8ZyENIObEIHoOSB8kDkWhutX
LDVWyvPYTEFsQmvxLIARVf833v0e6Y5PRoqItq8itu18o6GQzfqGIH+VhnSYq0lByN/Pxe5A34ql
0MvaRmcvr+Dyzpkfk50ttV49rdBW3mz7s24W/x8tJvdOa0SsL9gOV4K06hBdL2qAtwnQ+yU5kaDc
AjgtJgWMoKq7zwvzlQbqkFEzz674JwLz+3m6nxromlqRp20jCZDbFcgbViz4vkOqntnWm/JjyD6D
v6JQuxWLVCtNI1d6I9W154f4usD+WcVu92nkbUKjkgcVlGQgTWZHADkZVOh8cEcQFnBQBgANmBbu
ll8k/VxH/qodEZDopecGtLMgSyWHq11BRoEk2RjYR6nvgZ5brDzZARpDORuzA7eG6knHp1rQ2K0O
dL56JZQYa0zCn0pkNpWTA7w23uQ3LYkY+VxKJ6G1kVsfHCfWt3JTVxfySlitwQDb+GH10s5BZT2D
gH0q3glRTOeV6XqWAdf8XCh3oMw/vSo87KD2Ek/mW/DZ+qZmlr1yHhdlYFDdUrTx+yWDJgpVG1K5
au43rUaCOwsyqPbF05M/QHOGkMkVNdmv8Xzh9HhxL4INueDH6SVX4/mAwZGkRgFVg0UgZR3g3lDT
mvrwi7XXtgbjn2cAsg1ayiLaGcl2+cMMJHqEX5McWabjUGqc7fYKKP5cluiBfFPHv/idjYZIKwVz
ET7NdxatFN8nBQnI9dtHaVXPJg7QU03uRXt3IRBo7xTSK61VzUo+Vb1ID+fxMLx57hC7dTNSTcg6
/iiRkCxqpn5HucBiHHkdt5rKHsTQqQHIPyg2bOujA9CzaBJl15j1gs1389bC8uRftRMZrL5JzRoV
rj7D04pwv+HOKkVIQLKjqhmN5a18kS5CI9wEdqVhDFH44Ajww5BtWFnAZoC8GAhc3XEJ1K50L45Y
0eUtLRbN9nmSplVj0VLx6MHpK9FDqHPQiWw3QeSzyy2hgyRKVidOO0uNLMwE2iCPLAuD++D0Q9+1
4QjJiLUj5zn26r7nutBDh80mPgAhJchvt55Ul+/M1wrsR5BXlR+q7fOhI5bSNElMsEleId7VZpRt
Tn3B3+iEBEp3KlwWVTsQ1nB5Ov/wCOltFVc+yTJU8IeZABuekR5ylE/pF7AXsG4ve4I319wnm1su
vu4ZJ+oD8Im5rmOc0h0zqLlj+x6KkUggd2yQ37EfuHyzcVrRmpTguAt0dQoP/NxZ00elDvN6JOEL
dT2kXkKouGM5CFEArifsxqxPnNj37CHGXO2Y+hUHkCOdnlM76F8+AezqsbvlUlUQNGA3poy5SeJB
e804tIHINtDd8mqjBzWvBSo0c5wCW6j0KtpVMttFefrWM2MPm+drh/G2jNlI7dgdo7zu+Ohhl532
QT1BIIPkq0yW2sA2bFFHIHfgeZu2uFNot+wM/A0nmlyMPMLmB2hhCzRZWWfr03HSGrY/8Q6cAKtN
7LeU8qc1iR2m+S4ib2roRrsnRoeOAsQgJJafvKp6jUQYtnKyoqAggOuxpybtmptORT63ue0PIQ76
Tw68rCZBd9SYbsgbfuZQ8vimr+/vaUl0u7MsRRGYQKc84hNuvf+ad8XhXOsXiWHAynpUkby7Z7Ar
7J1liGAbMYtVFhl7tq1+RPDD4H0ztferWdvC14XYtpwead3uzw48pKKuW7X68Um8Zt9rX+FnFCvL
TyW4OU7erJZyvSO6PB+uvKyUKwma7NoFLgxy11OFUrRagCaieTOscscK12BPFl5eBCkaAYGhPlfB
RY7HdDwukY+kAjw4jqOQE/q1mqFDZxIXQ9lZFC7d6q0TjQgHrZaEmWPC0p3mpHoYoNz9Sn0UfNnZ
tAbdeXjLxgMcHjde0r+S7TYUhi1R3TmI+oBI6d0W0QaHzgO0vIHLW3F8OKvedz/1XtRuOwnPvxdE
1Mkpk1nj56V1WIXIS3i94/LgtC+Y67ULhjBnP1sj3TD0/qjZvQ34NS8WqHk4zoiHRFBFsc5gfFcH
YFeK5ZP1kl3cckScCx4fiYnlKIqzW/Rmbzzj2xXvOo9OD1HtLa6jrSob57d2qi0Nl7NvoAH/IUtl
nim1PpAWRDj2QPJgTpXMfkTslgzh5jn9SI4BWTF/zrFdC1lAWZ5Fxpi1wVcBg1kMKOpu6v+WfcEH
GtCerJdIuFrSGwVcBiDAx5L9koVWHPiZ6U6IAeYQu6mzhsNKVWhgXFCDJZrqIPfckl8tN+izAVne
XmCqCLRb7Sy1eRiY/bBvfEaGb01OQ1G0f2i/TPp4H4gWBZgqfwn+0fsxBL9mjNc9EneJ+fx3Ozq+
bHrooP8xy6nPmR+Sm2y3G91ezA04yTPTh04i47b294k16qi3S47FqyZgbmKwS9q5t1M3PREFt+j2
wrjN0gLFw6j415JRmFvVZmolQOQvvLcdxG0mxbr8psl3OW1uhnYDFoZtYzte3ADAcFQUqdj5V3J2
2rIhyv8Im/5C4sS50z4kjCvyHfWQJOECtQyPr8ImDGTzj9d6haN2l/bpnQUz2VhmSu3Ucwq769Vt
N+GB3LiSnrGWfTwBsLTh/kPGIM7b7ucWyAi2umCSLGTCcWXJLOgA1Pl3h68oimaHKTT/TTjSYtlA
Jj6eogmiVdDWLDxMdfJZIEZN0unxaKlz7gn3163DXfZbq221j1I78GyZHVALGc7yAoWKq8brQ9Zd
L19Y/VlAQ2ah73xaxT4muGunfzhgX3AfLZJcCQzMPBe9NjvAo27jMP6TkTwTfjBcensn3SaBN9ys
4VUY/9WYzsh+peLBLGSQ2FjLnnQZVUl8tkjhSXq9Bmv9EeWUT3+Mf59mXUNZ9MixjXuQkdTv54zH
QeAHzIcAvyGSEQVsPJcIKT1G0KRiNHbTzAEI8OV7auPTst2R8DQWf+xin5gztejph7EsU0IuEyTj
Dcy412t+9CZcvDys8OwR0JUKqgJQNVgpUyIH3pW3g1eGzobB3aULS45LLPEdNqGKa2RU5Lmn38nC
ayvCKOshTT8XVIJS+96sZuhBSiawi+iO/+48VmayTeViBb7MbeaXNT421SHl/C6vKVQVNuyEWTBM
4U6G3aQsMwqQbNfLV4ISG2Ted8ceKaBYjq2zMgly1uhBn+5yH1WInvCJbzyyxL9sjjTYe29rDohv
DHYrwHvM34VQzFxTASL8gF10sWGdupB5COJPOGWMe4eK7FQEZ4yc3siOPypYY+B+ESO4rF9YwWjR
7QZ2OOuDdwvU7kAxdDP/PlRlNuoGibg/US3hr3C+2csrNaOtaKG8U9aEJmwB4v1OROo+hdxeINPt
0fU29HjhJofkfBdfnY/T3T2QByagWm+korILJX/rzJyH6HSfY/5OJpq4jVXAAaipaFvAzr5txyrr
zuxq+4W1Kw/sZ88uEmPUBONC6kalkAeyFVxuglxgtNGvw8DGa9dSPkeweZyOzjZtyevDTNOsEmmu
KPKU7Cq3sIAUL+y7Fhl/xNZUHg6rfg3VDAxPZZg9rEVD9DQqaQTvI+JvdkaRidGJfyOfBj0X904x
ddEp4HDqxC7Maozzbd79nRb4HndHhT4mqbZnrONszH47zi4dLCrDJNGcF7gQ5BYSXeOWZIslVIQ0
Go59Q8qcpc8BZona+4oFtFdC41N0rlBem3JUE1GwGLxn1Yjb41oQbRjZ+FPlgG2Rm/G539M+62bv
ji1vWZnDdGoI7Y0l5PvKsDIx49tH//R6HwPrGoIDoHrepm4B8gtIAXCzgJSbbCofqVErWYA2WU9U
wI6aLu8SLj8uOOZteAanv01e6AoU942JrL4hCsxxw1JlidsyhaEHI7CLp30gfu4SKra1UX3/5awo
5dqK/yHF5tmFd2qtbeahl1tzIWef/GSXCqOVVeqTPzCgaZs9KRF8h2EZpXuaqlaklP+Nm+qg79rw
RiJzxiGrdfY9rDk+ii5TS2lIUWJrEV1tjr/Nkvvy6PIqPu5AkEhiNaOcRC2fLWKhAY6BQz8hROQe
1ZhLL7lc+V48PuHZQG6fvod5tg6IMqg/VJ8G3yF023ApBqCvGmCtxP1ZEr75cdkbIx80elWmr+cd
7MYvLmHcCk/w4VnWuMgSu0vZIUJNXXDW6yElV9WBjxP9UUC+bwyWO9v0Jpl7FUw7bu3LYrZm8JZu
XsaAh1jfxaeFEpbvZOXZypKql9Mo99zJHLABIz8PUcbZAT9XqmfIXqwZMbb4yZCQzkxAxMcNhmO5
F1mDdMs7AcppevSY3xsKHf+VuiaGbap5EVl+BQ7ER5hsLzt1oKBT6s9uK0fpBcRMy+oNDsX4bocF
f9xnTGFpn6dCTC9K8Je2s4kpXT47UCXFlIqn7FHY8VOQRDDtcMedoNIGOOQhK7Wm1TP5MEQ4ZIAp
nfPakrJ7FxMBhcFCGqqi7oE7c9HynWKkkH9hkh5BkZjIX+nRyz+yjFSZgdYmEZhXtTgNmLzZJn1v
u6ocJOHD82DDsdPY/Dh3SZJH9+ubmbKYSMs1EWlMt1CrPfdWDIeKC3Jpz1s14ASl1FHtzEwnOfqg
Ytm27UGZv35tlWlS6KHITFHTTEok2nFhZ3lmwRx3KZ89O+0pq8N+xkQ3YGmIo8qKvnzCYTTKj5PY
UvW0QfQt2fCOKUbUm4a001mkDDUMKlMVg2THKkbYTnj6YwMYxSdMO2aZZhvmGDRrvO4d3i9rMP/i
rhAZ6K9Sc03sDQu/qXOrcDj01OgDdepiGafcS4CUPY5B3OHg/YJguAbdctFn/UNyUzmL72+GwtLv
S62/ANOe0SlptInmtUWNFsVlmzj05TqfGNxR+y3DRnqq0CVg6yKEfR2XskYvR0/C4y2mA61rkrWl
sapPH9aQ8AugBT5DCqck/CGgZx4jqkKv+vt10gKVUMSb/WyyqiDfP3ijYj8HFNyv2+eZLID5ZsWi
daJLCLWWgDlX27t6whSOutOl2YhLJopar16fXTLvY/JLBKeIIyduDD1T9eFvenbZD/PXNUYaDP/t
EMeKiMz8zJ8Wl7vYQD3ar2Uph6dLrwXsbKTD6WRToxYqsyovBd3uhvsu1XL9z4IZt1/e8C/ATdx2
env6xW7Fe3kN0flRI476d9DRsKHF05sip+q77CwInv9OlY5TsfXSuKqWWlavJdlrME4MYZBE720m
ez20TivegI5FG4U2PWrlH6OHE55EQfL/DPGWRs86keXGPl/pjVvxUSUR8mdpf63bgmWu+9igXUXm
2pQHbZiox8pnspfXHHpix+F9l0B4++2aq9OW/WoxwbuWetBmiekZycOo+eXVUcTd4SfHIvQDmbIS
ZSeAIkz6Wb7kNceqCIoVM4+S8RDSTG+4CA01knvK/eQhYHKnM4C2RYBbaml63S3taoDqvZ1hQhrz
9njMod+7VxxKOCeF//2KVCe+gv7FQYmmQAgv0m8ept6pdrrX/TWsFFBW3vLSefTnd3Hd0qzqBhkF
YPwyHlhBs0yeXQ/ZICE+qINJtsSRV+ThULiRoDoIu09AsBv15Rfj3nfOwQLR5zsd6POn49Fihxzw
S1MMyMulWFtBdGqcMR2TB+i73/kUHlwchS9qtYDw7fDyLOy8N2bT2kfiumB/feff9WE7gTsNHVJR
dSojDhA0lKj8k/51rHelx4jx4MDH7vaNaAWQKK5l7nJerB2QbSHsyB/ncny66ePd1GHhssaI6pPk
mX9/G4TNIxYTYhdtZAmd/2X+VKNhQTfICMOBROdxjWCZ3kA7W//r1V9PDzdswfK+CVVjunMr7A3e
+WeR3AS9nVo2V2O569MLrsLGKeUL1qr6t8nZGO5bAkos2w+vS22hiuL0XLt2Ex3XKWJR9wi+Fhav
olWJjTlNaXJfj8hMP2j7IsOUjYO1Xv3u+Rtz4fjrZM9lrfH72NpkCgUPnJnzGxoMdYUfGrIG9UDR
O9j81pSA6hmPyApVCwQBe2UFyLcvfrGIbWXLohmLBixugbk+keS5Ym0yJuwGsOZNF6feowC/RcrA
HShiOyezVL7+Ujb/yoftJSfin/obWWdjRMS2HSTPjFWdqVr6W1FPv0UtZhJxkgadXBT17M/M4byG
tvEm7OAB2KRvjq+JkdlswLidsf7g481esEjjGdFf+CJ6aA82TJFDswct0H2bHMdiXaZ53xzAuNXh
ccyn3YDGmyWn//8D9P+HgjOGDr3nJEPlxeHWLPZNsiAj1eonkEqdTMwY2aRc8eS0zAGCQ/tw02AO
LNRWLAYAdmhQGfwZyj3iXBClHxIy4C3N4sQBeWk36Guc4dndWRNT7XEqed1ysfxuXCG0OMJvKZSR
7p2Q2erwxqgYnK3KX8yJa3LrQboFiHYfbJOiker/sxQzURizAhnuux0J2VfkG81316zBS6z9hkJZ
vHlOwpolKyh4oJBfr3vKINVZ2woqQEL8/SLuqb4em1dKnJLSdl58SFhl/IC5gCTrTFwVzVw/9pJq
tD58wam3uIYvnLDAYQffS3Ev6Iq07t6Jm+Zpy5/gw5uWhAqc1yOaVZE51F/0zabGLWAYK4z5ZnW/
DZYkknplFGqSu1YKj6Nx49fdXRvo/Yy9bQZH/L53wV7N691KbUcIrQXZTzK/iTxKHfkQuWR8S7D4
v5EMi9cxdBqYBtLnuInvOczt6DOWF+pSYCM/O6VeAU60TDm1PXb8cq9hLKwSumK6PUQHaytxt5Yf
yxCZgyAAm7Vd4qoY5FgT6Yc9l+n6MTAlNjVdrMDTzRmOoOrrx2VxNfm8x0nmpsBq+KlAvUCOKsmd
h4D8VtC6XPtf22vnMh4yaVyB05Mv/wJ5kTHsgR2XIxGvJzHwtlDSbwet+98xX4a/0ShtjotAw08a
a8x9Rc8EQz2J8ngvJWOldYJ5FG3Ppyz4aZdp8MNo8QTPzOKCR2pYKipgi/KCc8tMG5vX72zXKbrw
rsoryNn9ysx8hqjClS5PcnBKUSq14A2/d0NKHWPVuxUNGQT0f/q5ASO9Xo67ZpiIMGjCA4gO8qrv
fgavggtooQcipJf94vztD3oRnGFTQMpMcf/ym3CU7DBzFIESVVpQnJ5zw2jJ47FTTqMn4hP8lXKW
iPDd3/MCMEYQphRFpLsUfXSa16MdxPCY3CuOSMygWEIF1GbkTEnko4gq9AOmVKZyVVK4KefQXrIK
wftDPuDKA871udXQdeR1UoNyR0DKw83Raegg/b7nTBQi6ZaaQx2TsBrypYOedoOsicH7bNf8kVv1
fTIVJqqMgcKhSiLGnsJha6jLcx3YYDMFT7EwAYS1k3h4srlyKPxNuTnR7+sMNPZo7QOJpqdVMA9T
wLnsBw3iGJsAxqBJ1CBQCc6cDkfEaV/xU3stlzjzHyBOfM+G9bbXetNGcoiFVUljW7caNjS/8n7l
Wc2oUKBVyVKr1LRECddELnsnFIuSkrKmhtOezGZLGfDjhr/ZJ2P0vAfEa4m4OAwxB8nTDNEBaAzp
1oxoxtawS79zx/U9uD7QY4I2cdjjF8GT1w0LgTVsMfPHZDcvkUGqY+ykzVXyhNYgrRX1W0q3ikeR
cTcrg9Vk8b1fJK/LkjokjWIc5HnLCf7f56ErRwCJ4afrt6kz+ejHWlJ65WUl7382S/GMUOgicP/9
A0hAhysfundutZldSgtlpAlERycTliZ2O5IXqiz13eAs3StJ1LdOtFpp2ZBrbqBqx/qB+RQHvndh
30HEnrcUCmtnXsaVc0ssD5r8W2zOnwU5kmIImQM8yLz9JRq6MxDgS4ikcQH45aBwNKunub0iT0vO
SwbQTCzx+bTGMABKtk6y8LGTFIoF5xo6J1g2Stutohm9EyIqCKV6GkAgY1I5h5x++boIaMPxJJc2
gVmqjSC/USF+7/+MEz9IjBDcQO/os7EYzcvFPM9JqJPNeLwcRzx1GeTyNgjJjqSybTkZFRlzWFlR
B3C1FokS/4LnIEbvyLuiJxQYccmTYg5Hw8O3zkwVXNRnF7LXrtaXA3pKRI17+VHxXGuQapOO8J1u
p24sbAhUe5ahtW0muxz7bbUDuA8WD2vByAbavZEj8ruT17Bk3O2HzIOHqiPFKnxvsbi/rW6UikPp
E6TRGZfWipjbnxNOUSG4Ea36llpl83JJFWQVXa/I6aC9G2Qb8UikU5GmskSD3nC9vol8bZbsr1+u
gXuObstULN/EheyUoZGMNymKUyIIs5tbJ/Udje/+EeFXGS0o0bvt0UQXH5w4iF4wIW0ygR8s6LON
DqxQEbfM/swbycnevXZJ5c5iDPjAoznUnzRQZhk4OUUwIZTO7qgsq94ldY82JvknzKZqSFh7PxUN
LM2+IIgWQ2R6TKKCvZNbMRV6JkOLn2itQK3pm/1Ochw43zXYn14iFRAnbRWepST8T6liywj4AhYy
MKdZGZkXWbt1HXGTMor3WQR89LGI6v1ED+5KFvuEl0Tui/G48pf/wbK6aTP8ID7dE7CyXBOUeVWA
HfDl/LNGbfAMOyy/TsB3kkh17NU578VV7ewiQdvdzzYLmiif9sIPifGBFa5tGAT5AEeXoFSCYesE
9FiY+w8Ph4erkomV4IL+G3B95Af8tnnC8nzW/dxTwOFOaswvaiLQMez+wc0unbtMwg2pkbF2JEEl
fKdPkB9UWwT4HwO6Iexx/f9ZJGF3m/690/NepDnu+HHyCNm9vg7H2FBrN+/ns3j9PDP7EgsJYP/E
1cCtb7QNT5YkaIhTD9Qc3Ly1A0U/76jikpg9vt8Wp/A+5/2nrSXB+EAqTTsJ/8aQ+mrCXj/Wf4L1
lT3+A3KuWOtnJxpBTzlI8mwiTFkyLOAPDt6ju0YsZjTjSQ6gEXzEENdJfyP1y557yR6+6sWviboC
3bhYf92QXYZLQSPcciy9RiMHHFl2sR01vOBKyEsbpSSyWdcJLLdFEu5Q9qJWjTGVbpkPplDjKvkw
M3RL4pt1tsA8adsM0CRDX0/q1K0ivnwgVjfrQi83bYbp2Hb9KUqRa0TzPlIfJbjUUEDSsqqBXF1U
q+fd3yANuAQNhBN+ADi3kPTH3ETsJbFyisqhJ0DTwMf+j/tEWeMSXu6O8UuGhUNtxXGNoBKx0VqG
pTupJ5SSZSPMvC8r9U8MBLit6jybRFtlhIVPW0wO/TadHqz9G4cWfafBc/Y/5hXQQ0O3jk9QXHgl
zxJ85IBS50+g/WqbEZ0UMv8lgvW7Ul/eXOK9yWDyN3n5ye7OelYYaxhZM5McsvA6UJWAdFEYtMGX
agBNRxqF9pgV8qZ4yT/ooWQmengn9CXDdpIp4x27VsEams5+5JE/fAr5lzUPnb7M8LW1uFgGhicC
CB13doBSkgvLvgKNlksCWToDqHOan1a9v/pPSHxUM70dWw2FFU+ymmFS/bGO+IWWWygDzewVhXWj
c9eM7wSZ1az2KFviGeAndUyMbCSE3FNU+UX6yxxc6EhAEQfg0z+Aprxwg/oHICp46FY8ncbhpWGu
tUBFWf8t0IHkoEpXQG6mgcPzp6TDjZVMo0IFWSkSjvYcnN9Swi5UAUW6Wd8eUuTfp39jHvy4fIC3
G7PhodgkNnmqAQlmhcguoaCYr9nyVsdpHm8S5i96ksNReTjoj1uI/XkNQ2d89Kgs16O44tMBY1DN
x/1GIYcUDozE5+skdCWx6rhlI8eKCceq0PdDS5fFUX1lg+7SP96tq+SxfXhFUvgpKSQnl3BgP6bg
jgI9cGFJtKAN1QhY9D1mvWTI9+HLsJx/oyKOzM+K9OO82qjuB3oL3RXOCM5iXhyW4PQmLPPEb1uQ
doblZVM4cvWrwFaDA4Jsmc+z8CUCySYxilIV0XmOASdE7yqId/Y8dDwAdKGuCoTU3xazGFfA+Jux
GmdVSV78rxzQiKrWRzZyWThwUoFZfOVeVX8W2Gc5gBIovBMPVoaK9fSVIMNxXEtSnYrc28q/8xiS
6DrRtpIZSrLg0x1ZiO0xuD77ByskPTYsUFJ9UAV4/gK+FTlD6B2NBlt2muTkkVtw72hPtioilKhA
aZj1e14+hXG8G4hwkGuk023ON3NuR5a0lrg2ZJbS+QK3IjER8RuDyxw4Zc7xGcLlm7cgZS39VZVm
q8h3t6lEU1jKuf7hh+RAPaGmlThrPyy3jQvch6s/qQclzztcvEOmEOyickoK1FUBf1dP1qCsCRBf
NQFobTAg9RY7YHsQLtskcFGWVWZDm+JM6SgIFsVU1nMlwrdYt2GlsluPAWnXOUdJS63nvc8246Rr
DR/CRTKsVU3S9kRx+YvTSAR8q4Va/1LJyrPnFqe4fuLkArdNP3ZwbOEo1cImBXh2tbFLIHioTj8E
GPCaUxlweU4UwJpcZ2K6TEaMSob5IO1e7T9INgqkn1dhG39YVt5VdbQ3Sg0DP043YDqUnfkbqB42
9fpgmC0tdHxTDrCNakWUZD5xe6jN07aLDvGUpanuKFys73Pz1rnEQn4gAQBnoIWdDHDjhzg+Yy1d
co+zrnWcKWDfA698Pupfhl+FxydKEK73Z8QLFD7Dt3Mh7vqoMduVyQWrHGKyj03dNrAZttXkIEaC
TBsvczO8HCj4wX460/rEbMAvPSCdDVdjbRm/4grRdW94h7M+Bbzv6xDvr9OU4I51sUafPVmWBV6a
rVC8WfTy4uDyUhMPHz/5Us/SbeS+NCPASxtjsg2RrnvlyiRkXZ+hZq3GHv89SUSu0UBb78rCYtrm
QMlo31E0yaCQWyVx2X2/Kqp6rjzPSvBTzqmwDJbcOW3b2NgAyGoaB8fiAtwkin+X4ry7wrMiYzEl
ZccheuvnGc3hHguXMiat1lqTro1P4C2g0hcw7jQT1TmFLbWlATTKGpGKQguOtlbdRpzKhp31eNBq
OHrffc+b+z73xO1+NRtqtVk/up2qTZevDmOP43x4ytbUfTcgQpV40r70pKjgm8BboYkyhvSMsDmW
Xa00mSWUaS4TJP85054WeBBfBii835sSnAezM/LHFNc7xvOw9bKaPMGN1HHdH+ovA/MeHJoyvAFp
7EdFTN4mB/uHC/l4O40tTZEzoAXc9bjtIU6JG1aaotYvbs1Sre5VcLzB1tZe7okvTpv6/32IPLYG
9cVyxbX/D75BAgH0zBwXDIMWZ+vZ8ltQY0N4RG23qkvkw6mEnPJRV3ygUNXIuUw600Paw4znSJLe
7fay3HNntT3u+4chJ+fdgxVc3DFyOzmsFGT4NE8sEkDPn2690bDVI6xsIaarN3rgz5aySErHSnRQ
rpi/2P61TyHoKvS72oEJBwraCCwxF8y/QIf0gEsIZHKjn2nRWa1q2mXMbHL3bOhSnXch947cPXMi
RcCTwKe4TbECi57oHiPSufkQQc8u7f43B/KrosLEEE8B5VDNNpER2lvvCky0fjNNLJIE/CAjaaEl
ZWU53KxS+8x/XWdpmGU1Y5TT45EXY7jCFecuea9Ia6KDEotjp+i1F1UWj0S1B/ZMWuUijutEDz9c
K15iCNxv5qZWhIh2tNOsBGIci+T6Pg9/zkKAPEoqCr78yt23gdmZFDP2PDqjVsEiMK4EhkNOqh2+
kfhsmd4nkpeVrUkuTUH7h+tf9QmEo707qShHWEodOmyeh1RJMQgCBltlYa5sHq+yIgDpGBBrgE0c
YAPliSBgMtV4N426rVZR1IqDxZVL9xjIYj1MSWQ6S4BxqJjR6gTZjMUu1PZzONkQfXE6wddyu/rj
x8BkwOykiYln+CfwHyeDuKi3qXwQjtXQ3LrU7wolHsgLqevlRliWn/gb7QnSQWkmb//K+c+D5aoB
Gz4H8GJHu77Pg5vC0VZwkF9QwnuEfOnT0dSXKKKgqw6tMOlGkQD5h3xRo9nHUGx36EGRZkCwJ6zS
ci1ziv5SHltuQiip8tMotQT4DmVsi46gOl+EA29Dpd5D9OA2sDs0Ry/wj9axyBKpdG+aaJu3cv4G
aTS7xfSfUez4eWg9vi3EyByXGzTIoI9NX3cptMwy3kIQwr34cLw/tKJ170vKny2my9AtWxs6ssjQ
QyXQKMf5ygQjWR8pSKEErS7gMyMGmCYN/dRmmCS6lOHwjxlHaa7n0BR4jRSH/OLdzCNiwZYsnSir
+Z9oeIJjXKKU1+A74Hj2J/CLrrA4vG4LW/bSlo2bxuyU+obBSeFNdWjHGyRhfV49hfPF5zXyR5Q6
AU1y+3OIKmdG9QyU+W6SuWKp2TYjGvANhE6JiFjo9YBmllM/Vd/fy0xjYXWMDuyl3JjVjNxE/UtC
HLgGMqGXQ2YRApY82V8Bi//UjIrW9lCW4JDeLxpk+fClm3xSsistqlhSOTqJWA4pw1VbZXhVxUXH
1schYgA4s4x6pP3klF6lVrduYxUck7s74oIhfpr7oVz9e00ydBM1t/6WxeC8ID7pzAYSBLXn/FBL
8HunEbLmusZ08S2GBNXDLc1MrTc5ktgHGGsScZfZrn2m4Hh9s/JI5cyFG0g7JOmX6qAtUhzXN5L8
etzqUdKkn3q+K3X59db0SIOWyeQM2IVqFBfhICmpcOWQ7ByDSjJ/gdElCdXYYAK7wC6L6qRD+FgU
Yg3Tn9DoisFDrWLQWG2gfSHuBTmHTUAWj3b5YrEShrYPd8num14fbouVYcS4gTIdC9/tMWJ1cX51
CH84/77Sg6vEJgRXeQRANjU7zttxMr8ns2i2xJz1ZOK2xxKG8hSCkbt/SgPiuYLtXwdRks1xx1KK
baeUsniDU1gB/cAMF0lYeGQIJ1+c7xvp5asR8KQ+lOUjHsPveUCgWQFYFbkZi07CC+AziXhCmHLy
k6H0D0y8GYnQLG33QsJMSSTPP2HYYj4i2UIk2nXLfJ/fyNWuKHBav9dQ/dXW02TlYA5nIJM0ZHxh
lyRPJkiBWKOSAcncDgGKF3XWaYF5NW2VpcAT7syYGMdXQizdiwtczMePUgtE4r9JePyfaeZ1fV72
9Ef6zvejCQXJlhjH4izmzxYcXeUq+Zk1h1vmebfZCxrleeY5dHnsK4hsvA5YdJXCALQVvTqqSqlh
hnSm0EwxOoRka8MMqT8eTPGApJGYbQ6zBPC6yT8L0MD0t2JmYVjIRqFyqJKxi3yqKqAN1u4Qjfyh
Kogu+HWGgbrMN5Yej+qu3v3S3zVbinNElgYSkTvI8xwutMopv6ndyUIbQCl00tSivTs5LrcwhVWC
F0jckev9axIZwtT25afN5ZGNjyShDb4sUswzh/LrNRnTL0g95TG2lzMQX0oNcwPdqBeHzQo4arfJ
k6zKwdsR3HNmLokfH7zO8Eq+X/4nb7gVs5s+p0CmUjkbrodqnyqyFeu9wmQ3cZem5RpC/91TlRls
qy2fJudHc1ShDmr3CpxhXlmxH/4cQF8vsknKDrLU6RD0Z0zK0JjhYnnp45rQSqswN8Bn33Hwavw6
DRw3FoqCl6p3gr5JMJvPXMw7qX2/v7ollnq6gr0V0lDK+G/LDwPVYW5toJ8hSXgqC7mpfNmDo+QO
eiedha8Ipq5tlaTWNbfazmbDGaJLxAOV2eghsEup7LicuMuZrY3aTOj430Ex+g9Y5j4ALKVvijRO
nfz9Mdxti3JPbBn7/MNKWs4Lq0QsFADKhmgJF+GL1eBcfsRCQKu/ewqGodjT+OQd00k75+AteYN0
U6I69noxIol7f/KZL1MXYCfG0tsslcVr9Qh0c6Dmj6GYarEMMoIXbzpGfuIgXIOBQhi+Z64AdH24
lVBJiLtNMuczLB5XLviNhNgPwTcWPDOrrZg3IVp1Cc2XfJ6FdYLZdWVc9Fk9EzV/qvCu+mSO8c2s
AQLgH786KLL7YGioZCETiem1NvgJmaYgUAsIN8kiAZR0BRJ2fC4kVv3wWwrM2cEPlonTXWNQnKm/
k0UPZdAHiJeI1phGlm6GYOt0xafBraWnWu48d4h2ZWL2h+VhNaNE92Oe+zzI2ed9GaWnsyb/vzaX
blsNLBxCdPq4yLlqaCOT1xJHrHXO8bhOC2htu/mU0JASWfAZWUu3HKfsCtg/znx48kJzZMfrto7P
zrGmxWpus7JXYaoK06UvV+MjnSTk/BZCJgWLi4wQl5uJmRYf4vAaXMpsPQ9AqFwVl2db3PnLXilA
Mh6HqBgaHmIVaLXFOxjCfDileYsdGMVokr6dK+CyFfipk7o4DTmj7UogOglQJol54If8TxXLCqEq
ifGADuvf3QSVVEEMcjwVHCMFAtb8GTPiqpzw/lEbR7koP1/adfSPNDzQNi6mZ7FSgyOVspHxd1jn
fvO2YHDjU1wBdvhZhY/vN99QOyUF9TakyRKs7IlCHhIkxNpMBUXgcMGhS61qwu/QTUSyJBK7xhR5
FU9ry7Dn7PH/u1vcTmGAJg3f6WsMmEyffYb3ejCd9LNNu73TuGoiozMumZWz04fP0kp+DBFjZY9b
aAIqY0aNcMnWaEsvc9RrKLLrE40PGJ1rzGbZXniS0J65ofLhAYnxq1UJuNgy7A0ILmNOfM8V5CL7
CtEvzqims0FO8tpKkGG6egyJD1ojI7MlVm5Lck3W1tSbha+YSQVdJftd+aec1EKJRWB3oZLGYP6+
nPw7uefoQA0e5I88F4lm5A6hDXaYo4z//Wry6YVr7GEM6R5Bz/nANaXv3c3NSfnXKK6rriWl3Y8U
eqNJAf2kUTdm4JPBXVpcKSYp5GKdaHEgx/4ijqAQVugcCnUTTEreuWAqDUg4qI1vIEoi265oCUZV
2vEW76UQZRABNK5ytItskN478c96oZM1+YghXkWjhx2P3KgzJGMp/iXqVsNQ8aHxjex/j7syqs8k
zCDIs1T6vKrOV2BteaHeMPUFmNTf+QuDPGBSqjroqeZsIFZ7y+r53e7zoXa8C+30Jxb09afiGT95
JFUtw/u7Z9N4kR9X1Y/l8JY9zAJ5wBGcgLHKuddrFp0sDR8uxdZ6Rrd6UHk8RSxmXjfTP+vp34AN
EzhyJskiTp9YLg55O2rhENZtfddblLUT5JOYwZ07/2k4zG7dkeyb+qTOp8tgJ5L2oBQn3bvlewc/
Leal68Oki1IGZlvMBJA5k1op1H9MIiA+uA/GYja45dX4cJEcfzJbPvumZjEeK6PA+/gh5R6ndOSG
pRnMl3AMsoKcgS1kSIUXNUlqY5/5/xoSaec+XTJJBC0TLu6+dXnpTxo0nhGesVgq2Y2KJDsa/73X
jvQxtTYhzXzgUK2R2bse8f5VRciqSIXclNJrok5C+xpNd7J2GBjOJ1Mg/9r5h6tvjXkL6H2g2/XK
1wwbbHWsSS+780kJzBQEScpknWoG8DhP+EtU3S24rmOTIXEr6TM8TrkgPhX1HP+MiVNVUZ0OVIra
z2eCUhiYjHGuRhoGzPPlh8PT7pcEioAiuMhQ19SEMIV3w3SV8AfxQTggb6wY9qhunKmrRRx024xL
6d/neowKkirtiLjAPT7Eh+alqztIF3mYap+2pswE7OihA5faTeQTmNviPArSe4NTqnapw+xu+CFt
csyNO2x27KzmO1DdubchEVX8Js+4UAnAmVsYlOzydecX4akEtMCH9dH1kSMfCJueqe+7j41D4rtm
INxSsgFrnhTOyfVort71dw4bGbMY5uhLL125GjkQ/IjAubXtMuQ74+NXBQToWPoTbGx6AmsyKNjH
qe0YQiofmpvfO1PjklCLwIaAHK/MFLotaHL9aQHXzTOIphcp6mgl6uzzRXs1DZk3nbjRb59WkQ9c
Q00FY55ENWRhu3PDR5JzOAmfmHeQKPJiOxKiMw2PfH1YnzclBbj+WapW+7oLNiklc3WDv49jVdBg
BS9ubTfATINHjA17q0UFe9x+kcTSzIGcFohd88/6nSjOfZUx9raYNOHTbOJEeFXSpB0ki3L7hB68
48LmrzL3hMGWromBonC/WycRsUN9v8dLxCMVcwdwzFN+iubn5zr9WyK1zSMONLiCZts060tp0ZR+
Ow53mPkmULDbAoPalOib59q/UocEhkkAdMg3TLePQHmAG9O8HRLG3FflC7V0q8HJcvAJQXuy6eW8
7dN+WnCzz2LDerL5iEZIOutC0kzLJyhD3zwhvJz0VDHTDFEEcyBodYF9o2Emwi5OG26+WDNlYkfp
Vl5cpQ1J7TJKSGx0Thjd5bwNFJhU4S1IqE/cC962+zU6xSIz16t2b7C9wuphRC0L5X/VeKKxiF0V
z5MHeedMc79rAIF1IU4dQvPKtKd9JWQS/MMsFV3ixPdMRCb4Bm8DvPht6ciNhcdh6fw5ozwX2RcS
qGBonozwmV05vWx4Il8ECzHalFEETFNx/jnR+YG5d5epNmjH2pi7YwrU38PwPTuDj4JTomjbNpnC
CvcbI0kK6p9EfFTUHnX9fF/dRhJxGhgn+2nzw8VAEDlWmTlTM3XymjnPEVEkuNJh2ynlzoVJlcn6
BNcOcdvmzzl/V01hcr5smzg+39wjo7oD9/Fo/rImcDhYsYtNN/zyLjo5DvovTYIWDy7ZqWKew7cH
Xa4up8+9Y7nuDaDRTcfFh6z7MCM/kkZlrQ+dq1u7HK3LrVWZBEn77K0BMqE28ihh79HYTqaePiiQ
C1XD9557hH1SuOFt562KkfU25F3tgZYua2WB/SQx3dg3BGPKHGQvDWrbw9wyWyVGWb/w4MMSjkIr
LEMBOLWV+Dc+Y37PQJYidWHxSDcrQTAnQaqVgTwoXaRvjReOxs9Vh4HrSzqCZo97TvNWHbIlZZ3N
xekvVW7yjJ8ua4UM3qJAlMIeSpIekZbRmqd3riKEPQfcOnMh3S7u3kavMhZ6SoZH0fhrxZVYOyTu
KvwLYENR2qmi2hzoBPGjYnzsFOItCL7h5szUh9Jg4vgVRDXxO+gWQ79SzTWQll6VCj4hgl3mnSx7
bfEV/1HJ5J7Ci18G+t5+PQK+CFLvjOPs99YYWaoSbwN3U53x6a5JwFyCTt4vrwSL+yqUnG3WHs44
4NXg/cGrlvfIFTSzdwQJ7JlfY2aLml3IEMdRyt59S/pw3kopwam0/474Sw9VrPKqtgHiuHEm1QQi
Q7F2fNhyMiRLt8obv4ne6Y/3w2CTooJI5MydhZVvygA/E4POeXOVEVxGfIRYcsFevJOu9/tqRN0E
yLDfsMj1a31pvHWxIlF0Gd88FeL1MayuTvoNH2Hp0cxEnJ/7APVQJa9ShG0VRlh6J1VYfD/wvvhs
kTvVv/0kgjv7cdK+dfoZbLF/GAGOBAbLVfrAlN/DKvHgVuTvIbORvgOpCsNQGsXQ9ltPcYUXGW1f
asveVZyJRM8UXZw/Sl6tm51SE65YlVGFxsjaTtYaaQXmIBUAOJni8XZjYXdsZFYTeFWPFniBY6HR
mfxVPvUe6tSlLkzQBV6/4D9Z/Cy8HU4yF+7ZQnix4MWIhRedKkI79bxAbzl83qNlhP72AJ40uzHo
fOgJpzZ+0Qoaxt3kt7Juldt5F8sC1AtAaiGPz7IvvYf4NWDIEqfrOHvnb511XSjX6tBSBJFiTDj2
mKhcF5hXvYEyhTC/J5NYzo3pRtJe2tIK66BCJwP2TNVFK4GL2ZEoR019dsOq+j7t4LpjFrPaJ8yf
7zgGnXWERxQ2vbily4tWi1lecFUP97Ang+ITBj8qhdeVekSNuMAQgh5mAcJjW7cRLpPhK1SaCuwh
5pBM8MBpdlbUbQDlKrrWR1/c3/BZ7DLCKvTuWDxMUmrhpK4jkIO6zpYUIdW66i958dCm9d4nfp7a
gutsS5KHaOrpikPXUNpPb0gjjmrSivwjx4tGLejjW+iQpcJNA3uPmNpeLQlHw5y6QxXiLpFD83As
IEhqjHT15ZEohXXOvrvbF4wqeCNzQUJQRlrxakwSxiVL8lWiJGt5ReODXfxxPF9xh6t9zhIMHorb
hoQ05Yt+kuvcnvf/YG27wRFZZ1E7xxMXmWZgfBLWX0mLCQzivRQ+KGpnoIhGHFd3Tj76ZeHJrB79
IMAmm84fv4ymVYbptDt3JlTfiqGnVAmZrS2ksoEW10web3hRbtei+urUjPwlyIW7+l72hmYlxniC
vWTjiDey1jpOL7EUcECu1rzmO6EIEcuLKOs1HyUrrDL7BknsBLgD8rum4gqG3PYbTduPU0SSWv9h
ZsRo/lpu/usLDJ0d2gRmuPyznIU1i0WJaYsdhQAa3B1zQhPkr0yPaRR8eWiKISwuOrhPWQFf2s5j
E4WdsNQa5soGO53WlkmKwjSc9ZMAwO1dfibqpgacF4NhIPDeLOG6b1qlmLH2gU4s98LtsyyINREx
iAY37wUUwlxUBdAclch2rwMjYlIVw+hMX3DwKmqXNv+F/JhdrUBa3CBbhgK61XOfLK2W+kRbIMOM
idYhS62tWwOrzmrmc6AdNmEIS/iMWZHn/yZ1rBffGkC0BdlvIOKAS2w1TxEe0HiEolwC0jsCQQLK
/5HLpg86falqOqbIcDzQ51ctxQI1JLmRTxFUlviwJUNthipi56rWYMVNCnbK44gMUVjaLc7h0bOg
c9pKTPLCDdwgD8lDf3ChaCK0VMgiT7QOISAEOylwdC7Sv58eSTJWO+2s2tIHab3NmyVyo7pZGVKQ
sDm2b0VwMwLhvNnNimERYnnjXgvv585EwHboWpAxJ6wd1df0OqcAbvzhQhvM6wlUJeoZjxJp5m3v
aocbEf9gCZu4g6W7vvsfkhzq0rPa8O5BLt2f5SkhnWi5asE03/Z8z6MR55khPG4VoVA7TQG8TNE3
B24FNQ2CtamnJASWJHxNGotAKZCkLRquW7ajHrh0sDFG2gVe1+U+gHCAgBZJS8WALesViK/n0yK3
NM0SB8xmcDRNCYx9T3WhVUU37iq91M3P/VMA4YH+BTjeDKUIovGv4o2hPODjaHuyOfJ5QovOoZjx
cvnQr0zkcqAape8VK1UaXhIBEprA9fmzaK+c0W+bzM2H6UAZ/WsbS+QK7qNfkmkNjC3QZvUt9+b+
owhCGq0BG5pqajxVMyYgBz/lE5diIKLYls1TJDSedbmCGNtXPQdu+5IjfZG4aiiAL/VmIQum8hV+
2ETNapQxRHd61f1t7Ku0X7NJtO1cl3M9vx3Oq2Quqt4EZVeoudjopOV/c2wd2JNreoK4qBvr8J6D
UzHz0tBsbGJN180oyK/2iRJIjPBIsn8J3JQP6gFdkH4hdlffsziC6kYrSTFWHBK9Uzeq94ZoD4He
5HZOHrze/n+iaBI7tTUHdl3j7I6CXK59E+o9lb8dyqqLyJDiAJVtLKvKkRU2srfY08lVXoxT+/q3
BDTXEWrUK/gcbY2hz7Vbkn9qXAu0AckOp4IvGUSBy0kDM6gMrCvY5qVKVScZfLNNkom2Jueo7V8r
QW1qfBK/Ye+YyeZZ5ZMltpYpY9/U9k/ojrL1Ipz1fRaMEWNdNMNxLbBB2QsxTcZIbSqpF0RqAHQE
M+zKjOoGCgk0zzdKsIrj0wf9OK5Ejn6UvBxosGe7xz4Thn/i7q8PykAPQH0NRmgg19hjQOCLx637
BtZForm2WBR2+j+P+Uw8mm+l6CkvImMr+KP7h1YQF9gymx1o4IJgVqdmmVMdJ4XGqMIac2I/8Uc6
8Yld7I0lBmuyW7fYDwzEUHHE1xIBIJ2wh0wV12Qm38zn+FuEk3955cv6Ciu9HX7m+z22mEw5bo5I
YqEkM5lh4+PeH66FaEZLp93YlsY9b3ISjrqwxWsNXKYFbHlCFbF/0KP9IJiBrJgHUHmC2S8juza3
T5UPodHolxjkcRVDCP28qlq/VkF8uAWezhpLCOAUIRhQGb+9nlduR+pAx7vZhzt2NaO3QSiLthE3
2q/tC1LR/dvXW8g0an5giNIYw5+kiX5Ij4fi0AWDTSGgpTB6sQIo/M/3CYMsWyRKc5HT/8dH1Ste
kUF0ZT7r2a1siZxZCAiFw5qDBdtOon3ZK2ntPy/BsHe9zVq2hEnr6wIRdq/geedyRmk8I3DbKtuv
wch51fRB+KNMXyoHAgO+LvxM6MTzWY6bkajFr9GntkbQzrO2gPwCjB2QXZsQ4yZG8M5ovAp+TMzG
C7s3291g01AuYXBUL3pYAwxtrxiufs4ifeiGmXHoKG4FVH/8t8lBaVch2jjmH25uTTZwjgzB9KEp
v0g1FPMK+IwqOIXn5slAl0qC982YFaR9/HMNDRtg6+/p6OB/gDA8KNqgB228P+peeTCxq4vmtCtk
IVbmsv1n4XGAl7M40RADQ1noAdaItfll/V5OK+6jQDx4MBNxESCloEqU3FXGs9PgU+eg9XbbAxbe
cUwc8EzJw/Hy+O+9/6Z9I1aTVI/nKqMbchyX579v2o+gGR8fUKZNCToLTG0PsgbgGMbw9zQKHEem
zk6L2tgxkXzMh8pPwZZ7jymjR4ubYGKqRTdcGRDRWJTyNG1Jj+UlNvrWoSh2HaSfxnI6S0KSgI7o
nK02g7fKOb75ySf5nqbKMAmz4XOgZhBJssCBdMVHpJZG+PU+R1/kHJ0CEBCFP+zJxSk4DKSH9B1w
RJXYiDgjpD3vnvFm1ZXHX6a1ET94V4cq9XqHSHottzkAX3cm2fD9LSyJJy/YSipf4fI9ONRBTZU7
or4FZNasI2s0ULoErCiZ7YOwqUV8uqt1wHCTLrr2/VSTdCNXKhIDirvM+OKqHAmW28rmyHPM/w4z
pEmigJ58t13bMZ7T+XaFONzXLUAEJlNQt496+lz0PAeNYIq8ONJTa+m6/UoG0uxiKQBsb4WDiqn/
acv23+6K3aRPsStUddzF6QxkF9G/GZD9YCi40qnTVMSMPcjVZhEZZkPPHaC7ksNlmbHARzxnhqLz
LUiFinwbcj1aGLeTfqeob/pz/KNOxljLFLqGlviwhJmYp4n2Zsr55vcWb5ihVSfrcaQlPJAZuk0U
l9/VzcWa2P8tPDtQW6VT/XDNFavvVzWsD6QiXnTNRu3YR9a1olvas6NfLC8LcoI3GIHPAr4JR3p2
fUxKSD0fABncQ+YplpWBs49zFARaSZZT5jp52Iuabo7Z04HTUnWizqX+Dke2S5tirmLThTkQK5dC
ImTvZ8vgPEPrGAZ2nYmIF5t8eTIkyiplH2oKcmJbJMTYNS2dp5yua4QdjLC/O1Lz9U5aovATbD7O
jQES+AgBrDTvZQffukNWi72LZKrbaPdnb15ED2pe/OeUrSn3kw9DB+lxpvP0RMpDUJL55zq/ueJc
t/JtxxSEjBFhqk9dbYq9uIdHdEnWmA67xh06zmt3uYooejVLXghlGEMc2iF7P1+nXaoycuMaKyA9
/bTMcSK8I39FapBB7a1Jql+ySgCQjqwv+0mi3Qeh+rRRNR6DtKT5RtsGpYJKV39fX7shvllWe2Hg
ZbYcihupKVa6DoRUQotxhBgbdZgK9zCy5nRTAVnmZjpDmuYrLt/nmFi53++l9iVRkjU1EhhgMbHd
fGNcQUKO4fIQt8FeeWUXLhrqp0+tjBdJqcmC2ETNINtG+ZaWkc97S1xHb+0HdG8pvfUbh8zgxvL9
AJURtnIxwwqLrIMEtgpk9QA7hAt5WoR7wYPh0NyoOAfOBwmiKy2KetKsOjLR4Er7E3FdQwRXoquT
YJh06ZgAIgla/g0ygf2KGwHfn16Pos+mFCmabRhhKd2VhkPTktLNHRmjcZ3ZJpUdu3has9OBW/z5
3tLuFBx5sRJi76FO6eSciepWKWGxoC69QkSJzgjvbZiKKtoZeE/XE59Q7wX6dvbIOjIGPqoosPLc
uOuEgWpaLNjq6y6Q18PyYdyiBrF3k17TV2pWQW0pJvIzEL+RZvXfgKBPT+MBJW9jK5xWsChPHjmm
qYCMkOfjefTfnnKJd/FmkaZxQ0NPqoMvZzivSCD/WBDyWqHFPCmOH4JVR1FzKTM5tWuSj+a1Dkwq
oMIOlk1gRy0t86RCz9jSPvX+cqW/OyD1qk/lOWHYszgfOT/Jqb7quTL3ab+78z0Vm0BohgT0DYab
s1gaWD+JTPi5z3NpTOMbqUhh8VosvPcaRnjZoABT3elgfTSbGLLDrccIhm7BHZUOSZ3DI6JtRB7v
6PUuBg7aIcAnOGlxoVAbH154679IiT3b4nxMo5QjpndJG0lM9dtMW0kR3BH3W0oM61ifsun+64+T
uV/z45dY8uSda6cRrfYWutSQZQOGj3b1O6DqHG//H3dxulCPmcdGjrp+GlrTmv/eewx105qvQrFu
KT3u4MNY9RwbYhYoiEv+yFzC66e7eot5ZlJibirm57cZzWrJhF99bES3r1xrOEWiZwuFZ1VxNYtT
SRfxAWNzt7GhxA4aM/tVnz+2bmyD8Pe/BCUktudTzKDs1jT9xO7r/Ur8JKEJ6cz5OEnJrKsF8uF/
vTt4iLv2vdjDUBLIFs+8xsR8dB6Ycux5w83OgZgRvkHC4Dln0x9WOOrl+Lm0rh1nvMdsiZ2R+v28
BMGQAF14aI16BZ7ymXFz9HomFT0Dy7ixG0SIENsKQU8JldOAv1dR3COwRtuV1x2sJZIxhOkSsQk4
SzW/xroBfYol5WWA9j0WFz1hCSK7uH3CB6p/nTfSVGETI7PCbg+uf2AYIwbAvXTjp6A75WMZ4aPM
asYclf5IcD00agFEdeeZlTbbIQJgLQmpFgcKpNXQO0igVXLd8gUYeMGDV6gEluh+kr9XBnHtnVyq
4TabQZHvjybWmuTcfNrhm/7HJynxI543t7UjBqjOT87G45bxmfKgW6j0x3SJ+PTktfDidMiHSOvx
L540hngzQown624ckGI/EDGkMIJ3B+ERLI1URvNHUvxqWJ/ipXkyYt3qh1ZnpzZu7IKMWGIiNFQf
euYFBBkewQ7VB+dSndeGAzx7ahPVJqCkS7QpfXbRFKuIWOvv/QHhP0XVg9L5PZzAA/r7+x88qaaL
1KvUULxHkGN+Ml9MH5CnJGeIzEmUVJUwT1cX7IgNCva+Oxdyw1tBt6A5YHcQnQmizhnojkCPPreg
PE2IvQrg+G02koJL6J5h1FcH74xHx5VeNY0upRhMdmXRXBRhGdHBqZ6/sMsTOjQ6kLzPG2yXCQfh
+/8ZXq94EucXUmGdsGYcueLaSuu3Jq86wnQQWxo5ro/CVEyNZnXokquTOnAeSBejAwkPa+HZE9PM
XAvN6z0WoFs65IKnbwfvWpLISnyF6NsWSnieHPWGuXHDKrVbqjSEjaDJj5J6Z65Uc5tj5BcFqjR2
mhf74G+MrJE0hZqRETdj+LSVp1bll0LiqbjNSgY8bMTLsjHcniVbU1P499tyHvdlPcwdeAkoCxHT
lExrJfosWy2eIas5/uRijM266LZi+a6Fl8Il4u+7Kij+YrsYdX9UXBrlTP4CRc5DevK/2O6pu035
T0YNFR4yDOoNnHwV3Tx49cGwg+v16RwS8/G5gYodCBb1PyRG0smY5dzCuYyR3l9gDPm3gAL6fbaR
PcuURtYld5DGlX62QoFrnd7YqyZCLMOXQ+t+iq8EflLMa+/Xao6A2vQ6MMsjV8WeH00F9lFrn/RA
dZoos9Vr42i9f1RLyyWRPlW2Ok1KmQNz4JgHHBD1cLxLQDS5FcyPoWlGaTtwH3TAIZQQqTVrkuH5
6sGP7kzkoFBUKCUoectulUTBwTs+vUtkGOYSjs4uK2N+fzZN26ydXLmRk2NnYGCpOPsxZdcpo6Xk
/+EB7/1jfV/tUB6OaDEPsz7lrJZDwHsRaCmMl21FGIaM9cVqJ0/HJhMYgJ6HE/trmqo92ptdWQHx
ryN5GZapKn3Y9vLT47rD8WW2z2egozuje25U30Ni1Vb1Hkl78GyCEnSGo1aZEXyvg+PtVNl034jp
pxlemKJ60fxxZsURpJ6DQ91SMznhpFIXW71qSY0knaq7NHww+rULQL43Jf73w2xCuIyodHT73AId
pXoB16xB2G9YdljqF06du1teeif02drOLRjYyWKn9hsbneA7yRqKYZCR8EYxN9l6B1SPEJvR412j
O7e8UOXDNdcdWSr6kkxTyr9ELu4DPO7cA/lZEaBhhskAAwuoWiZYoEbl5PqF83wC2NqSPGlpHF27
R7YYu5rXEQAy7apv0OLNalCxuQOqDhv3aYSo6kMrzGLg7ipRTtojObGVM6IHXIH543ZHLBrDq7yD
oJZ+AMhKv06lOxGmsB1tJCaZNvH8tVvUZ0L+ubTvdnAseLoVvqwqX0Ak1FcVBVtD73HakNNmx4MG
uxHnkQEo7FjPNdDsbhHpwG9Q4eZvk7RXZbOIIEPhFS6f17qiAxUHg7jqFBJ5R/FfVf7GXF/49bue
pwEMP4CO6klg7DGjxuHTHmfuXXlpLuEUDVpx7lYZmu2AJaz/VzG0YFWj71tr5XbzhCtaqExcmf8N
dH2klV8RujDakg0Oma8GXYjO43MYH1M6rgKyzRVp4iTGiEx/c/ndl52FEaCKqG818C0Y9udszAVp
d7fUs9uMoYf/lGPRu9uXXDGtQRfk3sJkTIOsSM30aiB7n+aNnkd6tF2YNIonFxYQAYbZgVYdcqwf
ZZ9aquQSbIijjeV15IefUH8wwnfKi1LTVngpmH7f3/MzKJbNLiG/Tl5nY3kliHHSQS/UpxdytHw/
O37IxjpKIui5HXx8PvDC0/En7zITsTS2TAj+A2Sz91MsjpxCESSKI6R2ZOJVnYwOy35yeElAXBTr
eP0ATioFtwssHChE9SJkfEVgcKCI+JnAFdBxWHGc10lkvbrLvwOodshOcc0RiSSz1oeOe2IlWl0h
rMvT7Kmlhn4kr51T5TwqGIrUYAfmbpF8wwWxWa9t7loSJiovWNwd9D/dlC4Y828TdQWm7ctRjwkQ
7xjjqMj0P4qaZwJUwecnXVl/Krx94qovFstsbcBu0/64vo2Gm/CgQml9SXUEL3xTXmXfklWzjYiu
oHpDNcBqMX2goQJTLZWv7/oLFT07saPHtjrwWJSzNdAjVrq9gkN46KBLbMV5ER6KFJ8lOLZfmUeQ
OUyBN4Dy8YFK1ElI2F4/47bVVVPGL/PYl2uOH9Qdss8SKzj1IMGM+Lf6wmuhdrGbGRLbvqVHWM70
dZ2JymgsTUOVGHJ5BsDx0TI+dIqFDuYnTML+WZmpw++MfWT7gtlZBvkzTX1w9I8dIeSxN5pfMycV
K0LJAhxWyPJPw6h20IiEh8zgIIJG8+198ZPHzvQ748Pi8OuuMiZ9O1AQeLNFlrC+JyTbTlNh0e/Q
W+xhrx8EOrd/9RXkNtU7GxT50cIeIMNWEvvAdoNiTnOipqWXnqVpnqmt96C4lFHzTsoNaS51zYLX
MV1FVIWCGdERESZwd3dcbW3Nl6/hXOQxHt8zkeA0V11TTKupXXnJRg4+fO9gU46k2prgKXf6S6GA
Fc+bf9QYaNQWhdq0yWi6YGBc11ueWZckeVLmMf672pfD1AIyD4GdyfevEunQSvdWUBQJsoG3tuSw
mO9EYl0U5GSJkIgH6jHcoaV8Tl7DqvgDhL8iqG1k9gHEp/oJGuKrahraMJAKttVAQpYV0QLjxLaE
zzYF1687uF/ZNZ/VvEdjsVfKihIaxdAi1XZo8blLXIEXL6iqs3MGH2TG62vyRtn2Hz0SyzxDoosv
9LxM+ftc4SJQvAFtDl7SxieKpFg9bFvyd/m0nVZwSZp6wk740ZTNmMix1GgDaqesVhIRFcg8WKcM
56BKjnBwtNBk1xjUdvDi5SaNM0UHLyLy5As12KMEfEbAIlsCKt99iTzXnMM2UY4j+Cz3TpvBDQaH
qtb08ou2P7aaUFNGIiT3FsQ113hsAxLMhd5L4Y4OdA9l/vtGd1C9dg2Ez7MpXVIOUMh5e8+zUSw9
Y0ZAk3AfAXbrTe/6sX8z524i+zdJdJWTKwZIMNA1zpBV/nN8EAktd17M7Zd7p95bIo+bsLJp94WI
GGVsloAOKJkEK4m6RFXN+oqSpKrDIBPnpcB3Du24pOCN6TKWs1kk/n+e+3avXUQHchfU9B642mqQ
vakELDnbMZBW5TL9gm9/mjUwAyc8ciWg2axAyYVIjY+AF0TuoZ9ExO3EEq9AYK91A3lMLTDRTk2p
lLFQFM097QFpGJRrNxQer8TPr1eJzLe3mLbt/PTpFlXZWQ+GoqnEs/t1BDsq5QQayBrKGBPCueFe
r/u/MLoPjJjF5vgKjJbH9wxP5u/79zxICbnr70pGL3P0rJzroDpF+VG0KwEQ3+izZ+Sj8xZ/NMAj
9SceCD9waZe55izsP6SC46eoycrRqbJfGBXMOwouQsdeCrgRqErsPNgO/eVBwzd+O9Zi7kLyIBLG
aMiB8fOymG0uBRT6FG+HdQwQCm6N9Dm2dGrAv3oU5rYwRdjApdKIpW96pHtJArrtBlJnXyxZUytL
NnCqMhRqu6vkDCGevO5A/h/Vr/JxjBdXRE2yRNS5v9iHx2RbSh434cHdHi4bYlEJ0nCHRWWuMn36
TvQLjTT6SQoOvrlhj00YjvCA8Dp6KDoKgMIJkrw7avOSJb/+LywIhugUoKXSm56O6kpGBDZ3a6lY
Fc4IEGUE3rkqez5+Gr5fFGr49/dtH+gqmzkUWh3a/GEA40vj3CryJMRHOjLGy7ERAdt9BuDsm6cn
kayvIuHUKW5jj3iNvscnhDfypeQMkqEwbExVb+VdqyVk8l0+MhjJbT4lU1ELEp5Pr9+Rqq3tX4TK
k/hyS0clnj8mY7kuAaU59iR2O6W/adjoQWXLmhR5sCK9Pky8kahRbgwt66LciQo3s4GGaOfKJR+p
g1KLIXIDGY6HO8adJI6jrvPCIZaRkPoVD9AsNrtQP73Y8E/5FW7Qr9NzGLbePSk4iNuiSsnFkUmQ
Ynf5Xh1P3AHdkjZJKSBajzyDYPUEXgpN1k/NMKnXkfdcZBiVxeTOvZ1HQZW1VTNv2bqUQZGNsFxf
MNn627WrZ42ET3oquncyyueUdZJ1x17jXFuClhdz3QCnld9CAud8l2VjLatHsjOgzqh1Mb3lAxK3
IySH185gr+xMt27b+MYRxrQkt2AT7ZIYhGoE63+QAmA32kI5CqGumB3LgHVPyxQRKLIfLzdFloL3
MrYHzt68Y5Zx237lOHrTLYuhhNdkfFUASoO3eWz2Fr7Mux2EUB5LPotdcV1yFGYrCQLNQOMAoQ90
AHihbIxPyhy02GxaDP+5UNkhp+9nFNc8Zpvkc1I+rthlA7AZV+albI5qOucFguzvjUctaa83jBlq
KIAH9gqXHO1YfC2H/Fr/jnNBitbtczs6r+nlZ483aPiOcz7eEuLTfE+K+S7MipdfxhmJVgjN6gBr
nijvUTyx7pBStVdj6C1Hh+oDJrwMVfNEH91XTYpsnii7pDzjg/xgAtrTnfQNcG+iE6PrmPtPMyjg
619ZwBPfAxuSkZ6MvWsi9MeHamFrqS/GQhfMLREOJHX6srgjQaImA4+2cN3uB066RRnagAS/3h4I
epi1iZ1B7ifNTe9whONtB24w/yFsGVeuQZakBlBVXn4Qg028QV6Fp53jdNh1oLOGshPtFw4KVn0F
0YDUMj0ruwVNlsOiNlb2BqFUWYfHdM/XVX+/rVgdLzW2qu1a8/xUKtUDJk0q5mKXsnICoP8F0eeP
SHcJTfD7Lkk+J5I1q7B93pfnnAVQhjdVt1ANkTw9ELRirnXxH5DzcSKUvKu31yBNnmMcY9q1zT1r
QrtZ4FI2lWKt02+UcIbUSG0sifd9T59IOPlrzyYWVLymCucarGZt7QEctMST6ChuMCQi+URODmE2
UUk8aLcCTBVex5YHiEVlOMjTkJRRwALBe64/R8PTsVgiULpAPsBWOntqvxqIHYuyAqBmLfIqe2qT
ancp4ro4ERbfi41ElBxnXU5A6v2rFTJyjYEVeQ9CC18ETe/X8oxxkhHEzKbKeyli1sd7b1mF3uOf
GZSLWHDnW7c0vhzNIh017u97/A8voer0nraaWCDjOtmudw6etZFxJF1HcrAIYZ2fvUOCURQEbQM1
QrvOhqTdfwKZRkcE1EekFdFVrrfW0P5xNP85PS/yLejAcOIiMlDu0V6INe7aB0v88X8ct1/J+GBH
uuLplbtgW2g1Dv+bJlrS1bunVrTRoOyyJEzCVmk5qGuFeQLHThpVRGo4LZ7Yt1y7neZC5tc2ws1W
yFTKjHHRXbCXRdJwAQMDBSN+zNoTacZz0GHAVxnaXoEYpWUpHgfCsS30jyZAnnACvS/6f3BMCErL
ZLMGsxZIPhhfXo3uB5xJDtCCud8qdwmEn/Esi8cTibIe+/i+GoUTGKFLlDZaUE8nMblJ+7U1lLtf
MZ48CKmgPGaZ21iKIVtRFKOz4r3v/88s2JTBZavEpefIzt5nlhv6NZbUVxOw88lxEqPvPA3ot15j
GkOITbozrVv1PVUX2sHbn2AHaNH9Yt7tMZCRJZwF+ANVfmxGcPMpcOKwft3nYXxNAmZXhNJRrMCi
L4VUzzuuIQAG7fIxpZ6wNftrsDrAnDdsey5sG/n4XNRxz2boi1nxsXV9SnydifP5J6yCOe1Rog1P
VtLfkEGGAEPX6XQzRf9pi3vcG48S3nwukx9NAL59tzyUU8aQcVMUBAgMQz7crufBLA5UP5FZwOIS
QL9SeSlnjcPdJmfkEii/cHyrRoQR4HW0gzuGNglbox+NuWSsInZD/Gh8rl5NbDWjUicY6/lSHlXM
RKkB0ip3LkY3GnpOYyWcXYOmyhWVviydCqWAP2Kaywi/3GSYbCaPQk+TFAGVvDvr5v8WVZklJb4M
SCJeFsRe7Y96ErSR83wno3xlq0XxFKWru5P8XkV5n5jvaCVGsZtDUFcUAdq0SxvtpjrbT2CCEn7B
8uJk9dJegUmOHv61OlCjDchH9LZ2xvNOAUi1tzcj+AsI0BlswMgUTxxtezoYQTuhEf3tLgECbS9b
sOxLCHnq1ccyuN7xmlEj7TXTvBCodXGmpJx2/F0BDUaPy5QPjfIyHTD3y0FpBGeQyBzrzE37n5Yn
ivA38oa63wb3zudR3Z414aZj1k7/LNzVuyIJbqlEzWGdADhpb4EIMZjKcNuZoZOOairr/48YHXYj
wJfuTROnYvnkQX/WvKfjU1gtJZquKbegQsE/gYfVBX5wIrXMU8gcmcKZt+5rxR/bVH7Yo+hYWxQM
KE+pWr3c9EW2WUVWennApzx9Df4w8wDbFspyJA2bLyd4r3zicoaoWc4sp65E4X54wG+gZ7Tak4M7
L9tUV4cYmUa3kgnW+RUx54xZCu/OWR9JL0FtJbgnd0fvGtfSMkwj4l/w/Ues+mDx3i8OEYiXYWeP
A2YVz2GCU2VMkpUnzR3KiMWkJzxNa1F7eJHF8+TVWf2UBpaJxHqPcHdfsQ1wFWeWNZuuSAK+GP+M
mPXsM7LDhgzcJbFOUKjMnU5wR52emiuHbQtc+msgwq6FbX4P1MWB7LD3eY/0sIcfcIwL0oWAo2sn
U7ozulGtXZx4d0bwiL55k5duW+aMrKxv2pDNNKptIJwjSqvNlJblhK+13BWAyvtnWTiuTI4Krn56
ULwR2vO06yHKDjI7xhOtxCP00sCPEk37Auyqg3Cythn4XUG+1lTFw3tNerC9+k95ZSpQEqKpvsWL
iT4gV3Ja3cMpL5/C2F6k53Xa62OMijpBf59y+TJ53T7XTQ2DdI9DKnQpC/KBaNidiq0WQOE4Z7c5
2ny+B30aPZS3JPwNqw/mv/uJRX7KzZkCndDFnyDEx+PcQ1ZHm1pH28eJn7Zzsf7x1mo5G6Q0eNEi
r/vXu/i+5SFmDuMszRicqSnEMBRD22q+tlwpSzGbJWan2K5jOixl2ofqafK3HlHAuLGebBm/hUVH
jFrv7HwbMdTRzusdFnXz4erapzQXPPotxuPKm9vX1M2FHWrSGWZD5TyFYHgtEVZOvhopSz/A+0zD
jJzUYrCGhqghaCcH8O9YhTcVleLSih/W5EJepI8qap/gT4BBKGlriHNTMepY0tnQoOhiOMMKz4hR
9M6Yy0HjzKh3YHemdVeZtgzJC8S7ezxUnFVQ2Ynj+HPImo9IoxctytopbNs0qmK99bUhzT1rkBlr
0jmmWTA26j0RCJht6FPSHtPeBAq7WaNzP/eopGb9cjvRsCseBfYGNH0CqhBBjMANFLtIraSngOcd
oZ4XPwlbx4kKJfukgm+8PYNXlY0HnlYwQADKPhUue9KkgWjdd1AHOpRTkIY/GlfRxaWOSI0uJv6i
Cwz9BLaYen+nju98QoqLHM2yhO33ZQyQwFjMyju0CUCE1wcLKxwXlE3L6yBNsGPqkH73rMi6nqih
T4aTUjF0Fq9ar/WZ2rRvoCuLir6+sfBer8Mi7VCjDRAUaJHFE5Em8xppwOmFbsHciInPu5IPKgkp
FX8Kb5DIO5MfhN4oLibBv8Zqs+OrSzfxHfwp63Xe5XCTJgqIxtNHYlN6kYGGwy8wuU/9QPLaVC8U
lrnA5OZ5WqWyCnHIG3rzC5KMpA/4XItiobUz8yQrrxA2B/RYgXKHmr+XXwO0u1aUZquo8QQBXAZ1
3v78ystO0V2b+qQv+libklxTlRtDsZUIcVkaIaFYyGptcQbpHV2Y99mPFoYYz8F0+GEeoeYQEC6v
JJgB4eUFjZGeVciNybKmgOtI10Q3YfA5nLdaolfyj2HeFqnt1UliRN+ewreCeLIbAjEqzGIkwe2u
B7P9ZAEXUEhWFKdMjESzET4ewgJqt8tIVw01vn6rV1Pgk+EF9z6iLNNlCXmgf/mMvxjzoaEHX28b
KIzNu5LM4kK7GfsYaMeOeRmYc1Zy2Q7Bz/WAjQd4ajewW4jB6yEnBWBL1qzPeDQBZ230otg6ZC2r
CZ/Wpulwmd7BZ2TejZYRdvXw50jYOnG6wiqA5C64QyE6yAZgsrB50xgANbpCcbd2OSQ4gU5CVYV1
Zw/PDSQ60+bYShfZ8t+ok2h3GT6qtjZH5jwDtOknk6QoAPrLBKQF+KqfmRu38TCkWds0nUNzQVx/
r9kiXxKdUzr2ZEgD3X1f83kRRCIf1/zttP0Ps8BNj28+sLhbauwnxFT1o0tTq0kbOCxcOpCfKrGP
ilL5Ch0S3GXyhywSf6d44e2gnkYZ9nbn2VxQMUZDIKBw1Ylz7A2ioTEVC6wK0ji3RtKi+TudjjwM
L2HwaCVUaMFXyZhsqyrtClgqTvf8XXxSPuddHsNoZJ4wtu3vecJbpXwrUlaoawT4SyuZEfc7U1mV
TUniWFaAK2pQWG2nbvrA/g8QMgDFK95JYuCEe1QQHtxcigO/OIjtaa6b3APL/vQZpEQDPaFF8mAM
QKnGf8WBT3NZ6BjXa1wMvRB5jE7EnHqnUhWMX7Tf6AvcCAB6dxK/Jc24RQL8VNfiqfapJKv96DX2
anDwE0/82poCJeOoGpdVz0ARQWnnmxuIvdW7dxD393twO1zLuMjFlGnP2/TlPOwJx9INWMoIwJnW
Hg7/BSKMGEW8ggZd76QPNNj9dhLB2RVQOtlUHOsRCsNIl/qrGkouJF9HrjGCxNuY0QAKFQ6ffrG6
PPv/HzZMrz94QaG7lXPqYXdQelxwdNwgLNu2Q1/GOQ0eCojcdV6v7Nd/OlOYdbeKMpAkcyBEbOJh
XFPLo3kw4mRZFlVrNzpNk9vUG/LwUHs07TfTGUi0Q7bPcpyB6NvKShaKTlId7kPIX+3420EPmecj
Hb9LdzaWVpTTbeNvcSIO5d4Dm4cnK9iGMf/hfwk15t/uvqeeN9s4qG0UudAmnDglXhQ9NEop5q+t
hfq6cEyz/OJWRES8on0s3cUs4ecYBkiuV2uC1TNH8f7CzEiv8iDB8EMdh5N5B96f9zfe1wfOj/f3
bzbS7aDv4PltXYr7HUWi1OaobvZtFVmD5Frh2qdE7mMrdz4ZQyK4XyZocHcEDA0ULqDOw12YDt0n
vd6ttkvXSS7VnO4IdhKBgdMTwB7wcVlbfu6qB+lIbOFmvCpWlMbUopfJ9E+u9Jqt8nSVb2lb4dcw
oY/XAmjIw4+ZWZ2QdH4TuS33JF2zXOlK278Ltqv09+njdr+6I4vzbuVP4R+cg2RZcp+2RZ8b5Qak
fjANi1RQf2rwUTxfSQt2oSowhrEd12NDpgxFCAqUGC+pEdpYqg9nscKRA4oBA/KTtZY08RmLCMdw
Na4l4LCnIw1Gu4vJu/K9wM4viNpKbg9D8N7WE2k9tWzl0Z5md0NRK/+X7du9cuh03W+099I0M31l
1/gn/FMGLqmeN/vUnPpNY+QXLlAUGciyHrthc2c3fh0lRZ/qkoCuAOhxGBTJheop4xAGYmdkix1v
3/HUDJFhCIbhS9tCcn7umDXAgm0L1Aeq89wuu7i587VIgSuMXhkuA/OhXtImmyziI9veDI5nspqY
C2GAE47TLxuPZ1nlNzqw7CITbkCbEe1m9dMcXsqdbM9Z5ZqXbNupywtzXNXwFSVN7UBctqwh/0mx
9WjViAMHk9RvwHoGYlFQz7xDAvlU1WNM0APQ2hmD7RP8I55dkEjG/LWNub4tDoDdz39Q5qj13NDb
hlGcoL0oiHRk1XYqY2B3O+e2RdeRBeiShZK4SAIwQENW+qo8c31Yn6ZYsCAU/Vn12JqQVd0VHU5/
ifee1L+FHsN8CLt4nek3zaiLMrM6TGxwEcnJNHliDKU32BiiyCIhS6wgnfhVor7KoiHhP+pES0C9
uihmk+wbufQ91K+/ymdxwMYMB7j7/y0RPU4zPAvwOs8gdVu+1UqgxLWFvgJgvSF9NCur8/OhSy2G
ul6mlt60k9Cri49n/1xrR3t3YnxAwQpwTVqDR8NnMWwxQ3q7EgPBRYZ9f7xJoxmuNFRXSuxE3F2B
tIF3bax4qseO2TJmpbVeHXcPAmx2eGvjNG4n2wCCMgYdJ859uLTr+ROAzBlsxZcLvHDuyLb9vHjz
EFPMM2rpnsVJ1QeEIUCSLnzYGTojJ0jXgSZWGwKhJIWGgHUQ2k8CVQbhOKNNzNg8EoNy+Q9F1bvb
UtZNkd7BwTq+VkXqcmxPsfCa6Iz9lT79csq+S9Xv4m85yo0afJd7h1dt2kcwaz3h2ot+u+GnjMa/
lBr4Fe3B/M67uRJRUtTFWS/lLj/BMgf6JF4xQ6cBV7en6zsCq2Fjc5i3N+c0bSgNqV30nDMO/K/W
/mpdDZrZoDT3+EGk6G42ZOfDecq84nyTeldD7VqmW4tbvg2Dsj01dHji+7apgQ6S1LTg3cojSLPp
YYQ5P2f9/hkKw+Jb4HLSkHPG8jJxY//+HA++/2MiTJH0VXyOqSogitUK3xQJkT0WRBte99YDQYI0
GF/NfjnK3fprtGALFQgYeOIvSs+Ar2tOp8882hW10dE+0sdxcpSynXOK1r4X44MBvSnkBHvguszJ
xpKcrgi40/8/9IuirA8lFflo2SYLNc5j7sjwgcecSpuPfE65WtZuNaqj8DIVBWcqzGtDJZkla1X7
UdI8/FwjrxsuF2gAyhSpP9C7wN6bvZgEXjyIFSBYf9bJVAS0x5sXFiUMFOryoF1sX8gbJOAyacR0
PhRQkbgGVDYtIDltyr1NsBCOsWbYi2eY1uxXv5N3ZvByuglvaE7LQSFxuaEpbtg8xRJtgUjVHmo8
/dyodKl0XG1j+uwHnVvKWTQZebHrIQhhc3w5YCg22qzT8T9FCNsWA1rT3ZM8vsSz4lUD3Tbo9GQu
FcUOY1eh3se6VQxIcS3vMDRUvxFzXlQs6Zb5DqlBNjUTvg0OcoVDZ88rHFY/E6yy2YuKgOGQhia5
UUPgMDXA8bwYqddiMxSKiB8Seoi4b1b+tRE7qrlQQN6qBrQ/NCODOI6Nq4+/SAN/nyHtGfiN79C2
O2IFKvqrpXnFhx+8BJv5IEKzuUtFtVh1DKuTs4XVU8V4+Ggao9zoebqtd6T61GKRMYzcVST7+aIo
7a9tB0BwkjhFPN3FEYh3f1YXEuFjnbUzYCmYtLbKvzOYd1Zg+yJ9huVasfSrCRGeawR1KGXyk695
29JSqWR9YmrWR8eGYIH3QWNLoxugM5HJCDVW2wXievSSOmA750X9tWqGXksgtlCIYjYOXIJW2nhq
PSO++6uRG8RZp5CtXs3nPTWCN67BRUFLHj7sSAzxEh95gqe4wW4XnznluexAahCJP5enIZUVwPkv
pgsLqfAH2MBHA6a0g8wdLDEDdvMN5Tar+Mb9SHMSdnbE2qVnQAfvFZjKjsoMBSh+5bkXgNf282Lx
/XVa8u8m9xicbtBlgrCdEtZJXc6VLc0V4og4qKxtrfRpfwBTfZkp8ZJV5adAapFL/uQZ5EDX4Z5M
DZV3ehBIjfK0gPYdwuEZDJ/e3L5F5ZSI8c0Ewl16QTkX8TAKVAfs9+JLgX3S4JXVtqhnVP+58536
xOguYEocbQQ96jt682TMA3f2T2HYj/Te46jK2yXJ7QlnDAZC7prA00PTqy+msZgrxT5ocBxob/we
JZ+K/DRfOtcDgFmKEZz4eVz2K4Jq15VgIHlnS9GOYUjzkulH8awsb+uOegQ2M4ZBfAQ9CI1Am80r
7lViYJAwo5UfAePgY0e7MseYDC3xL2/4os9gLKORkUVMGpYrbDEOVbHnkOLyRutKilRpqA8HrqJ3
I/60oQNt/mviHn39A73vbLYmV/WZXVEMkozwTcNnNHfa5Z5MvJKQ/gtaIwffm93oEN2BuZq8FhDj
6NYqopqJNJWH9ComrDYK1kPsQbE0m2Qpby0ZIohuTZPay9oDwF5Elqp6mp0mI4TFRiOPPyudP8Rm
cmELF6vqGEpfaPGNiKAIKw7JGVPUkkFQ1t/ghxpaMNBH+s8R8f0lcjDiLHtNnq6hAhvuD9BwuPIh
yjzyDJyAcOcp56+DWR2nOdX7Ue6YOsgFiSQF/Ftdb1WzTKdo39esMzW3j56hMzZpJjwcUDKXUT+3
wjwiUoCQPubQtapyuyRzN9RJdJF9ZyTRSr/5hQ4kVNgkmWghoinf1mv0n+pud0AdJ3JpVdCrKemQ
CTzSOEUUNVVkfo5xfvcUc21YJi1LUWnQXq443RSxokp8QY6Y3eBfviEe+CFV8agRcQdI9RVyn8tU
w82TStZMcQ6TP1Z69hzsCdqnZIB9Dxe0lzr3OSnyfj9OSqtaBSb4+yGy3rUKT9g1csVue+Cb4DzA
+MevTnCy2+Tu9UCNfZ+5ISJMaDcE3DKmXeqv+O9TpwktORq60JixBNsslNDk3VnZhzuM6BbA4eWI
3+cBYl1r2mlRXnoXFCxWSZlttOf1AJXHOkV7Pg93ZnsBMmfTLfm5HxKHeIoR5v2ieJKxVVszLC3T
XwEyxFKjT0Yr0ei+pCXI+OK6teNiZsfY30rpUobdOLr2NnaKP6f1Qesbv5Q2eCjmMDliNnvzvd7x
wDYQv/K+pOANCJ0OrekTZ4HnplPolqH2lJnbGZpNJq6JPtWez8Sz4qI7vif3HqeTHzzpGkNZFAVM
mrsvDtGmps/62V2RYwlkAY1ptbMbQ1cG8c8QeW+dUNvrziAjR9XzXyXE68exMJKM8RO5GslIOh78
3Qd1xgBGwWaFZjT1Q1hy3j3L6z3nEOxbxufTs+Lh7t/x+ALXNB9+TGKdCo/vU7+VpfqXhNoDwqJD
UyBXkRo9MqZcwRHPemuOEI0XIXXYL/amUI8oBsjikek+DanP/Oz6WSXlxYbiSC9H03x6DVpLTifi
y0Mq6C04DHpYOkZGQG2qgu7MTDUy/hdmo6f4ZqKj677N0q7Wlk+/trJGMEL1FU5nAQwz4IiGNg89
PBeVVxxWYZk3DZEKnaGM9wDicjnaVUQAsGagBjowPV/i+M0/jF+ChpFCkLxfnTaMr/LfSHtCEYtu
K22G4jRkPIUmexMSI+pu9VHUK/ok+pk5kj+Wob0UXBMkbvkUiEk+nKdaCpsDrk5wBCl+TMaTlro+
a63rvqCDwJXDwTC+ksyALc08rmD+wlL8ek3NblPzkRCzcqqHpBTdEzPjWUmIfRQOXIj127tNRglP
yyR7UVFjBpiHMcpuHsCP+NEH5Z9nyc1g+f3v+C5vN0lp5IohioihBgx1tdPZ5JJSFH9g61S/YPPn
hJC8LzuFXnpyZbAnfyG8NkNd2hBIoXj4dIlHWSiEu66ybBd/h+Tg0Fg3dY9Q+oYqQN7zfnvRxRBi
NIUOkcNT13ORWT13AXLlsXSvClEIh/DV0Z6MI853ysNiZ29b+4Sskfx3ipwVcUGNdb6r9xTFKwqb
cX1R2VknCyLhT3mAqZ2k7+fVLrvPY9uJxBP6Pz/L76Y370x2Z5TiYWxWT+Obl+HpvTSccph+lt0g
1CCVRTH2+Lfs9SVMNSji8EgFrk/PueCPwwIVnI6zzxQyh+KmKL9hD/HHVf20oNdhQdSErZ0f21IS
kJdgJKWL2hrfVev4ed4CU4qIPe24MASpA+P3M9KCbkVp9GaWJXvtBBfzg9Kj/TpTsRY/6wlQbDlA
qyRRo/IeIkSh6C91HjEBpZHEzJXnv4iqdNV0psdVtcYIT9tBlKxztUg5sxZmkMSLzvLtX1wyRYGI
OB1qlIAgcumfLVddUfSbajNOitwr2wYfG/n6YTFO8k3kkFHV1af6OVnhnG1Lo9xHLlSsrTR3HsVL
CSnaQvjut5i+jxJol0p4b4W0zokNhomJyA70CF/yPDtLa50HfFOMb/mH7IMIP8ZlFuYCIZd//eRq
uEI/LLLKFdoaMf7kgqupo0jDrAUxacsSuSe5bF5rxQC7sPCgEstB0/94KKIrNPfd973mC+SU8FMo
Wuq67pEwSMdeHGvmfKvGUG47OuGL6Ry4I3po4Np4GXGagRPqtEuSTBw3QZwN14L8dMZqeucM4FaB
Lyb5P+tKawQs/joR008kyRt8W1JeXWjO0pT5QjRE5mhyjFgRWJtxtCsJ+lGb6xNoezum883QZNtW
NC57q8yMinx8zoPQqZnsjKOn+0SpY9xeKxZfiOEDMAmDRUKKkUxB+wpjSIm695MF+zaCtRl12Xio
XYqYvBnt3sKdNE4RtRs5ysMcSvuIVbS3/5lxUR7VO7DdOOwWXvPpVRgZ111hmHvtks4QMJIbEaHC
IW4oz7lgS7q3vc6hlFzzcvs61tbpy15V8SJX+FTw18s9IsqXyV4l93MuqqWv3vgWIyjnlhFVDc6M
Rmije6AYD8md+qG7b3sMB/VhX2EjVCHMkWm3exdDTN7aGfApEdOaHrv7l6GxSp/yb/zz7a0kQuaB
upYx3IAgWIdPhY/deyN3E5gNG/1yZY1tipNkBt8jkfnP4w42xGuVwB9aLOM0JCbgkxnFYeYJNU4v
s6WyyyHnkXrRDWRlu+SJXiGyI1otnigdsdzHZzzEZLqTszMWAU+ZHVJx79wAyO0Sm3xQad4zD7mj
c9RJwqS/uxkLh++i/Zqiy/UJQiGCp6BW4YAn2wgMgWzGjmTlp0joeCXz774VjQP1lS1/7fjPjhLi
G6rkOejlmeQB9j/E1Adr69rxJ8GR2UPKnYHhr52odxO4ufqiUgtRkJJlHiw4os+ypIZ9bkrWSNL5
5HYiYMHVCV32sZKfTalqcAWAIzGI+G1MUWTJuelCMqjA1nbnaNmUEvrWkLGVsWbIs2aBmO8xsnPP
Uv4oQLJsJk4q1vtq6oVFDIi7zUDEmy90hwD02saMaU8HzwbeeSrWWPpqvyC40hXWuSU7gUGLp7Sm
ldGkBiFdxF3SdT1oAAy1f+Qsz/aH/0L0vVwt6kbTxo2qXBwJmriJ8+qytKrwdt/dfEv2COOusEEa
Yadv8np24Oslh6AOwF1tU2DJfcyUD+76Lv6zjHiZYKA3sve09KUoQaCW0HpNoTXkblAEPLvG4iJe
fSQ+SMDqYxHQEy6DoXAvXpdAJi1Gq2ZjqBeo7Ms4Ht/694J2pq3p1TIiZkPre29GqxDTuHcdkRv3
fyAB//xNKRBjp7O0IJKgn0qEucWCIKBIKqflsYx9zuIQH18hiedMI+vmk/M9YeH8yXBSShfB4gSp
uoMfA8oJlZUSzMFQm2CAhWUFNsFcZ/cg9n/q/bvTW0hwcupIFMdljxwfxgRgwKIOHH+8lINIyu36
L4+CUhvB0GPH+VZFL7yIXWeAgMlJXvNTRalEJlR3W19UHw+RoFqyxhL3IXK6H/c7pMeyKKlFWOx2
sFsW3cqc2GQUnceWZg9cpwg284S/Kmoed/AEPA1dp3scjzKrWdcvcEMs8GXZuPD+J2SSoxHd6Ts5
3teJitzLfHNwJKuTvP0Rku/r+x/3bIMC1S/nlCC0tdSQAbODnujPoa+D8Wd6O4t2kC/1sfVaGO/d
ZjZk0nuG7+xzZNmLSM/wW+polg6OcHUO6N43FbDRWXy3sI3DsQUWNd0RIDW9Oe7gFKoM0BV8JEBt
kIm6faaL8S3IPZRNEfLsh1vvhxcSU2rR08UPU0DFhfxoYl0lXYrUW/Ye8kgALpGe1vu0Ma82IAP5
SZ0yttngbF3fYOMcNRYMj2YO1Pj+SLhrjW2myaII9LOdTnG6/5b5UXAKEH75F3ZHL8QPCrtQiJGV
lOPpUxrv0qe1fTDQXF1daK+7keFWOW6V7nOFTrAwaCy0TephTaRzAGIQjjX/2kaJ7kZN0ZVq8m8Z
IpzLiun6WeBIZGnbgTOe3T50StgoY8TL54lL7giDASiGW0vgbRhyq+ae7rhPFWmHM+wDFA5rIbdP
b1JNiq3+VEcd625TIQ7CoFr04z2Pgcf625YWl3rq9nTfHOrcIgr3NXIrKOg3iwYuZytwUP44bLnX
SxcccjfJL6gMrE4IXJ2SIe9jP9vHkH/g44/7EqiPaiiobUHj+nMWe7ezI2WXykYQrB3q1pyArS2L
GNFipunpzf9cauhZKe7vzxcRjPcUSBnzZx3xzGPLdiPvdD+b1rN/XWBgFUosj+OJg98ximGsY6c2
fKm/972Mwk7LlJsesKpur8NlOe6datnwCzXi7QismXD65b2ztL+B/Oynf7apk4gDFVQoTaP3V4Jz
oDR6EMviQYG6jWcWo+zkDTxEw3mFSZfsI4w76LKZBhY+UnJcnH+58lgoLw09IgDn+281xxWtPtFA
J1J3rb6Et247cV9juAlDWmINx8ulHK5HGIQAm1v4fsrdjlKStIZTVOqglmKM/4A7mH9rJQ0FG32R
HSemV3VeFKvLGZ12RhH7jQ8Z8y5Ryz1UU+W2h6gxhm/DxzQ7RjktlBSABeq9HLWQ8xiVph8iBfkS
Eyn95VDd51VnTSwl5zGXcyzvhwx1cdtAwru10dEEx4tkJEa3NcWd2ho38KyZVfJgprrDGZjJAKQn
ojYIstT3Gafp1bjwqkkTAS3Avq1aLouda4K/kVxpP8PhiLgI/AGFAIyFLOy41UJNgqp8m6n7axPY
h74++Ft+KsK3AiFnzVyid2zMaCVM2efBZFvM8t9AouNrHy0Ch+lFMDT1BEvxM3G+7RE/fUod29CT
zno0PmL5sgXwKaYe3JubPlKZD68OUuLj9X5I4GqllzhQieyUpGJSR6EzsP1bWzRFn38YzKsoxS4R
5tiDrqFpZYeFAbTFP7K0Yv9hdYdAv6MlY40d7Y1l/NGHT3QjsZwfyGZ5OMcaRBj2GSJl5R3m7rJR
CQOfQd9kntO8eAxwI32IxMR5uU/qnVATGdUqDC7YUWoo8AcecsP42BYWJXwNbJxp0WL/YxPunjl7
XHv81gQ+Y/Tqaxjl2YhFrIylFBIxzV+9rQ/TdQxcbXFs+/oXQVuowmer9BndvKb7W1bljf2AQT2q
L7siDBnJOY5ja1ka+9TLQL8p/KaZ69SQz/5DuGGhH9dOaAt2MIikXfwrgtRUVnkqBtfxIz7MYSqF
o7inidVLj2r9I+9UhXf3LYY2UCeNcZoHX4/MtiTdPQoSy46IzGck0OwDR8eC374szIcez+uPexTI
XHh7g9xGZyhZibU2mBzFWcX2Kz0ltroCXpYWU8JIZdcDJf3O1bmVH7ln++LKu9uAKoAZN4nHn3Qe
r4qGajfAERxVyfqGZHarKDwYTM2Ky1KXX0kKcsjDUMYl6Fqdw8yR6AIOBhCm1OMb7d6l8foafkDo
Rxtn2wzrDznayJ0/4FHdtQrO3ue14Q6rQO94bPPhdDEAqg0C2HHxOFrvZXf7n/8Rwtjt/rpz65VG
bnB7Tr4vMOcyhZI5PyVl02YUQ5GX01vm17GL1wXcfNMaQJ55HYTCFviUnopDy7PRtvDCdnJzhIXU
TOC6trJaOG1/NqUslLtM7179tLi6Vldah5+QdXmY4zVeNvXOv3Ct4PMDzCMb+OdJgJZoErQulXM0
DG2aD7mKFD5P80ljmrGzRQ7U73ijcJq+PLuTsMYu5ThiO4wZM7RVVBstLzAp4Zl3lOHK3+xV8BRp
53CDMwjP92HhowKDi7S5gxRGX5G7+qrmoRsIFBxESNk2ZjCOzFgB9eb145IkePiIsuoHpLoY1gAx
TAGVn6R5D7QbHDW3Ijg5xEHUSf6Zt4x18HpPvv75KtU05DjqucsrwTzz1sT7f/zfydH4n74sLi98
xG5Uw3NJ9cuOgV02yreoT5YQLRS0LAS2vngIHy1rG3BaU46jilVT42x1g6CfaBxnD+a7KnXjz5V2
uYMpFmm4fjhcTdFw8v7uul/e9kvqxB77IqesLmeyrp/n6uWeN5JEIJskERbSBf5lBhAIeG9svtEy
84VxVEOAy02906TI9a6qH0pUbXBn4f0KUwnLkvS1zNGUbBbUTxzot8KE/r/WCZYPBYFsq/bfxymE
ZIw55aP2uBmePmNgEhV7BW37udGy8vmZaVY3tNTDERach1K6khJW09verXV5wf7rpHBnAa0V/2ct
ruZDSvOqgmbeFwCZdALyGotDP/FcuL7LND8kXOwLtgJBKxGqhFS/jLYN6chCh0QmEmGGaYUsxfoS
uRapk/tJ9HCW3xQTD4IkXqV+Cnaajpz1S/1eK5qwGpa2Jff+aItHmmcgXvZN+VyNZdNEkMRnOyar
CmJrcGGEKNNANhqQgMkoW77jyQjNV9KS4Xsa398ICYbNFP77T9RoCBm4I8phACfZThxMFKGKjR5X
3HpdMqAT0PeXkc6/8rQ67HSkfDustlbRM9oTsdlo6is9YZgUrzXtBB2CP+dxYZgRWq+HLrth9Co7
CwqeW1rKTsbjME1xJX+S/FAtuzgzvZqDefgOk3xTpk/y6v8Hu75prCqkpuePClRZyGEc720I1I3I
y6p/gkEBI5TV5pnHIYdl83u3nUPkHWLcihvCLkeGyuaZ9Y5Ob8JXJ8R/JUoYZuGc+5aKHN00dSda
/SH3W/+4U0OWaar6+dYwQnojnFHLDCEFIX86bdTCLCh5x52T33srNtR/jaiCF3skOPFWyGy73W+E
qIup5rYWe1mwjQ9xT5JE2l9j1OK5hLHLXoKVhgoRfmRHJNvkmNblFEPqU/2TCKg5YrbMgrLvoyJp
Z+1cWeijHvyzpa1M0JVw0vA010EpSqaT8Lt2/MXF1s9MeeKyCrzGfYTbEuY9D4XXrrlIIIW+quYe
5sWK87Kgy97vO+Ip6uDJNdm2xwhn63gae1cV0umO3H14yF3hOF3WsOnu6xhSC6kYOJOh5KR26Stp
vmJRNxFo1iUpFUCoU9ekO2IMZAAT4hkvQZy1pdQl4zOJ3uwa8yeOZvGK5SD5QcjJ+G6TQ1kaOi5+
F+sK2v7sb2lVDhqYEg8yl1v548mBdmi+TYyViOlhf2NCOL0mu4W3ur8MAehF1HuQ1ONcj0aoAEIB
J7+oG/u8U+HNEUwby2GXSH++qkcux7/3D9mcHHeRNPmjkJAk0XXzHya0xwbZNSAIQ6RTjFRzEvoX
LnFge7fsYi04NvkBM5FaHMF/xcSGooelcUiKAquJP1X3cLBG38xa+EpfjiNmGXY+Gp4Td9YO3Yqr
KnUpQKQBwMJ/tnWroWktPbwD4i+6xzYIid2hLvBgZ3A1YYMXOEubWcY5w9/kM947h4CPqXPudJMO
z1/9XbEuwQaEEnLJSQE7CqIg0UEuCZX8e/jSvZHqoLr3iwVjnCdmn7jkH0ZrTGThXyw2gAcoIJ1+
aLntjZ0YOSSlXq7Fh4CQTXcAMpru7PkWE3+CVISVWFrlAVAehRYxrvbfJw/VJdqc68CV/OV6D5S5
Kxpczk8Gk74zFW/F/5IG5DcuELM+/zxcLPql9JA6+exIPi4EZcEan5qGO0WBn2+3ebp/3xhKcDsY
nbNzAKarDWeX8mdPhRq2L2edwF/UJdG7bO1/AJ2T2cJp52sdnDqh5kinRmaOYI/71cu5WPUnH4h4
Aq6VBQugF736UTCi+9RhvX15IST/rV50DnRP0tt8mqetWKpaUPgRhHAViTts23tYUHjetd6+qrjJ
64jQ4YSGIVr1c3PbzoH3hjK2+ROIaVhVKL1I2YmPskLR0b9YDL/eSsH6oCLNNTdihQapLTr7mLK7
Bs/0SZAmGOQ7J5IGPDzKOGHDU4yyk51nPn/AacuKE5JqsMoyuZ7TeVpWh6lSKIaXz/bOZpXmBHug
+OPxkuYIF00p65w+FMrmC0tLhGI4LaV20E7TQaT4NdbzrUQUv5ooYSwem+yXzCyuPiHJKGXT82Zp
LodlTeYcDG+MsEtjfrB+q8eg99QqUb8fk606V7FiBvxQpEjXZrP0rAwUdqfKJtouU7Q/wELlqOiG
NRNaSWzAbAS0jI68lCPIs+dmJHE35AgQ81f9dVWOXGIklxzQ0eLxyxllhseUAFsWdD5+PIdwlvDI
ySKyvo9CgjWb+tgsSnZstZWqWnpRH0nS9e0bZbyzHf7ckuOFdDbL7YBsV1a9UU2dAXEYyAwaxjtB
RDx3Bq9mksIBUPH4x+RFb/45VXikHB5CJ3oC7GF097SpYMbM2vQvYXBycEUcFuR5ISZbE79OrOSy
aRtb0kigusNuDvvNHYYiAWwdLI2BIl6ofVNGxOIq7iBtgD0N+U0BYe0At01begVA6ERcCnmfYjos
HR5gphn7dReiYIIUjMO5qN/99zf4tg0/oTVDUKsRKHelPvqG3wqOrzlOrzMEliXe+n40wsBl9UxT
uTw86skubJfozoXYZa3wsNDWkjcZvHxyppMeqKXBSy4HLMKCndJOj7n2GNSveoDm82G/W9n6ie2R
t/vzXKC7TiOsoznv1igSL1DyxA0Kzho/pNdqGwIiJ87K3aVQJ11zIhpcsnBcZhGXDuJF8/k/3iGa
LrbqMImjiF36ia5OJRXMd8eyOJ+reN1Z4VxF2b46CbF8POpWAVlu00Rmhy3qP/u6N0Z7+IZuJuQg
3B2hvzaM3YRSGvoc2LvjLVmV9BTAOjw9z3j/p7CjyfmfUhOdifsKyz1BBG07fYwiS+nb5VPpNFTM
5BvttXj6AR+qFrW9p+MbwHAou2xEIQgt1dJF6s7eYBrblbnEf3S4uBY3Pt1I2DM1I6A1/Bd3gPIr
OnI7Q9B97BCmRzePX9+7uxGYv78yLZmDnD22jD3AzfK5EKsG3tUe6doccXh0M31iyWiUaUrXLGo8
kF0TPvPwi4otv+B6khhTL+K+iimOQZSfIthh+7aYnPiTu4L4f6clVELbBis0D1xCiEN7jnpTlWBf
Wre9dTvbXI3fyfZXTl9LJAjPMiNhJ2kyAspz+PAVyyyS+hYr1KZbcDvKTKTUio5i5Sv5EijQZM9F
eBtcyqpDG1humhYgUciKyvVRVvcLvdglWaOeykdFE/KhVH0xpDNnbP0N5slfiuclfNjKE2lqFYu3
sg4krLf33uCQnFkytXiNv9J+R4MsvbtEcl+ghb/xxX9GYLjcvhq8G30FRXIujp+sIY3q5FmIh6gr
3/DFUgSGZlBonYjms0ttw5NJxx1Wbp77vURqYcB1P0+X3tTfh8sYsRxfUZGVI65xJj8aZX14Z1eo
RUAzYlZrvfLYBZFH6ukRDJapRokr6t0lky1m9zOCD2sdU3J7PVkiyr85/AwTvbD+zxS6D4E76/zf
nvwsNEP3t3EhitvkmRUp8tWO9NlukQF5D6KZYbc1yr3nojCYwVbKbDjBuhu8KFlpacdEvr7fIJv4
8ZEqyn4eqPCvW8OM3/Ok5s73177lOIexVprfsPLh+LHb58UWNCjPvGEySGRqCjh84je6SKbz5XhJ
qQv96jMR+m/KXcObL5vjJanYCQFxsaIpWKbDiGvoZMShgh00iqFtycjve6BaYlLWpP4rwfqWpYvc
ElUDLD5jXNeg6fTzevjCYVNENF4F87ji70afao7IuM3DchgNnOPjIT7T0JrryRNXAuDr9vf8v/Kv
OpZvOYIc5TP0+C0xnUOZ3AvuWlERc+6HRyPbvNrhPDTQrRAAzNAQmkTofxZK1rq5NQ/OKSe8hupt
pkV6eAEzCCmeQJHIINJoapkhZBEt6GIW9gJXa+jXmYW7nnRzGtySptB1OlRn4IHcJbRnyykIXfmN
sutVzG1P9plipackTsLpaWvT+pJWN+vVfUp7nDSRX4Vtlp4H7BZfRQD8RIokwjqmXx3HfzuKRBDU
UsmmShtKwluxql84ZUb+6vVYm7AYYEAlGWYSFspWbIvY6TtxnncVEghmQghHZHojV3y+g3+E9Jo1
u3I5mLUXkjSyHfwaxo6pqPLQq1lIKLrsnsaL2oElAP68AuiB7pqNMCS7WqWHBXHteOmuG5v4QYse
fXN2hhqXF1lgSlHMdLe92WKdL1OcV8I4RXLG9ah+5M/qtmRqaOScQXyWp+Et/ZI05ZW5FvSBfP26
/oq/pekVSP12cxmK8iud/5818A5KyQ+ATZ6UsjWpN7Pjl6LBexFMJo32/WYRVWb9uInoboJut0iH
9V5zykIYtX2vrf+hLuoi+ufE7TQqzo2GlQsXOwQ79PfjLE7+fSHAuH8oAe81C6fXz3LW+HtNufBM
1mtZPCOpIXoA/NQgRHkmxdD8zoskAI9Meu3IyHBhODbfXFpwQn/K6iZtpbw+ulcvwohWXR3TpTd9
OeW4e0I9/AvmDuxumNVDhXi/KbAZaSaJN9f9yiB8GHXH+k/A3fnnNJuUaWFecVuR8sgyLIGTf3TO
ysvxhHzzDS2A8smMOnodu/7pOzf6D4YYoCc7HigiywLidwYNmcS37usvSLnZb6IhMb7+5T7P1cf/
tx142KgkN0E75eTZPEBkKlk18evMEm0nUnXtZ6sV+gBYJ2P6osmVRaVgcpWIRwYxziWjDCXeCchp
Ak4Mqu+TGJ/AoWmExKcVLVxMfYZAKUZzPdxLlAOguyPTIqkHUksFjkyNjR8Gqycx+n3fdTpAqKbJ
KE9Jsx+y/jbN8vv1ITVk2GvtQOOcL6wLqCsf3xdOvigNEOYLxc7IkRTw3HEUESHey3Lxq3RISZ9I
PIta9rlTVs5jLoCI+o9a/YwsesbihwZxkAb9Nc7xruA5VTG0ZOrbqYSCzLbq4+AtalC5T1QmSCeW
TZQWCMmol9IWFvCs6Tf/xIoRFHnULXuBLG4rzvONcj6YGKZC6TxS0AcNUSW6t66DaxAOa661QP3G
snG4kLIbFw9U10Vp/kEVcEiwvc3A4Q227j84c0EBu/lBHLazxLbntNXnsNAx9LZh7WTuFBI4lD92
7FSDVtVwFtZOA3a6UBQeL3x5TMuAPqu56vdw2f6nyAIZUPZWpA+qhBSyWytMV6HbarKz/DM9XkdO
W/utdv78zO71bCm2Uaorcg19jG3iibnMp2m9/bltYm25Mlt7gmvX0tLEZGTwpVcK+KlmcpyplovD
ILPlIsOuB0r62myiagtj+GtiKtSjy+Yofz7dFM/qYApCu89HTlE3vso5iD1Zsa8S3BbS8hw2+4eS
eH+OARjHfbq+H6MLwml2TcaV3G9w9/6wH0QhP0R9rwMdlBa7E1+i1DxOzSJbTuxRHoYthDEzIL5Z
Ej3XBBaATDFREvCeaXXl5jja/KdnfqE1SizzYhDDfNmlxsoGM2j9/idk+iCpxgnbUTHqDsMcPGWo
cVYwk3q9M1Rnx0bmwiizB+QDmFeNhJEnvHg/ZKBI7G3b/yZGWHox+P2LGYwvJ+AZ26WTNcZ0VVs9
NvLMgmv8uxL1Ri5OKJxBln/4KXOUwaK9wLf3wnaZnlgBuMkg4u8CSLi31KTEZk8rL53itQ++AfNh
zrIOBxiMSDn6QKeZvLusnbPqhuPP2FpZSxJOcu2kNR41ODbnPjaOCxMbUdzRFcZw1h8qSUcIQPsO
fDnFz26XGE+ax+fgl0gBQ0IZFmz3JUTljGWeSTch8OCbG5tP2VDg3BDSHIwMLoWi1Ay5MY3uNj0n
scGyTy+lrMA7nGeog/QcnG5PVEHf+BdzFgl8qD/+Hhtsa60ccyzMWFHZArmZPIAYQQALothigA4f
juFz0f/yVr9Axv3SytedP/SJ/cIYgq4jy52aoJckGTCqax5Q9BifWCCQcVtSsRW48u1mXELw91W0
bPQEsJFh5g0bwfvhDNCiUZw6N+Fz0gpOIfGIAgpoDncYAEPB6wWHwaL5D9WxFp/939fSzWStlF6Y
CWwhLUgELYBB7rnYzIwEhpu1x4lpaNF09uINdV7qt4r5YRUr2C6zcl0SYROUTvFPc4/F0QEhnvyx
hC6WP7TM9FM83NCODbBjhLUk4CVNdAY/VVgwjE76v6TmFq8oMC4obJtTJcYfdqUK3a5X9fY+IN7h
AqYlLlCzlxBNSx7LQaYzH6aOPj6giXtwXliRspsXHxW92DrF2rlrCL3euR1Tf+jreZv0b4O2uEHC
aOBlyEBjTQ3DMhtmv9+q0PJ/T4LnLe7oY5p2jrZeXW4HtnA7pfCO95fryby0rJaiLPtSSEa0hfP6
Ko3Kfk3q2QBXc/deJgTsvzt6k7t3CA3ADxj8sS5G5SgUydLguKX9eVylOO4T9bT4/mp7T3ZsSaZ9
3OFNHnTnEDuItffvjgpEfVQ/ZOE60P+Fv3Tndjvsh7yfwC26CdPO/0W4W0ijjKv0xeZl482wFRrv
pKds80ZbyaDqjIu95+UOGDcyTWBimJYJc0DaREupqbwbaAHIPUCTvGLoZfgu5L11izrH6c0jDFY4
XzNwceFPbSs/JXw1APquoDyQajViBlFO7csGwxGSpAmwd6JUsNZgFZzMzzFBeFuFuF6x70nbyULi
RNW4HBUBxNqZK7b+OhkPo2vSGfliw2fhTQwbN0F0u7BltYEPWnaac5/yUx+AxdSQMmFjNlhFcl8K
0EZ9r8UJGrk5Q6/vwJ3wtKuwQNe25VOZyYJlAt6MVOsWs9Kjt97DAIHW5XkrJn0uDQqtW3HF1SE6
5m6tz8M62htOf6GQcDt/8qLWw+eYTWKjBA8LzWYQEh1NQnAES1CME7lueOPTC6scUwuXKPPZ2Fr5
TBxJfRgWvJ9F+I+Kx9rxBSkLkXovoLwBauO1FsLLOG3U/9jHK0YoqQAELCR98cOZT56U7A+7LqKx
L+9FOtldrWTO6Pu16HSKQCEcscANWfkcnuOOs35OlHVyJIehscmSFbI2iyOh8Dv+piP57FEWV627
jmQRB9SBwIIYXxXCQQYUOxpoDJz+6lGNikEeSe8RwZVpFyI0CzPxetEuQ9DgusaKGaCLaHCDeka0
KfWwb9Cd+4aftY857B1Rm0FPvSpPY+jPMK+EnHAW7BAjV3IYuCh8eG4LiOmKtlAo49bzp2KOKoCA
ezJ5SsK3pOa2JzI8I5Ls3iUpqVIJ+F3gneHZimx/WbKpUZkNcdcplrOdPUpKiQNXQcNbd/PUB5BT
mIdFyuktCM+vkx6x6letkIjqZ3pb1+IhEynJTez1s1ZkL9hb9yKgTop2OTbRVJvGc3MvjI3piHCK
Nm1eiausSo4a7LYldJ1hAkOHTkeZ5VyQ5/T/wx0Vny+TbI/W8fziCpyySOCQhb5XDSHqzZfpgCrp
uP3l1/xnd90qX8C4ubc+RWb1UxrbsApdC55Ilw5jYMA1M9O6fEJzN7td8eSBWvmSBXFRQluxrc8R
NiZ+nXW8UYEup/q5vB6QnDk+pBxqeCwimRlvameXeQkaTFnih2/y10DOvOV3j3L10DywN2tk5MZK
3C5GnxXuxeAexnNiDwqbCf65iCO64gtjAPrNYo38yiMPpRQzJkUCRN5E4mmWd8NYdiMyU+ES0l3w
FcllBqAdZzidI6gXfrHHzK6pUnjl0ZId8xmgpwzrzfhNr5Rvrd8asp/5iX6+ph30iOkToi/fjqBV
SA+JpS3wu1qg4Xz4DX5unEd5rWMhGMS63SS5D1Sdq7OsSgyUXG1CL2JwUfVd7zHuzurEXBejEaVr
a6FwX5DFpFyWmmSxTZRPLLREDEvBJR62CAKWBgPZ1kRBaU1Xc517DBDFJMbOmMjxDeoSFBdwlbv1
EU6e2nU3UpK3bwsJESCzF4s/Iunhfgsol/zrv8+PlJ8i64yrQSRaM3mamXSAfweLHYwR5PE5Z2hG
pwq/FAvUFBIObWg9d0HSbqjPoBtNNunA54q5XDH9dSv22EGK1ucyTAxZ8HPMH61R0BuD28wIU4O4
QWfgTJlKxg2JmoUyOzRQD2BmOANHCVzkEWLeu2uVoIzYnhNconYCaMODMS0KzGSb3zY8tiCOxKK3
6tKzp5PASesjZ4iGjJOpazVWGUFwCjhXLQrV1FczwYygwOEj85SpI7h9Z8xW1UwvmMTKw2CD3+f4
Tdl6xx69F8plVenbHjG2eS/ZxPf8XMHrDZlaBuOZD3VFJOSWj4Qp8Hv+LsY9oszqr5W5pP/WRL1r
02CJ33L7EMKoc63L9Pxdne3AYqUJpMNl+SFmgfhcBwelKS4oF3wYZ/w9wOtlAQZQWaxyNOylqUFc
2Alam6IEdp/Q93VW4NLS6yhaaiZT8RiEj71GKeEAyhYldOgN5p/lS4xGRSaVx/Pw5D+odhMzahV6
XFfj3IjcrFucQreHDOtsV76mK4GMWbFhYQkIZ8rH+1cevUxY0mGMI3+bxAsd2uNv7/EJl/JRLgJW
XcCZPICozJYP6VAKXw/B/FBrKpUdlSd0XRI/0cNFNsx6hRRyAYdobW+re2uK9PvYFqFuV0bx4Kxq
B1ZJNFmT3N2+s3YRJ9YgRCYusD7eY1exGopk22FqO1cvTaYreZ70U8nCk6akECwhM7HuM87V0ntN
FHREcPMeeHBua05i5cOCTVIkDiPsubUaFjetPWryTNaiDZe6zv57MTwLzeYzbfjUO26pdzJL4tZ+
6PksygJTWDqCY91JY1mjaFHsdExuV0OgK2aPWoDIwcCiAWMS4QSRWlyZ0dtKitn7lkuVoSN1NNjl
gQ5xtwq7BNDo8v95lzsIm3GI6BNUzLnKXHzsfR6zveBbNN+GCWjsyyQNUvTIyTwzccT+pC9f6hGY
7gOkKSEMZ0RqbtN3HFpkBsqXIOPI5OPYjbAA9GhSe4huIXaUYWQojpP+2krrD/xubLLlqSiDu5Ja
kByyHp3VX4bUiyBSwpLY9omHuRPr4iAJwDjy0CRILBgEostxA9bDh1TYXfdRDvMsfMc+siK08sAE
phGQm922WMiB+l1AmeRjslAsFZdaiJMciCb4ggw99xgxFGTKN2jigId3EGY0locicA0I39Rf6iq1
1MHhtQvw2bCOXj764jwx4xDxLzLp64x6B+2a/q2zfCO5iMUMTrIdLr7hOIcK3Rkda9mX8Jox3q54
a4uYCWFX0gXCxZiAjYUojlvykbu5dV/CW/ty6FbCyp6oXhWWqXMnSIQPZdjjsNI2pQyY7MH8aSbJ
M8lM1BkqKZ+rmwEYB09O1N0a6Bjs+s+kooOph/Vcth08FBfJLep9ZbpsRD3Xte77zTnTMY7J59gW
gQZ8AmlabnIQKAyVuPca0722AGsafUYzR+I61WvsULtZ9pa8okEOZ4t1zi2p6b6j+GLtNoU3SyqS
vOwsA/e6Gn5pFvnZ9Ux8KNxCKz/T0A3SbSvkKbRl5TOp89YKTscXTK7hpeLJ60O/MPmWIe9BrDdF
1kyvpFn6DOcwg5VPxpFUkaBiG4RytVWJgzFr8O9umBxmsbDJPa7l8PG1+d42X4cJ2GAl7mVUXrdz
9ShItgWLCmPvO25lUFrGy7RCLxogBJkFWjZyNu/dpXx10BZShLj0fMS6LEUBN0CKPJEeCptgLTXM
B4jRST757jJNVRHE9X+4kAO/RC+2Vhg/jTzuISqYqomtKY1CMcSoiIfCz7hdRrIGWI5pfCTf6G2o
lbFCOoLJOluBK4KxXWJHVVEDYFPfLbVCPhbcop2wDtUpRybXHx9tIxpcwDx4IirWqu6SqmTjwfHS
uknt9DrAhcKiENVAMkcaIWvdPv19yCf275LGrpJMsvn4b4uqcxOD0ZFEFTBYaNgJsGmnY7m9FmsR
54qvzrCMRn3jNNxGOvyA+97ks7u2G55ZicMXLoKD87JqtH19CsXPYfCj//71cwDkgbksg+4RvGWP
6TNxsJouiqDxaDm0GmmUCIeVRoeuUoEr5ilFCfM9RChubRxy0WFNAvKxcr2fhi0RmEshy0hWzVpA
/2sBnMS8ojeLPHYnHH8ExfXyCYJWhm8EB/JbtJ5mzYRFdoLnZXWuNRqB+eGtKWSP5jlYiuWDlNkO
VMp5XqDLWdrLfzQiCdsdy7mCH5kdyDtkQbq7+ajR0pes5F0vcYWLmwCogeUOY/F7wZLwjvkAnZu3
arx2vYXxOjh2N6Dhz4v5XzAUo6J8zCzK8IGGUH00iuqvi4fyQqk7JrvEC6oYqY3HkgtkXaWIuas/
9oUVmLS1BpW7ErD3rLO5OZY5dnV/MFZj2JISh+cWoL8g3woBpnsc5cDLL7kvYWFwS/ZF9939gHrV
58UykLR7GAIu55jUDINUEAaBPvG2Eo3dmQjOXy7XeMu+DAsVx77bFkNryk9u4X6eBeyVf7UtOXek
ASgKNfQQIPU1UzJxlUdwqsMNaI7bc35xUJTLhjKX3ULAfT8LKF3FCM255EODA75+UaRsvMYoeBbm
sUS4DbVyjmiCphaN8yGzDh+kK4+NfmU/G+bQNydYABlJEYqtmZLeV8vEtTYWF+NZpq4HdwXZWhyc
E3VVh1qSvlYdGHk2p9F2uquR/HcHURnQGhLnj/7E9lr+mXaKWMnBl+8Zw4QqIORWNtF684ZrMHur
Tu2n3JEKy7uvkjmO/cVb+uAYk1uqPOEVb41oOh2NXvt9GauejA/haz4qJHu8ecQ8gTld3JsEXVUI
wROwW/gaffg9IMX36uYI/EABL/3sL70uOrVY1YtgB+YgxKUSsJyS489zJT6mI8wcKZWBxFUj2Bco
wu3z4cxPIx7jhL5hOLCoXe1V9AT97Rp8brUCBBWG3HUpLu0LuV6Ui8l5P67JRsyFRtsUbV6kHU6U
bYDfPIwYyNelqvXPhel29fFSHxIwWw9QXSeXAAzpq5OZGFkVpdf91oicD88tfh5XCMLceSEEqxgE
A1+lDq05yCsgsfc/9rRj30h/NUeci/rdBb4Id+s9jEv67d7pQxDvPbeEXwJ6ip1y1kU4zy3lxzXS
EYJfu+o0BhCnsbr2p+yx0CjWs4ecCu/EL8FGSBCYZjEGvNTshuxuOxRuvxbfqfme1IJp/Hevjegr
d0vFRzqtDLygPmzlGC6MdWgnwvcN1EY8aovMdtR0M++cEUUq2nPxqOeszO+WC33PLT25jAC2Fpqt
cCYahviKERWzdm3/zMJFAVvIvuY31JTK4Q7rnv0Gh+XZ4AwzndO0CYE0dkkawqkxXNFiQ2rOpOBB
1rFH8sF0PRSk4csG+bJS4H/J9z0pngQbBcVaJ+HhTW2vGx2U0WQ//Asfp4wsBwDaUBAMvgRF4dXN
FLp2S/oY4I1suTK0PdqMusQc41JcAmYjgcu/I2gw1mPh8xxpprOQDLPAU9rkLVnWrtAa2ROnkn8h
TI6j5gWG2wa01FgP7vtm1rhbIpP1VpxT9/+gKghlvGx82OCV7Asp1J+JsdFs9JnguP8g4oSrRW4r
9NR83DHTCVVk4IDjw5f2u1HAXzClQnmBTt6QcZHUae3r5TC68hXXzSR1LqI6td/3dr9Lw81pZ3xH
xh1KyoaEcRDkq5dedb4MppMBG8UjZvZxfeBoN4qKEZOsKvEWCOZdhLxu34/B5jrk3uJ+EZwHA5Kn
sL7+Sm09PqvYj9M1kwjTwGiBFglYqPc6BrhC+IirwH49UpwdmhdKvYtTMSSs5eXnkrPqNTC+CyPr
OfxMGIPyz87SCY19XGmxPYD+hc3t2J812HAf/panhHR9TEA+9tA5sfkC4cZAErsfFagRx5KfKG4z
qmi8hHqNWB5yudvZJDDsaC7N+v5CwmQ/LhtBAGq5XBQ3EG0oI24+tx9/khRhBXxAJFRh7PAOrCKo
BO1G29/+WalhG2NnP/BuM+e0/JXic6s9K56689roP7jicDV2jZhh85IM11L+sQl6eEjQ1WIMOKFn
tDKuP33u26hcSpwy08Yij0l/XY9t9YmRap/96lU6SbyN63KAmhYCLzEjg0ePd9yRFHKA2bkl2rIL
g+hkfWAiFueW/WGo+wC158ob3ZzsaUyslspacIV/4ejGDW38RmWIc9xXuAwFHU1VmuuLptihsYRF
Uj473z0GavU2wiutga7z6At3owV39/1U9xRLwdHfS2jnitdlOTIP7/tR7dbv922xbCpyK6+lYl+X
DSMbQBGd+IBWfD6Re06KwlV6jyCwrQWmp3ddF0JtxKONHKDa6xYnb9TdpqDxG2zdse8WZITgtKpV
yrx0tLRnRor4pPgj/9y3hEYmCuQKLaOlbcpOIPsH2KdG4Gg18BP2lSkoDPt0FA1+zYN9TuUUayqS
Va3cDBvHAj/Mn3rSX5bb/5PigBG43isl1x0GDGewnOEuQ03K9StSXzPbHPOUR70yNlsEzxKa7F4r
1FP40bv9nQNYrmqc8q0ZPUAT+jhlRX8cH1azVXxS2KV9ADdlE2yzuPQxTw2nvI3PhRMLaoeynzkO
687wZ1n07FndnHV7mThfzuq4vynji2LtOo4vgnmn2TYLSeEMmhKAZX79niJY7R38bNiXHjLt+4BE
vns4+Q1H/LGe1TKgosU3bs8ZGsSOXiIoXpVNAfW3l3EuUHA+b8j0fh8cpNoXPbBhYQBHgcykCmJe
QJwhvUqObnuSy5fX7D5z50Z9PKhGMzKrjr6q9swM8XruLiJz1YfUvHvXhAWDKs++mOebwhugx2X3
iekUVzxsYWSQDOwaC0MGbh7aWM+4Y+1ftYELW8eauwE2fumq9q7n3U1ZpZrwt45Rk/1fe/CPSF4G
X7E8QQmudqOWEjXjRn8W4ayCO5q716CvhGhMU21G8d2thI9TLwEsGqyPk2d23eWFshXIcF+gBwtS
KuJfmxT3VOzpbKz/Ykw7sLNDp90kRYqmLgzBnpAOB6Yv/pcRGAqjA7f5Kgh9WaYEIegPxTdgf6/j
A6nlEIrZTpj8BggKhQqOtrwFkTgPhuRZn5eb0rnP0R8h4wdBROs5KkzejfWJFIYovZ/iYV336Ah1
tdSHg3bQCKuGyxJqD3U+TmfeFn0I2GPla/OmiHHSVxIfxybROvRpDUugJpP+dtAn2K8KdPXRsF99
BHKg9gNZ/DhC3ZcVeNLQnKpP9YFywvJkdJSDywWjJAxZcKDnQGv4tVorQ6JU6eEoJt3k7w+8M8RD
SD2noLzO2q9KnU/Tohb9bH4mVQwAAChg3I5Tw8Plpyl93JjEAM6kDYsZjr3DGN1c63ZFk75e/CE4
mqGIkH1ayFB6JBOeGrcECt2R4jZKE6OieqwRjeEczZn0Yzfrs8jIJyDVurocATGmX8nU7PsQAC/P
jINs9CZn3aMemykhcCVQJQZuUmcJS2e3YBmK1hBmudKKI3z/PKgCEm91VyNZMhfBfCGYwcGPhpWx
4WiJku8CrsI/9vRBSoXRzY8T42x6xiPIO87EXpMsls8TFCAM//x3/i/QSUM/miH7d7q4J9+wMmG0
2yC4k8pO/D94/341Smt2ZehV3V/s0MPdg7r1g3367PVmEP4FGyQwARretDI3oWPh4GYVXxTWq6dR
knNQT3lLgZaAXka6pjLoZaUSm8Sx+WfuSeAk68FmmlGAoCRJRtFqohk+ELytW9L1GA5Nig+7I00Q
sLp+t826QAYwcnKu0F2XhD6yR6z5+vz34E5OOFcD7wz7VrNR74ojqUUkIhE3iGoQcpyyj3bMQ7YW
7P09OcUHnGULBFWi6Oy5T7MWm0iI4T0gywxcPWRDjk2uNkBL5K+zSYYo99+3ndSzJmxUKvNEHJ5H
pypOsEY2OKqNTNucEns2ghcoZufHE7BhA1i7KxNGjLwYHFDxrzozUXOSI2ntmFA75kk9jmF91sPo
RGtAVQPWU9olM5GG+5UXVf4YSLFmp2rsZ3ee4Mk+6BWbSXitsUMQZBBa85UAXD7gPwsWRkxQUJx7
Q5LUhYrnnpkRSSdV18pfVvmEbtEyozDHUcJRsVv0mMzHt2Be75F3gGoxhHqtEk7L9sUVktQhb7Ag
CTUaIiC82Za+oCWQjTQxNmV1HJUQ974IC7NXJlFHISbdAwhOTTSEJOyz9gkzxRzs5Fk+DUBc7xmE
DNIU+CWTK4XoOFIcAgMD1SUR8MNHHjCX3nIInXkBZVohzFGHkE2SoD21VVj+Htxyw9fsoqxYeiAx
46WhaebHJ/bE3E6SeQk6gWB9IUR+eZkkGd3/6D+61BHttxsUfjdLCwmkk75Q/HR0UJkJkXc3yG72
CCBjr7NnoqPXk5EgVQBixVJogkLMowQRy8SKUbwamyOrH0Oh9gqNORIF7vforeFBeQ5+ZImD2dum
EqCnJeaPrnSuej4spy9QTtbyJWBBQ5CErYV6f3E5ZLVlxtJAu6Jlm6OKiPWCBwiUn7XLxm/TGTFC
HsFqGWVFH1tahn8+tnXeTtRbjNKLJiEeNo3EvqxQsv9P6e2QZBJogOv+l37fUGUxQ8lXc8FGI66O
Dfc/hyQGS0spBlbfIZDQzakxiiaWw94s9caspOg+U02VO6narHOlI5Mz3KicVvdaSf0fyrHR7jxL
efAW6kl68tsqzzrNPVXYzUj0tnfKZpB+TUMtxjbq6HZtgnmW6zDyxQ370J5Mnnyw4wPzddcyZHxF
l98kZLoW88FnOmqWQ5/D7oAEEcA5BpyoTy0Q0uhlP58zKR/a2bi3Q4tJPr2Qf+CZbW/fkv9NgUmF
Ip9tWI9FoP76WllJgu9t9xPYotLNMDr1Ez2rTt0J+UhLwRNsA489XNVHcew74mc1bGq5xtRdORx+
vbVINJi+G2KDKckm6KmFDs7HpZwMdpSYhQd19ZNf5Hj/sKn++BlPhw/tPNpMenbY30h/o60MoqBV
fMNftBtj7me0+mUuWbZj+2x8Yp48jhvTG3WmrinVcPFH0MpU94iFr7eCuX47wRH/PNXcK0VNeJ04
Hr/qi2rHb2kto+MQLnXITjkdV5a00IaklEz38lzbjAQKI8+dEzFiBU4C4OOLaCsvlzxayAttD01I
diXnp0DdHXe+CbJmKLhfSUEAN8FInuvNK7Hvhv2Oo+XemnKRNUomdz5xKhcac1cK5TMOpokoOplb
jtb8ybij9Or2sN3G8imWzglp1vIKD7jTLpMFqqwwiHyEIBhoZaXOpFP8FnfJLcaxrOTx5QhBt7t4
6z3q9jnVGaFIR2B5RxBLUNFPRJNJQhKQdhpaL6xFAiyjPhwDrftl4hu3HfJ90saSyJVhGZxOuDjX
bnw/aSs0yb4dTHVb1ykEkvSGDG4doVMGCI8FyhfQqTDVc7ADGxT1vuBxJGKCXW+oo7gDcYJxS0Jf
susKd+WFK+titiHO7JY5jjf4z3ywreRPgahUoKOcAFHjheXMMbUXSDJEP96w3cf053vSTZDQN1oW
ZSKDbNrtsgAfpV4L1Y7mxVBu/8b0+IYUvfIbBUiqDh+nvekSxfaGPe8hbej8tdjzFL28TYJkAaxs
3zYy4hLawrVvrKdk6M955fatctYDTc0r6HztQLCx6qgCj68ei98r4ViKhoyX7FejatsXOpWWY2tm
RtsERwWUUkmBYQXpSynBpYT/dYkMHf2yk56TsBP8WvjtAUlpt1LqT6QFNqRUNroT//83hrYLtBGy
7en3cTujWJ0qezh5jgqoBU7rLOYLgg1o5nsTGkRcmzDGkA+5ayFpyxdjr3cEZaJfyoHw4MiV8Azv
1cR8qm1g+By+YqdkhvvKbUmAKSr5OJew43il6s6Qa+3Ijxq52YZHxR/QRsW0Hh4RyUxQWUiVavjH
3/m1UrXpUMjkKuRy/CZtY25bxP/Y1g/7g2FZbaBwGZQB/4HYFtLJlj/p7G7XXMx7/T4xFK4OvFPS
0GJYRBgqiZwmtZZ/rQ3v517U1B/yo1qcNrdAKj7HlwJ0KF534/kKpjMcW+1v8198Io8w9ZGjqZ8I
6bCt+TwmN4teTbnaitWEmqpGLP33PdkOsc1WnL3rntffbD3KTr3+WRBMTs1ERsyOH2SnTD5jFUcv
q5JLTYGOnImssQC7rLbSO5s236y0FlFubhG1VPe7eG3LM4pnWiY5ys1p20fpOkcxWIJD0aBdTdcB
r6Mw5Nh0zGeUhqu0Mm/zKtg9bjo5BKxMsBPs8BqfXFVKNeVpShDiwhyNtf/LuAZfkiBgYt5/UEm3
Qd2P3MseTh0DtxBNH0DC5zwNAyEt2YWEt4HCw9Wepub9KXjN651HQxlfRgwof1cphTa1ExeKkqUn
0Hw9Szz2jBW9vIfG5kdq8srzWfWu2S2lytEnyw/YkrRO4ZCHL5w74+OnR8XWkh5zvV8hws8Q+U1u
4GnY1UJa4Qzmabdi/zF7S9YYxioB8iYPHnvHFHhk4kw60uB/J3fDxkI3xMocAXIbjMSVNR+oH028
yBEDXrCxQfKjEMhSjlOT7l70/pSXjLBHo6BbN/3908z2zWu5ehWh6BEvqq62Pmeyz9Rr3mbDhSKB
QE+/8cycDAovDHtZOg+6ux3tATI5cgDmrsTG4c4Ji/H6V3d5m0pPyA9zNp+xQFZcMUr42gzC/VVb
e95uBFq62v4SgAYLHKeNfpjUiGUqFIn6Vj74VnGoX8Ki2YFCjrNfLmwyoY18S0Kc/yWd2X9T4u5T
/s3l/dUdto4eJhzR6rQfkYdJjDcn78ezgp684m2TodMRI+tx7lXatg4u0LhVLsFT6CAhHOeJKluS
V08KNj1y1Sp7uBNrOLAgJ2+W7tRy4JvdxaOnFc7B9bJAN0dCiTP2lv7G1DysFoMYJejmzn4aS6e/
tftGPHLml9BuLxuB0TA5bHT+QgpZg/6LAJogiVpYZf8RrBA5HKmnjfsnI5iF+9FXrW/4g4J0y2Y0
xqWnY3B6AxDdeSV3dVn0NsIdC/+HIZpVImwNMLRyr3pI4GbAm0CCTfg+7+qVE5rG91RYWy4or/Tr
PICGJpXSVgSA3FBw4HQSo98BeOcSFFzo5Sv5DxlBN39EUaUU2R89EUAXaGDYM1eiXM8dyPOqYkwZ
61oozZDubViRb/Osc6QwDK5qW0zlLf53ZEFozBSSrNBysDOVhXHkgpI+cPOqLHRXbf/G7YAFViae
oQUdJCcrSjMhW+0wCTqUguZDDEYGU7DdCLExZM5tDbklmpa6zRkda51Wad2qYx0bz66d75xOQaLn
karXJ5uq31sXIwphlil6WHaOe/1MLDCOUHws+nGsgP4mrlJhkACFBaqhnR8amCsAUE1brU/+St0L
EM0oQ/J8i1BTq3keU6u4ZKTYmRYUe0E/w2xrwvwXYh7T5HEtQY0+Q+SJ6EX6R5dRQ2IqmeJohOKP
hE7BeZyll+x9Xa27zQ+/2fW6ML/Fi6h7HODC49a+Pm3pXELji5f8d2wL2ylwcZEy3qZmJ0SpwxFx
9LEqFIUmwLHX7j4bLUOK5pnGv3V1qwxsXipzeh7BQbaU6EJUdSJKqWReqFa0RGgoeHflqfL+dQf1
Ys4o0CWrsqE8n681tFWPYo2dhLRZmesU3Mw0VQmo5a+cysPrVfmgt2l3TOBFCuWLszGzSOU9VTRm
RwFpqGy9j/ighP64epirwZ9PKtbzPCgUwoUWgAnWvE9MpBrNxPxGPmngipcaQBbU0Yp+Ik1vCFOm
NxWZAuWarX521x4vuQsxX4MhV5FZyluR2U3Qu/01zldWqVkmM7MIsJAvcR2wMKQxqsIZSbNhSvDg
X6Slc8r6ie9wZkheAhAXsEgzN8U6HL1eUXR+tEKDcHo8UzceWmTtvpN2ba8hJEfDAh2Gn18aV+2D
opVIwpGOwWVMn2wyf0glXwGsWe+Rd03Qmd44op8NTMYcxNXXUt6BRIO5xxzqhzhthJK2i7t7fHaM
ETPGsXZqzqhPMYPAzKqcdbDFdeitu67iMKOBWWFmbCvWPd4I6gLTh9r8HGIWKgnyS6rTNBKd05Lh
qwEN0eJIsQDG6yHxN1y+AfgzVmAxkxNmJNbI7Dl0DgpIsKiPuNkpYdhaExHD40aHC77ryBQqj9rs
T9p0OHjNdeyZdj1N9bkn39vMrGShQtHe8QMXMwC3MIZSvGvj94xyyNyprkMw0yqPAsX9kmYXUc5T
vSgr9uthvr66km82e4F7hmJSyDCKsiXaoA70mDY58cibmsBLMfCwEQIYUW3gI9kYq7/pO+vkWxI6
CZfLf44vCit/Q9rbQQV0Vi7/mLCbfzTlO0DYrJXXsTmZ6SF3RSg8SAOc8j3LOz9QuGSDLJlqDF6/
8zBuURx8b3WWwFnOgUvC0AOMchLRoA4kQha9ERqPqZy8OGoJebUvR8+lSK6bQnlVfo6eBK/q03KO
UTaOaARGamRG29fkUgkbAoWw7KVs6JuChiBxR7EDo3SKaCUU61lZNOJh7KehXoUAnQe6gYv4QDUc
EwxrIc1Qru8YR7KyG8p0VGSUoQ1CHK7oF9eeSjybRQbWTLVoA2FaZ3DRx46N5WIkglZpnuN45b4O
/nkrwzUKf9Aj2wuVEKN8dnif+YmdnPUpsnydmNvpoqGsfPI+I4b17+Nv2VtrzaC7tgPYoWh4jfGC
T12iX5IrV+2yKl2Dxe7GaGfANthCsEvMcBbkx5FyWwTMjpAFeSlGxzUv8ksEphtow4HRjRlGDW/L
SYdDPfyFsDN6sDRK+nJkRU8L9JAo1xoKE3hI0s8lxBiRrqTcynbBJohvflgLET6SUWXTGHeBemxn
riNTFRxRmF1i2Bxt0+qh7zdvtM6AB/shFioPfRAq/n/Y75HY6BiIL5+3Ika/IRyYPwQEgBYv/2q5
YeZCvoU15RJXYG7V7Kp/dZ4OG8WjxqSHS6tx7J73QBCQeHpFTGJk8iXjTbpLa6cidxmylrZTUwWD
VUt3Eu5yrBAN3E7s8GRTQrnX+zbPtvVklkTts9FG0F9Ef4bito2b9sqJ70UPZCtW5EJgNLkyPC4t
HWewpvgJV3JTrvqfxKw0JMyeaMISKtqv1bCXOx8p88xgGLgbYjhoc2CsOzcFrjsRmLPEhOMejzyX
q+CqvWfqQ92KeZDqEBg+d1lVDd9XZpVhIAwNCd0niGgfbAqa8x9bEbKwKQGZWFYCbMVV2yw02dwN
UK9Ka/frmmBIc0VKyqy0pOURhI3h6H2cGQM7JPfI8HdS6iZulgqhlMFUJhW6vfpyxenXpBs+TER4
48mkF0uYAM4TekWGhRFymqjyjVUnzuT/PEpRdba8xsf3KQiPL+lbuBLJ8q9Yry4ulUE+jysk6PVU
w8Qx11avqRZ/TVAR7QgjuETkjmzQjhcg4Txogag2AmxmgnuS2dcQufFq5ByIEotg5hageGyzLxX3
P3Efexhv79nQGmBHdg7FAE6gMsPMCy/xqgdSea39cFh0tzWrS36L3kbMLHKxhDseypQMHAiKDf2+
IJWOllMk79GGIZJYGNiib5xXtwTL12TAClArYE+UX0TvLoNnfcAhNyFkHaiNndLWLCC0wx6K6EzF
+HrZOnL3YGGCs3T1B52T/pa+pbAOwz5NcCVqGD+IewN0X5U+ZHw/a49qEuQ6CWxqK21MuMP4r6f6
HrB5wDK83KGm3Bb1l42BNr6otjWzBOeTZxB8DKrlnfDIiHMDSgO7e4e+Yh6F+4njSpo0ZYFL6R49
PyXT8NcdIpLmrtyN4CLiAXfA/iXR7gPqg6DQ1vYs9Ldoyat0VntRDDSlC74C1kPiYtFuMtkjuIij
IhO3i+FIT9Ky+BMhSWNLGdM3CTDjHIkfA79t0rsdb7VdIOA0fdvxUnxfGPkhvzW8qVECh0Q9nI2C
Vf3JLZZqgfip9EuzP9YpMYhvdCydBjBG2ZT00jXjcjRGR9vshAUOFSXMesJXn8U9ZdXKmYEA8csQ
/EdqkWNEcks7q0ElcIDNZi8Mprv+eRXdrDLwrPfgMKMdvozeCQdLkoNjZaDCUXm/oGLD8EUSXQk0
rm0U2OnV+gnr6NFDFyTKxXN4DwtjhwdueK1EEucZTYE3IOYc+D+mDVd92tpj4d2zVkVo9IFK2uEq
kSdUchQsaGvsCq6rK1U/PuEijHAay4wA+Bh/bRDNosHGKe6sfYzUd/G9cjrSztc7Snktwm8QbEBB
r6XUsOq70hqWYAGhqas2lerhKvKrwvjLPrOU7tKSOuUau4nv56AkQogn2yWOXgojcT9hxsLnEYIY
x3CqVYOydJ3ZS92LWELdiv8Wd2viFVQfD3V9L7JQ25iYctVXoYuoN5PL21cSq8fLfO3+d5Ya5MkN
evNzXqu2Pd0xHTzFNM6ZCimj7ffymd+Z6kUDRdPWk2YyBH2kRuITyAMvo4xSibX9y/pVwf4q6ngU
6kkFx3hduubJI/lZLDyvm94s0zNGOwFfmGijHDxk99CR/YxIFQmeto/sTvanrIrta/2U3xfI6EUc
X9ngMnXb6sInpJ+LhrTKSQasewYurPUpuI2AjRE8NnEbuv0aw6iz/CJbgvU/VTdHo6UE0T5I9ORG
zElXf1kb3J5/KR2nzhlg0w7TpqQiTtsRZ+EV2wJZWf4YmSMq2OZ7rMOAQ/MWwLL2vkhoToA+1u46
aEGjycLYKvaFK/7vWuTbgtjem8oTBU3EoO7w48EOV4kZ2qY25sys3VvyYNWkT1SE6NJHc/UlDmcB
s5JZmW6NHYtKB1/D9YynoPlO/xuqj1OH3pfAgWV3FI20EoF+eMP5sNhdMJ7hmdtOcbcJYjPKprMt
ryzTMEykvtaqRlaig1XHWS5OvyUx3WcHXti9yocTl4PdZCbbDsjObZ3rlsck/EZ8jr0LvUmEQHkU
VgnrWNE7qI6VX5t9Yehe78opy6Lob+z8F1RCVPHP+wvrVJ0N86C2NyuxyVAEhKLFmokKfE3hGBj4
V6OIGw5pDY2sm+0hb7s+PG2UF8OiPDM5D+2RZKXEXo3WH34mNg7NbZW6adU3Mc04cOqxx7UUDkpN
ARs6C4Cb5sr1WXrleZ2FFcrrk8h3FFrNFd8zqMYNNlUmx4JI+koPtS8K9EFaZOYqCI0MnM7CjxmC
MBnpmeoadhvQsQkcLtxY6cqJchOwzF1MDUeYHVr+CkTXMPU7UiDf6GIhEDTNkgScF/kRuk3C6D1Y
ZRB5Ol7/1SMAsN4wtDgctIz/HnRxk9GB+WJfsXF5sWn/e8OeWcIyz6GdgeY9i4o/MVpw/qpD3oR1
jprP3hqg4Q1FU+Z4D42hcA67fh8tU7O4FkzBMaA7sArx7RxkkkE2btvbHEdytjnzPtFi1AiN2N4a
pre+Ymt8753zBZ+F9ECFeBIGDR1f7kthTdUH9Z39eCo4EU6SzAEyMiu4KVlkBSCx1pn++0M9kPaX
dlnzbc2jvTi2LQNaok0AqUEZGsp/I8ZczTkDJfGs9tLURCvnQJM7yCcIFI9V2SqL/OyFaIlgrVZd
Mluv0T8/hjjneOmSkNrnfZANNwbMFXvWos6k9HZQM+j6pOqd5LNjR/Qt8g20tAsydSvIoQIBjQfU
rr80JGmAccHUqbGASAMytgKTKA+RnyWcxfE0FsCWUVw/myVbgEWbrH44xU1BbUTTX1KyUiOkfyJA
icxXpnnfv5RjMH+uIEOjm6KM8d1acjSBT8+adhHF3KyW+2dzTT2sLinaExKuQVa77Z2upqjDSJ7y
Q4suLq7C1A9d/IH+Dr3C7dsGnFKf23np73oEeH6CbXmiwDKs3uF250R/ai2APoA0Btylgm5mHcCK
Ag5R+8kfU+A5p5RmCkyhIfHH+IwVVeoe9UgwUUXOnudjru4xPlD76rBuwsEmJNglG5TxF6sALfzB
/NUJZ2ClNbePMoNrxCeIxP2XYbbNDsZGn0hR4eInM0+4EoG0r7hymUq62UTmCHZpu+M94HSP8K6A
dCRLCNoWEiYkA53Em7vhQ6/7KNrwluJEEjmAf/bME6IXWy4zxrBLTkcbx101KuEjLKerto64GpMW
d7LWHPD+02KaTk92qYrBHFEnqCf/popB1pWxa/bDbypjJ+IR2iUXiX9/OV6AXnGuQVTjTbwqomhg
N1CZeQe0q2CdC9KA47VqtXAFsOHNhIvUMmvmhntDJIXelheggekiwXQnG3rEwuPYEAqsGfuncjnn
82mLv3YLTbHbiRHT64beCCoT6Dt5djSGgC0SRGo6vw5hVlY1j3I4PRddo3Dxq5rzCtUpiXVAMBy8
O7GsxjQnjV561bo/mgVYphBbrmYbCuNhRhdzvUXGxsZ1aT6wXoh/205jXNqfJa71Z5hKvegAk7EM
tz4AQUPNdiJTobzHhtVg1eyhtx91Rh7D0OV1guwE1AMuR0SqBfgZlNlWcxeD66uJ8ft9RA5jyd4H
C5F7fbPDA6nUNkOyhBiPQjLB4AeSQtClAFGr3p8Bz35Onjzj4su70KuDEPUzMYs6ZhbLFNVlgLn3
AFPNQLup1IeuN6znawi2429tGa6/fPcqXQqRcscZ5eGu7cKrhgro6UPMQXwH76AlVjL52CbTUMLN
zNCh8jTcUhEwBU9VfmSqgmabadcPH3rIYUVVVhpIt0c2LvVCgrT1KRLoosZ+CCmPGrzyif7xFF0o
p371vEdyxVpw45ww6siYaG90pFCBj1XksXXyh3JVz7WiYNwz8B268Vmt8RJ+OC0+m1VQAPjU4R5S
QdlGOAnQmnuQRQ7EKSbOqIBlKaoZyCrVaurP1g0vOS40GNBIs/Jqa/R0ZVY4bxenG1zGLskvzsok
a6Le3O+99XBLza1jOR66ItrMHqBSwvhxi5xqWHTF+T3q4G9I81ckCeaULnswVZXuFpySi7GIZyRH
MZ+0xuj7B+0/sTbUy0j/zrXIveFGH6KHLrbSjKb2xMLCSZN0QzGuEQBm545V/yt0GuXIQqGCF2Wx
PeP+1rstbuuj+4ftvuSm61XNc3bxMYtCDsVetqeyp0n42WhRviiTmDykJWWeFzXwEdNi/Y5i4HGn
i2TEF6DesdQ1IUz23zfRXSveCo9p6+yLD3ZkjG1VS0eNyXTI5PZ8ixtY68kPyX7tCtnm7LOqmIow
qmjBSfK6OWN9NNFX/8ZL+sdgg3QKOU+m2U1XbBsu1u4wOpJL47dAXOVLIJ0uoVe55HXqnxlm++wF
fvGHcoeryLtEpcflbWzk7oHue11QTtvvkCWhCuQX6t6K8zBTBvtZDxCjcnLpf3uVULmRvQ4m26Xf
Dda9Mo3WI7X1hyyiNs2KJG5Fm2PySjdw4zxRvA0nQNKGWDebIYhnFugk+bC9Rszjc+qb8vdTGE2g
tiKywIlk8LAEM8pmbMddfBupJrWLlZtoZtFvR+OcAPN5MNPU5bBbq2IkX55dGQs5+3/vPKnfL3xN
ATkDio0ETxAHrfHHEkBEpFw9/z3jCRUgRXRsn9h5K9RWBOKcTQp7M8RATIBJVLeqwWyvNLKwSf5T
X9XsTywvp1xwqGcCVpCX8e+mIlIj434A97EvSEjPBh7omyFRoD6ftgRTmCDyYpSbiFvV4M+VuEj8
z9qj+rJsAm+U9O814QqSSycJM2nYjeRDux7b1IifkzcYU3Y75ypx3qbkNoZOJIPmXFkhVSdGsVax
nZ+aJRkBpcCf2IWAcUf9KbaIa4X2IOSkycnu/qBpN3XYUYxK5bhDNeyQDDPWYuzZntmDgbs2zDGV
THFca5UhrHhJfoqeND5k0z5/fFAGWPgT/l6pLHdeMVlT/1ZfzINlRMx73Wwe1MerbIgZ26hAscaU
E6j/t7urRBcg4/MP0iiEwzYdzWaA/lZ7DQmB2Xz103zCB29RFDoq68YTmRTo/HKWx7t2Mk4BWUh5
EmnCWBYXToTMiwu6sc/2oufnmIj5ojjH5m9j3lfjZdUSxjL/cjIvOAPpoFA79yqM1FcT0AzUmNlI
E8lLyl9k7dUEre1vCNTysZlHLunvN9A4ywtniPKeR4dePqC5Zic9Iv3sNHAMkhCBxLtiZXNXNiBs
ClvgZrM5gin15XaWbaYvKyoOYDZ+55dipfIu0SlDx9wG0RnWideRcgIfcHH4HqsMRXWVRsix52xI
8NDV05jN+d+TiRBtILZAo6qJ29MKCwyRuRNehjv6XFNjlOMHr1JIIzKDKlHBYoUBa3nFOSYpBUwu
ddWaXQOIIBu9DOjCybJcwkMBwSp+Jd957uM6o5icQf+t79yciGFt9UJoOtpyi++YSNnyDLi1VZRD
t0NmdY2NBxtpBj4jUVYREeLy+iIfqMXXAA4JUNVsEGQ1kNVQXTNP8TfOmOT/28eUujIgaIx6+B8a
auWBfVm8VG7bJ9dv7ibX29mTNc+xTg0Mnrv+v5kqXGqDwJD6T3/agLRF40/CIYBZnx0mof1rZh7i
5Gbwe2Q1gTMWJ3lgjrgqXVpp6HhTe4dXDazsYoBlgR63w8/A2d99kru1CxvYHzF64723pesfYg3M
kL/td9jMZ9ZWx61p9i2hAR4Qeu/D7G6AmNdUFEwakoldFQuvdnBg2SL0NgOzGlPrOU/fIWprLO+V
Kg6HF981Kd5RrtWFxmTtciULuISCDU7hAdANd6rA3PhkBNtgU/y4GK5hJcC2B6LAFJRao3Zke7vn
8EWQphkJdzK9DcBZlmwZCd+DdHVfIaEC1CGhO8e6x/hYmFfwlyghws5ueBbH8tNuXmxLDr4rUmmo
6QVtyEx1MNYAJKq2pQImQ6w4BxTmhKteaM0x2U9FQCfG0RnOjJd9XJSUbJZO8FEEGgZHCHOAlppW
pvAOaS9dqx1pGxE8j+xRrYsDKglQXEVW9DFCNOZoJNCAn0QlatZUasMGRMiIw3tsrU63xdPgX1H5
MTNkQxcrKyYIo+rsWlPWCt7q2OZCQT77TeqGADA2kMhAD3bZBpygk+823cK1ATjqnODexHE1HjSs
Uz33wL916cllfMw7ildPz9lUu2ELEp/7Hd4Hl5vHMbCLKPIpfRswQiAhAJ5fjPAottWYFflQo5q1
hzjebxWYqBUMUrDiZOl385XilePAajZAkLo3W7c92mS/5swDogoYZN8pZ1svC4eCnv9b1Tg6zJ74
w568Z7wNQMVuX+LbmcAYZXm+E2fwc0pVIflz+Q3FAR6xN0pnI1oZ+o5Qefb2CJdyADiLPvTuFmhn
edG/c/xS8PKLe/yvzPmA7w8L9YOeH3ltVSFH3nlLnlw+T/kjA/dybDL+PP2vq9KKwVNQjWIORjae
jMtcClyKIaZUhXw7sBCO0nLsU0u/QwfPwxlKccMQRWzw1GTrsyFkwZ0FII3zETbaHPlIfSUVjV0z
8L1fjHhYYe/ijU9mcDmT7lAeD3QnkZ6vZAlL3oDwcAEP69he6TVjsd1l0EZViUpcH0dvA2WCxXsQ
Rc61jlOUGRB9dq1QQ659kRU0OcgqujHtBEpqmrPpz21vuXUNIpxpXvIaRRdlk3AA8i0UVuDhrWmC
jZRDtad8/jGzIBOrm2bf7g1rtoeU+7sjKwvLX5rW8VDU+lbB8UNJrVxggQypPovTY5mKPwCbVbrY
a3f7kLgA6PTLqsRg5csZ8e/JQ3BHzluaBI7JZ6QWm693H+oydNCr8pFHaGoXSowwBJY9HfzTs8De
6lH5vh+r43cFON1N9cRYP/vVopH5R9B/eXKEbh9hwg2hGFLHKUaBabPAzYqlX0my+OTFvuPm9hRY
zfqMg10WRVkuQIPg1TcdVvCFOomlEAgEsaAk7+mDOcmj3Bzj25tTXfhyTTzBHQV7Goy+ZETx8+fv
boXu9j6CRSK0Ta39DY8R6ICeQFrTfMUo2dKqWue6UgmqASt2zNgHR6q5nnIm63fweoJKAcwk26oA
R6cdPLlLuP2TlCfTzUpJOH96H9byB8PQiCENemlb2NKfwBgL6KRKMOOpmHJosNdDuEYmEv8kCRk+
ObzV3vw89HPzkvYUD93vqhjVHRlCkjoKv1QU6MGHq2M8FmUNQt/Uxdstw2vr5RIvP0OZO+5R66sR
3S2BTzjrNiG5oJaoOY/UuL237oj+tGcvw8kKtLsJiJQPITEXZW9qZgSs7wd3qQcdc5xcQpCzjeXa
UoU6DgYl+SOi2XhnJK5NeF7EnMOqric66IH9+pxdiLpt+lyKQvFavZYQaqeIfAuROYdNn/MhlnlA
c0e6LnUSb97WMEhk1VKZE5Pm4BxWdwcyY+J3sYvNlBmtqSFsLSRjmFoSBAptjK668bKa0FB/rVUv
6OkYcQOo5a5YoQok2+nMqaGbQnj3RAenWBy27sv60j3J2vrYwBXSCkORerd5dQ41dg9Zewn0TIpN
oWP0urZLdfMwY4pIXYKDZXTfmFefiYFwior347SOi+6q8tYcWjlhhVTs+hJQhrN8fLhDBKKr2fM0
UjXoN/kgRu5JqPNOz6lj4IYJ0IPsxLgnO/YkZ9rOAiuu8h+2bK7vsQdKwZxjmSf03cAsdPQYpIfD
cfAdtnmmbaElNrRFEydcDGL6sZesb5BaIm1xsIigO3kbLxe4Jv0TbdY5CenDVup5r5Vk8tPt7bEW
U3UtB+IrJrE0NHAiLotZE4WXP2vP63cgsGAzRr7Vcuot9jtRDXKLvazNlT8nrLlrkSvVBxWkIhe/
Qm9BMcoT+JPZD7WwUi9ZYn/WBFosyN5tJ5K+esiOT9cMdMi5CB0xiXIDTHPqNptiBm4ff0HbdoSa
JxLrosG9f9oGO4qrU0ejOOTcn4vDRTEOxLvyUNeNqfudxTebK2Oh+KedW3La8iZ6JPaRIpegtATB
HqZjQvMRoD4LWhEK8WpIFNjXhASHu8okuFc+yAFlnLJkF6+sodv6FBf9HWhSF2Qc2uL72NjXP8ww
KuiYfpeqG0P/fkzfyxAqNrvAneerYHj9Qc0TEcjVPEHZzDjzQrn5WQrxtJ68zSTyrQPCPeTjeB2J
YXfrWGSLPeVHCgH4dDK1/HOCNoJx7Y8vryHBYnuMb3KIX4GAbGphL0xFzSJOGKw6AIwxaGQ/mspf
L3IVZLfnbR0aNJbdgarOceWmcKU+aerpO306qfGrPCmwDaw1H8nLMz+7ZzY/XklVOuU3zSrVUYZO
nlzAJ4JZS+v0JgBSDu+jQHKF4RlJmuMCMnG357tUulqL+RrmjPDymW8ZsKbGGD5Pggpb5UjNfb+i
HSYjXTvJQvge5MdUoMDyA+3QC+a7XxR83GIGabfGMpbOcoyUJwVD0RtTnbysmS8bbGu9IS6OWRqb
gaVPBkgvPNnN9ELSoAiRixAfcZnLQ9t/bfI+tc3FIgqVzgeBTGICUK7AKDzuNaW2foqde2k5hUS9
vIS5k8LLePDfrxscZjbOnyiYTQSlwEaZLwJuoFBvjgzk10HoA2OvGrg7TTQrJUGfBT5t0mHjRDbZ
UJFo6X+An7AsqoJT8aXGiYevrnUDxpteDbZ87l2kDGFjHPGifi6d/pkFAz9ayQRxvXUyxv19r3qH
m25hh3Y+DfFEmgyzUDbZBLCNo4KAJ7ghX39RjlrbYGugHy0hBpTaKkRlaA+V5e4NrXXw/Ey7eKdN
4AQ4Lnp3kr8ULyYE1ZV/GA050TUhLra1rEtJmwt9QUaMTqe/WEMcRqV1LV1PhTY5dG0jDwCQG3PW
bobgfuuajVrMqJD6DfmgIswtqw3tJl7tExmlZxSD6iDfjsSNaqjrd4GTz9mxQmHWRzwtozak1kz+
jqFVwkI3V4Smko5ZqT50CiIDWPS0UZ5cr+sdY1AFpJqAUM9HpragJoXp/pDlyKLBJrp3mxGpw5WQ
/+pDnW7PSp/LYLtK6aF9A2jxy5A0FR5Ei+UPrWU73/6hcJkemIY4ix1CbjF6tYz+cOElgpFDDnij
ha06evw+dYVHTaA0zYXd1AJPn5V14B91V5ahCjSWn34htAOEMpTi4fiSukafJTmuBAAjf45BI7qn
yol/EOMqbvcjJ+fiy+K9eWI8UCSJYkLM6NAxTKU9OZTuftdFZAjevgAZY3MTI7tGl6KtB/MjBhur
e6o7xlji6YldDsf95CDcZE8aYJeeGWuHrSxvpWHV6AzBYVNC0DGFuzK6NcZsCiFmckV/yqcrzBzP
KPrLc3RpNEJr2iJvIjxw4Lg2X+5VAMOzn4VnHbqM93SRIwanbyF3bcN9fT7cFRn/pO7fP62FDnhP
jRqMbDQ2nEwDmT0lnfhka3qbwxqBXgJ70AdUYOvHRKzdyaSDMIA/XHaLYmGl9ugZJVGnjZzJ+XWB
dQ79/qKhAMvVbSI6xbZnqkC5XpDAjTK5PWlZ6xF/I5DjsjvkRboiHGKVraJAohT0j45HzuOS2xIf
M/51tWVyw4Z/WO1dXPCgFirAirwgplSZWXZalh6eGyBJMRB/DVB+oIXzF76LgyRve9X8f2GYC657
biQ8FXe1v4ibLyp87c+RW1DIpDSRnWrHibaoLRTxbZoe+ni1e2IObri2ztM5/eHFJt61o80PM0dR
DpV/ULcJnAO6cYWL6prdLWRdAPS56+I4fqkj/U9OiYEm+88HIeTBJwl01CFlcI74fuQO4d541LKk
oB14OFXkBmPommIAxvHdZVrchHiOU8ksZRSWD7Xc17FQe3jcL7sZ0ai/EM0sDKrEspAHwFygUGsi
urf3Eah2OAM58X29NMs5rY6bbSvscwirKohot187PUIMeMet7CZku760dXxQ5SfIHSa8qmnDAZoL
UG6ktTiKyzMcqKrE3ppEM2D/katjoSxvSzC9GSibN2+VfTPWgDirXlGg0ITsPfw8s1SIuOo5b1d5
QC1ULeFFoWAeol2W5XEdkKqy5mCbT8St3060A/pwm+JUdLZzKDnHcVsc5wH9l9m8tMs9HVgZiHSl
bjRn0i/1/dOap5bp92vHzC7AlTZKChyZMVC3Zi23fOZxhwjZKOrjApkGn83vd7+eUjT4KNjTPR3Z
R6ZD/43cD6iYdPRZpc/+ytsYD6YEbp6DPYZNGE705cLC7jCB35yShLLA0TmEcmzkGVD5C1ny2JUR
PTc4PTZT97QcuKfoBFLKGKh77u0R6soRAVDnUbhkqJj+Jfeh0Z15EdXnnxC4pvHbsqeBpYvdMfUT
WVHeG2eLuHDnYIhkGH1XDsnGqV9SLhxhffQ5UDjItnp0m2KG3RkJEq2fORJe6G2TXtyBDXqemMwE
iDG0TyvHinkNAIC6NxDIEVYmBRGRVm51RmwzEqRCwcIX+AnaOY24+LLhJvVBbBUKyz7l+CAXDTnG
iAT6ONXXYs4ehzcaBIR8CXmHmAEEVMHl4IlRbq/s8I/QtA92Wj6Sp6wNPZxZE+MX15HHekzY8ztK
0jTgMQnDjWDWjh6qm8sXMjd24nPBlN/RLrvHbxKoF5gVlIoId4+FAYoCqcFSbZHBJiW24AFF/+7e
qyOtGqDXc8OiTeEunX+45mIKHdQOiI8co2c7kDvfpPTCW7yFOHT2FLEzeWyPtYjZMot6JyzbOrZZ
uXxa9l157S+R/ybmHL+V1Q1oUSnmhh8JaqRTwHMF7AtSrDzhTgKwFEn3Qp14FqfqMPGWe8DQzinq
gvuIMnXQgWSsNbf4vNZFHUqURlcADQ9h8gQjvgfRWQYUCRew7RqrRI1W6XjltAwCHoLDR6TKuy+w
tfx7VPMyyuqjys/w1/ZCGyMDDT3k4H/qwDK1z4uqR6SePogmffuG4yDBu9f0xZrlAEeLcGz5TuuT
C+6v2DWu/2p9pP5gBSRht6X6cROlaMzbB7VuecYkvDoJ4M9HepvUH+w4V6fKTvsStB62PHJ5IP6I
XAqRA4LWAgylDe/N865k//FVJTI80ag1BbD3m1vYHGQq6ekV9sbvLtSRhzxV2eFkyL91YfOafzlq
RQVVYWkBuYWbUCLNSg9I8ze8LVGgdrZyCTTBixCGfjiOk6R6/hLhz/XOlLzeEl7BDn2KgtzA+2Gs
y+GUjgae9INcDvN+fmfLWQ6/+G4+tQQvJ3uuHyPPSpH1WbKK1qzZHmYql2g/WzkPYx2RFSrM8wd7
MD+jmm6XzZz8SR1Wco8Izv5prEMe6qcT2dNZ79PybUpJzn0OIO/C3d9SyllbJiNGHg7iCiGyRF/I
bJQeY1+8kjP47nEHPrDp3ElgSJu35dG8E1WxM8752uAdHtQqjQtwv0xfCC3SpStkCvcXKCt1Hv4V
ObMbV2zvF3eMT/mJXIMmJfRC6S4JxHP1/A4uI6WWoN2R8hI5nvkxcJWXw5W9fLIb2Kcj5oVSrSGs
BCvwT/Zz9GGZiUoNnfoynV5K5+eSeYAFKatipSkPXt8T8pZfHUjTc0CA9OSiD5daCSeB8iLL4+cS
2BbtQXqiwJUy/AZGlt7xRcJdYIpK5zf7YVyhx200VUnoYhOH9nKoqbVV8VHYHKf+LS45E4jwHuOt
KGy6s06PNccyl0AI+XuTv2HOxzv85cZtlzjTkU2ZoRD1o/MVUJBBOAWdc2x12HuSd5dGPQnesGOf
lGa1/RDVxi8rXcRc0UElvbvHTpGBUfrqUjn+Pyecu1mMUBafdHGTyCGLewEcoWFSNSxvlJ6ie/qw
nCoNl10QVh6yK4MltaH7dAVwuqzg1n4SDjwhucfem123Y0ZaAqUQWy+eaooUNv0OoEpSRXrrqIF2
RV4stUNN3uEddl0Zbbffyyrg55f7S+mMFtqzNzDg59oT1V9rDW4CevcPY6z0KKFxzs3Tajf1RN9u
EQUZzalPDcKy/qDXyF5b+nw6StUx/jPC1IJY78TL/WPJRzvhlTdQAjNzGtrt5wLLULjgekHHaQnx
nQIhZ+334L7E/ajKgg8ZjC5WRlth8nt9BHpszwfYMN9EmeMRoC4anRyssvci5EH7DJZCBiInBfcT
DW+5kPOEUeAQEUeZHtUwmGLZV5/RqsMjdWrS9mglbS7S2fwaMp9pWQSpJ/v3F2M2TL9zump8Ytt1
FrJmbksXp/73oU7orDItaAasMG1M/S2fqA+pYcBYETTKa6TbQBaQQQjj3vltB/cUmHD+EOrczJ10
JRevbYpKyWqSgonZooaxcfIrdpcyP9OHn3LPeJW4ovlQzVh+TTMteWD4NEDonAoK0ZzyH3ZyUPi9
MQFVkTGw5ZizsXsqO6whwlFy2zxqxkOlWJV8/cj+bZKyv43/Skz7+TMsQLUdRYoCQsVQub1Xu/S3
8eiqo2Pw9YDRjMowY6VC6NdzNa2Seeh7iiFfEAgLV9r0AeaZlyf8motNnE1rXmRaiffMm1kVo2P8
/TZeuoAt8hE9UtJSwNNCwRshbZn1dy7aCoqslXC+H7ZbZEbFyH3e3Jy+nOczGRz8gFWDWM0f2oWX
KdNUIDi6MZfU2yZ26/V1LrYbJymscAHBqh4aAfZRmVni6XCubXnsCgZ4zkmX9V/EZVKl366xTsKG
X0vIcvSPvHrfO8pUsaXMx7r2jklxvbAIW6HEjRZ4Yck0utWImIpQDaTrGs2CK+ZKk+ZkP2svYdr9
ZZCD5/IuQYctYA82rabiKm9TbR4zc8tU0EB7Z9onJiuAJWXsgqmw//qfyYWSYAF/wjxKLbF2aFvW
opSBG3ynxc637+UdQAcc+sRfJI1kQtxVHyOp4rpfgY+7cWcXdQqh52JbsCPXmPPpobKYKMVeYDCb
j/LYMFR1EuQOEuZPJUvDZ992D5K8TclyzXbKZhBjrZke356Bjv4jfuSKa2ZbNFV70HoQ7nJDlXR3
QzMfmLlWSl/mQg48temGN6vViZNISE2uH7Jpi+DiEmV1T1VhOwazr9B30Ykof0mTnyqv/YU2tJSJ
VRlqsWV8JaFiunXnWcOco4WLcDrVi4EnHJNMtcMAPgUhDSPlZXLJfNEQ3IZ6ZhKyLsO7aNIeSuca
zHj0Xt3Dtf5dAYv5gFbde6ZvDU6v5EnLqKukngeHNh6j6D+i3oXSNoorzlWstaUqUM6ZrSWGrfe0
0wBpjiapl/nnYOHMo8qnwzK2vEJBCgv2Ru6AJxXP8QK2RviKOFb8KIB8CoWOyFsIpSH+RGDfXQZy
lmpT5/dRow/n5bE5GZald5UGBS1h1/ux5fMCNg/ultYEI6MqDR+lj+P1BW+ofGpSYbCpXyt/pT2D
d5M77dYsva9w7fI0fnq2byzIEtROAI5d0a+tRb+w7cxHqYx84/w/pUhmJb5BkMHeVKpLba/rBABv
T1E759SSjNexW7CqeFJRScrNwaIwtW6Wb2m2CE++A8ycnRlruOLzbqIo5WnUPmct/sz+FCPMYnpP
RPdwelz7NFSYduV7ci9CDaYtOPmNjJvPjx+oBCOMcV56Ic0xrxhBVPCpLNj4m8txeoS8l56NSMRa
LZCm+5qkmlODkcHwpu1RCCZIOstc45SSpNacnYVdhccYqNIapAAnb8q/lKd8JzGpDn9EvgkJU8DZ
4gmwZDmUCUTcv+RlNFfz4jGgnHlXuE81wxt1GbBQYjNeA2xk5FQwGcfIgueb7M45cNKVVPrjuiLy
1dNSXApBGGKJhA8Lf8llmhJImqDMgSRQfTnI64WedJKVfBTk9KzP7K7D/WpaT5dhWzKv1VFXs7YR
dHAP0gWwteDjPqkvz7WEC05oIokKxfU7nIU7Vy4NPQWasKeXQcNcky4veG6Q2Oe3pHTOVKnyp+Kv
/JwVza7t4H41ZPBdb+QU+7xRzCjbiZnYDmg3E4zLGI6j4t4JE9jb6gJ0jxlq1jveLq1CRrFuNhJZ
BE5tiX387s/mG6Pla9lVTnWvK4B5skizTxsXG7fS9iJJ0qy5Fjrcipjik1nhbOJKFUPmuLDR0GEj
peEyeWO0rUwWEV/n1OSMZ4SWJ7Sl5MSpxjM9fncYvTY4Yeb/cXWpKzuNp+R0HqICx1i7ElMdjRup
Vqm6BG7qzq/JKb977KTlDUrQEUWnNJMtADeqe3SKGcZRNA18Pk/oWDhBrnYC0MxY68IgF1fNm3Dn
1iShWWLlCLXTuqTaip/LUEiGeBbfEITccU2gUb/pdyBm4FsoFoCplX60N0Hk49ah3zsvne+Ih4W9
sQ7Mm5OK3nKfLkkF9vZjw2itrKnrAybAeInsI25dZQ7jVt0iDJgeNxVYOoYVPqmL6kdt82ZU0z6O
Bcc0yKcIINqukUfZ+jjxBPET3GRHv/2XqgkI9a+v7UdGhRgkVVINI52GwmP7DyCkDYE/I2SHs2Jw
ABYqMTmjul8fkCp4YkXo8VnqTw+yZHeDpt64xu0v8DMP2kz7G9aC7e9QVzmBtpuO8z0+XrutgOYT
wg2ReJB07z5bKkhBF0aGRb6rN07e5PQuqJxMzEZvqx42931bN0c6T+4C7SNSSxoIVJXvsdnlIhRU
+6EIkbDW7x1+vOirDJbx0kJnTuJrAdCE38VkSvKY/saCWogMD4pG+ugXhVayV9O9PKQEcM33k1CE
327NwIH3YpEAvfmGczWnjdGfGuVr2trAk0+nyhvZp2GNlTZdJYFd075kqrrLVX+0kAN9Lxa69s88
pBPkBI3QaYTYO+a4GLNgaLf+O7IjEBTOOxCv8Q5RP73iD3fPLXfeApjEouO+LmSAYN1J8ObZmQQc
jLjMNXZzChcO8Zr+avJpH1AimfNf0WwJJ1jdihXwirIxgP/4IKi6dYbHSYYCw+FW3QE7DIFGMx9l
n8wrJ13RUvWE2F+Md1SPVBKeAWMEXkjQSDbzgFcIHZSbU97MlcTLZlC5CQyWOPtnCbUPxTAxo094
hAMCqktFUEKLBlScva97F4zfRU/YRguKIdLBzCkCi2hWgHUA6mf+x8CBs/vNWdDvPoDJJzP9Up1m
KVGjAyEioIrtfQrWFLTtjx+EGNvYnYsG7GRv+jBP2lAZc0MhbCWSvXdqhFuDmI5k45zJmR7r5CFn
Gy9H9s+cAwjP7SLwgLmxNwYcKVOeTRP7QHGeoXM3HF1QNj7LNKjAVN53EGO/xJKJXlTRjYLWod5H
NId4q0+RYua5NeW5Go4z6+j1Ye2T/RyKD5zVParmdckFkCl9inwUFAo1MrLKcJwfoa3lQCGZJOev
G1YwiJCsAg2guioj9jYXk262WGbRsSyrbi+vy3Je84vGiVR5ny40NKyLUt4o6NS6ycCkxP4Knj1z
3+1D/rDR4E3SYhcXA9/028hPhIyy2XXZKlgswT0alVj7LcItgHl9U0a3WxRfHDBLGSrp3vWp/TqG
vytnNIqojhI8DKB1XWLWq3R46U7Am6SrSKD94El279/avofoApAWZkfGeyNZHKbS1d5f/YVIwrDL
UnNe6X2f8A4/hsUaxDqNtsYQoKLQS0bIG8Z96qtlketOT0LkShSCNANc8lcTYztOAAvpXH6XKIT+
Isa72FUdj+Sc66a3CRwS2bG57cUr1KQt0rgoTP4VlJ9hz6gNjD9ZIMoov19xnnDIuVbHDbbYra0l
Gn1wFqO5CZQPghS69ATwn22LXFhAwyReLdxyw8GnTP5UAEJx/tGSzKahDUGgtF16Xvi5TCRKv+Ui
nelCFJ+qPgr6/yOVuJxwPBrCqpCQpP09KpI0JZjI7Ep+KQUfdpZZ8eBKsjaOdI+qngP0QM+gNNvv
fK9rwD01GQYAfogk5GKFwZ9o+RrIGAmKwb0rePh4KflBUf/mwWJS5LsqIYQPjKeyVoGABIkGgGRZ
Q0eL3QsB4qTEmajMOLsr9xbjdFeM68ZQfs0q62JlRNFElW5BQIrZKxqFZBsrLRC8w+vJXPgamadM
ivLDx2LDKathcJ49GzIC33Q/XBpnJgJH5gt2t9K5+wt8zSUrIUkWBznTS5/VvyGYEO+IK2fsP8Qi
8QLXl9FsPL8x6uXpIkBypkweBqUtrzuAOLeZS9sjCO0rbaGzhdlBjfNvYih3YF6YpnFgwMHCoT/z
kmAPJGDZb7tbxmKwmlmO4MSG7A/NN5dCf2sKCF8GhGE3VlHRI1Wc4PoM4Vect57nKFVqWymhUgxg
HdqU2jU1t/KQ3Ju8UdZTxoQztK0J5ju9vA2XS0KbGvGI3Fso9bDQHYkHNKYCEaV+usn46q+mRhLJ
2ZVNIdNPaN82vJc85DFiGScaPKsQO8ELzULWVSA54/A2SxFnKnfJUW2LlFgwY6QoAErweAfI87e2
ASdGJlFhr4+swEOqibQeCS9J+38rCUocbLqKaC2EoFWRFhyGSJUuS765BtXztnlgWkVoDECLxIXu
LW1PwgyeYHmXi5ifUDr4hRfwHrOu77he0/SZnDD0RmexqVc+1ZaD6CX3lnd2pZ5G8YirptXlfoLR
iuuDqJ/7WyBLzAyRnezIByU9UBDmdcDBCE8cwoNowqg2HHlz02B2sTuZmMfo3xlyIZip72C6r02r
X3id/wTqeuP8vM9MoiRWTwW+E33myNPwru7Mcnti7eATEHpYezEsy2bvGsG5rcnuDltsjv+OQxWp
oE9KhgEHboxuGRvWUg1ZpyvfpCCJldoIC0I2TFx9wEQcsGWJQmujaBkF/FoAF+ek3DBVSgCF8gua
njwvt8GuGvUPj+ypd3O7X+DQpIEvi/wARi8a0M5G+DXGkhIMd6c+GI0JA8gE1zXb0Eny9oGmdkiF
d077m+P67zmq3QFHw3YVpgBKombsQ7KE4RLE8I8sa1Bh2xUyekNMSLgEkLqkhTX9p97XGXvSkRqQ
WrKloCPoEfO0F9ldW/GBBIYUQlxEfVq9IzdaoVt1M6W+KErfjrTwinrxKj9sVtTafgSw/liLkn3i
/sB1PnVmKrLibN+F1uL8lckm3gxRy80S3i91QR++oy8hQ9AAxxiduSChOVxf2PM1sNkwiY6H8FeM
zkUnYr3+qwuJUgkbo8JK5H9TnhfaXvA9XxZfS4ynt/pMWggp+tRT8w5SctnnYuh1D0rH6MW/caXL
v8E4MXzKj6LENhTYz4X5toiREcmZ2uylJJTyeAxMvNMuK4AOEUFpPYadgKMFGZDTfcKRQgss6Evc
+EHaWzReJi/beznME6YkmRHm/+vj90LrLPW5LdzRd+/hSBL2AVMBg6k7+aZQ9wt1rGJ1LhkM4rjW
ZdbgwVPy/ytKuaEuBm96TeWb8st+uwY2BBYTsjabn+or0uCDHBTZu/o4VA/u262aQXcZR7azsdie
wtrQCHGCMjXBIrtvcHJnhtTElH9El/QzcAYlLBiZbTX9fkf4azYjI08SB2za8vfo2GGcd5O5wVqK
4so0ba+9e74WzQTvv4p4KtBOVTiSUV6u09QI+C3G1Elpzogbnwigci/Q6478cL3Dmyyavv2Gr2b5
6OtQPa3N0OFOSHXzaTglQfSrzbaoXMuQpV9VdJ5SbyyyGlOTqvx+VpTe64BOG2B+HawcJe0Li+jQ
nZHwLb4nH0etppXmVJWy1MJ7Ut6Gplu8aCq+8ls55QeqQvJWHHZbDX3fe8ylMHVeVP52EUdK6b70
Mvzz1mQVfOrtzaBTsRqWYtClVVLH6J8gsr8uZrhX4d+Ws0D29M2YrSTeLHRnXviAzYC4blM+J+0Q
z9lQzhLZX7MIk3sBzeSHLbVaDeqBWdMAzbwLNMR2sbIFy8/53Y5VpkB1yCv1diIBbfrpoK1ILK54
f+vNNn6DluGbc3ROlKj9ILxT5ThoxT0ERnx2il93WzI0J6OaCSxTLSsuLZJcVojVFfVAXq53w9x6
tcjWcuQ1dtdy4o29qJbjq+Yz9LSitsl5JPqSZEaltRht/l/1tiCLVjvzISXstlTGkY/OxA65R8Kp
c3LHAFJR/SNM12k3Mp54XJ/V6xE+bYMHeYX6DgDT8nCh33cs047YBCIQEbIwbGZnr5bii4CjSiaJ
9RgnRhKXbgLfjKPBUIhn0x6QI9D+9201R5XmDtAF90vz0cSpMmxRif50O/51rOuW13Zb+V9kV0lN
BjcYpNX+gKoP2fPxwTb9aq1AoN13dFGgFf0RVdVp7bi7yKXXDLAHXBrHdg+Gpp5y84pHrjovAmgE
JsCdhfeWVjA0OO4f0mj59XHawjMzuDgLkvUt4szEt0Fi55Y53YTMW+CaLN35WgCqizE91HsIt3d/
/Bo+ASIHWRE/2lbbRXCUFUB+dqGH4vuZddCKE7xeaI3dW7+Hb6/xL6SG6JzCqXgAsqxnc+euN+9G
iKOchqsTb4/hi9x22nSgpqVlkXmOKPSTxxeQYkSvf6nz78ciu4+399+YiPC5cIWPopHLGUwf4Y8h
QERrP6D2mWGZQKwD/zyBs+4IyhZoYcHaKmyPxC77jXJKGpbtGghoDLJ8vmYbprJLZiVWU3cbgVCO
0LO892csNnaO2u6CDsyWJVhON0m+x7C89OTZEDECjqiDVOZyRD9Mo3VDzrs2OHczWjZtt+7OthN1
HHvgSn0WdyH7RxCgJdHGHLv9DTKREHGurEeDjByub+8Ci1hw1yYPoTbH1nqqu5uBk2sBL8E2nvUM
N9/pQi5gU2SXW8HBlcnBVEBkRqZQz5kVN4zGQhqeSUlxt7bkCc5Jyu2craZw7dnNid1OA+l/a6EM
+e1QO0IrWYydWBdq8gXcMfgy39JBcRKbNCH1NqHpGd+dCk8iIlbelvQqIbn4TCX8ONuRzNGaiFLX
75Zp7oVZwH5uNg3A7ujmnD7A0FCjgV7MIDU4K8nd7d2N3wT2iz2oJ+v2HttzfqLBcIl8fbektcWr
oIP04IU+q+uNDXIBtI5qmjSmkiiBzGutrzhh4PaYZl78gxZe4zNIt9BUHZDmDIUgzpJkncKQItqn
iYvBaOAsNWsN0vc2XDsZU/SL12z8RrNhCIbQ652aEl9g4V3HbRpHHpMpStcMh3KhnBgx4J7+X+os
X3/RFZy3FPoncvRHk6avWtpiVvQXyo2xaNc49boFqq4biKFw6l3z67TVW/PJEejSwvK+wr1EGXSb
T+f9HkIi8iM8y4rN5aDHL1yZY/qObEvfS3X5PHLCDRd37H5Yh8RnFF2wmRGw8YyHSQUBHxWfNSXq
pSJOwlnw2efVHPPHnpfjcLyotJqtMDdgLGP6XommxadT4evsEXLebHa57qUygoGML9n++KsGPqVE
tDjojh5FE6lRFTXCogiCxxBhKekqh9dlD5W7JS3VskQl+DId2Mx9S1MsKa5ygGEPFEPb1tGK24eB
SAhLr3RgQVTAOloyQDJWsQEoq1WrBUDGxG/IYj16dFQzNUOny14XrMtRnkSklV154p81oNZ138xG
OM6PRGWeoFnarHdNacjL+1BEPC0TjqfDRxGWnv3pvOs3z08RuHuVosqnD6XLAAEwv3p2DR/bRCVo
/5i46RLCbqvR7lnHcKoUDUttxxVQAVod70D8lxR1cwnkO7TwuT/mXh2QvSPJ3y3yAEeed8LUudQ2
zzs3nJNax7UbdkciO7CGsNsDmILX4j27Ph99zdfySQRDcFRvYRfrzN7i1h7SoL5kDb+Sd8tR/r9C
pWiJYc3BeMgzR/Nxhv3USrcknoiAmIB8cX25d8OFEOReKkRFfP48dZKi4yIvUI8jkPTS/pedqHLx
FY5+VL4ZkUwEmYwa9MtRrY9SV6+F1e/hxaByrJ9TM0uVAgrsWtCE1sVtiXbHngaeJFNbMwU2mgDO
cLszx59vaoEGbtT+5dseqxjHQxltx2z3eR/zOQMAVuek6G8/fARZ4pw45kG1yeE0hNfwIl7sRa72
ewECgiFpy/6ZGONJmp0T/Ys5fLv/GmHrm0O5TtewfJ7DKACmSxnyK4SqEwgeVD9YtIKCcfEGMCir
xoyPt7Sbg+D7Fsv7mdIYOxdvh0T1vbTmn5GmBAkT+BHBsHtX6GzHeiHbaHZY3Uu1ZqBsdqDVCV3u
bKcq4XqK+tn6PLUuaztwQ2Vqew7+ifkCuGwuuxqtUHkJx3Cdoey7kmM8b9TKwnG4Q8+07Br0Of4l
TpZ7AW5gd/qcjCy4LUUWrRStvHMgY74jHE7mhz8WTvzFSn/Tmt1Km176o3qYClYolUE/EAL2Sg9d
GC5B+lYGhjhE8grLlzjDpWQZ576PQFsnCOQyMU4gZC75k1Llp8CC5yWupjBq1HwnxMKGVKojqK0M
ip/GuYP9pWyxGZrbY1fRG+71vq0F3B/tXor/1rM66SGifePI3xLG/Gz+RvYH1HvBMRR8Xh+YdFRw
2V/7xFq36i22a1Yz+/rMpaU0pcdKxdfGPAA3KlGc3a3eeWuYqtWx164rxTSZs3RSEqMccnc8r7bG
rpbVuPO2a/BkLKDhqYs1WHyMem8O7pxR2sua+t0hipX6BjPs6kFFYd0+19pgq+ep7kdkI+DaUtfO
s51N+PA+X4D2JM9K52lcjERBNr/lo0D3BznEpHZSBQfpdEurbmNmi0oOyowdl6lxgku1bsl9FSin
wqaxNVLbd77QLTa2J2UDpRLl4rXTlIe+VSB6NYYJ9nIlQtXIZLhKvH6P4kMC/CfhQ6jcy1C0dSRm
H2rQsOJ1Oze2N2LJSgnUs4uR0EWmf/tY6017R8tkN2LrL/MpBHokYhT6Asxsyd4TQVbStb+9s9Yp
wHcjfgQSkic08zfVsYpZ/uCNCr34Fc7NU7q1151eBkww7s7h6nikz2Nc/0DWahKJMrm5rRLTcOGF
zGTZpILl0wC5NtUkqvhAaAPvJA8uCpZ9jnYFqpXsUzcBCUwpVRCEuxWc3IRNJ2LDwqcgVgNXEGXS
zSQeOE4v2xW/8FXo1f5JdcN+EASB/O+itdibRCveF9q4BHi+/Vyhw62eSwcIx2yFKrJ3wKzLzdZn
4iZSbsVrkBATXp1eeCCNur/izKRPcZ64/41CAHf+RsCTOIjYqLtGai/eY6NAQqEdaINaNHl0ti8o
z79AMzts7qhvWw0ZRzKKmimvx6o/WaO/gw7MLOvTagODGJVW5hqoWu/9kjDSrupFO/4Doy73LbZJ
J0MXFFpBDlsR44Hgy3+wi94aoSptR2ILkzTSMdkJ3m5bKp6FU2yLylrZ40MmswhqACKypou4MXzt
1bIzryjMwD8S4xgLmY+lAFI7UKg06jOlu3S56ciTfq4FVB2D4kza+XlXtV8wl/eNIiL2d5+d4N5y
n7XxoqCRixlhSc6pPSDLJORmt15YtmYqaHrXubdpFFU0ZkQtoEUT/8yJQYOz3O7dnGWadfnsBTCn
OXtoI/WTfs/5rXeXAZHBiIAIvar2qYzT1MBi91iWE/9uH1WRfpAjmlQhJk+NiJauZOx3auuUMik+
tSdrSCkmu15j3LeW14u5IS0YYFV5SHsOkSYF7V+xsQWMbFUx22H9N+7ivMSn2pYWIZ6/sPeyU072
IKJ0e1ov62244wvuQNXCV2aE5rxVQ3qHL+JnE5/17dKrru/+m3zj99QGdIuF2A8q7iIahV9CHjNd
yU0s+e1E3dxyOm59obQ6AWgAqWnWPX+y6E+asdg31Ib1r39BjDez3pNDe7rBSU20GS82OmVqRWk3
lOwVALt3+xOxW+zxZ0NJPrbQBhJE9s8i6abqs7EvRP4N9GBQRfBAiMM/lEbRLnT/tmC0mypB4J3u
1RBOC9kCPNgaEbUtv98fd10tCtTq5OMi5rYe1VofvzikJzMr/5TIxKOJ3mmJDIVt9kholh4RKGrY
otz+PuiIo8k6mFkEEKuenP21W8/MB0skM9T2DviW+gRQPe5w6y751s+kQASLT25yuBdA7oj6Y3OX
vRvQKke6ZLe3yt6Fa97d0rSseKGptvt1m+iOAwbRrdtbubZCBRx7Od+35UJ7c/SgwQfGp6lQuI7Z
LVg/0kxsz6mFUn/L8pmkc58pzjXbqKLfxZ/TR3RFTAmwMtnydRpMvrucySdfcuqUmoeudzWE+T+b
3vly7CcwjKLdHueWOp2y+ZpU3WU+lXfmwxGPP+R2ac60VfZK18KDcbRH2yZKVuqcy94hEDT19ZDg
YV87I92by/PE4rXGzDonvQEwIaXD1XRc9xyb5HTFaYNBAtE90JPk2q5RswOWUggu8UnHmKCk4dwm
H1OFH/J33Z9wlleL3fe6KUrUiw4tpRAN/CcIe5SccMPv9Hx7qeCkwRIIK3qJZUKcEqtE8bOqjKXu
mBQCK7/iIs6nnE4UB/izw+qJ5XJeAmqttnruOg6F3sEiyRq04pwrhrtAVPw3bOjuSMQdmy6zgKtd
xkXftS+IbvB+ooSH1izb6ziZ3fZqnaCL6Q+mLkLCAgUaX4SGQ0+/8aEin3YkZJFFcECAy5Og2CZa
bX1VC/qqzsw/kUYlVXXS4rTZH5gqTsKBqp8lBTnUIHSf0R2S+l7Whg1HqdmfHqrKopOcfqpVCRwc
CecLj8h+U8Lcu8sVnFy1xudS3QlYmvHDe3GqCZMguEvQzk24Ulx4/tpsXjD3+J8D44CVIN9LaWMb
rJPX3plhyzwKjectEaVpEF60nD/qgORBPB53/XEYOb96jd0D58T5/2jKbi5YJ5rcz9xHSHmeXXXr
tUOJN3x+6QVNK0u+THtoI2dpBgouEm0NhNk6sm8uZpq5uGttcakUfB6mZ1EmuvIs/6r3H4zlMsSX
IKpQiSuIZNlAkjtviVVUjzjWK2jUSK1QKtBijdCgni7JvJKqQvJjqQCkS8dQPxWw3+CXwrgt3pcn
mxDfyA6y8CIjaR/hQKhcPeEMkW0f0skCenNRrBWwmr+h+tqEW/lZ0ql0tS93a16ZAnhGkhr1Zqo0
Lan10PKWheYv4aMpFd2Ck6b0mANg1yCsGWeEh/iQJ9sqmmTKO58X5lFtVsn1WwGx4M2Sr5S171XX
P74A41Nj8erTkv13FubOQA0s3dXtKbxACiol2tzB0Dt4dXYOndrG6t4WHqNtUqFd6fGpHo9qeVqd
MwOsFjrYdGhFvSeYziDvEkPVBbOonYsoZJKQ2H0fn8SfexOalmt4q1LXbV3tZu9bbT57BxlKYcys
RKtS5nmp4y4qdROR/X0TEw07U9USO1qRqQIvD6ojAMPMKjm8sG5942xLz7R9+Xe+M0iurRSG4Bcw
bcktlFYbxnzExnY4jD+KtEWu9kcz18GrAbRvXNzyhjlU6sdJPS0c5abRKxX49w0kri4mcj7UYLTP
INGKFeeTYVb3bOq2lSfRDTEe9qAzGHbLdpF71HFWBDELc6I3VvbwZ+rrHgOsiMIcIvbMRVQf2uuk
Y4mfi76TaDZj++8q1R0tXi0PgbVJWkiicH948mxeYxbt1610EgOThW05RfwIubnoAntQSA9QuTdN
0MJ9BX4PDyWyDhW6YXyc/sbHZUN2z4fS9OECqnM6b+Wsj+dgk4xRXH+DOKtcsq8CB4rZgOxArEnd
kRai8P+q9DBRyIbPNBbuzAcB1ZoJRTwymV/8EKpHjeA+n1VQ5Tq3kcucj0TtxMoKExfHLxrlyorj
ytVodngLwlk9vZHrL5TXB1O3EVMviJezDtbTyQydpjQ/Oxba39QJnsfU/ohNZEdKbq/bLmly1zSN
fjOXADkv7pGB6nLcJQDgVhr4J2fTqmp9aTwro1/WfjR75+b0lT526UBw0J+30TeNct7MaltOWNB7
RyJIbX1THvnWYnM+vCZiaTxUZtk7KdfEivyNDuIcmihKnhY1YHiMfeo2OW3R+JmULhDrK7hZr+i4
xs6CM/U8TIprUtW98CH6adRprd8fP910BYGIHfSHhbrmojyqWv08yH6Ilzjst6Obk7X5HoPSFO0X
ynfw0kpNtH/Muz1n6l9b9QTIrCjUEG0BsZi9zX0Bj2BSdSRZ0oCj2RvFWdwfj9MMKDYGF+ytfzxh
6SCIMtJvMETQ4RmYET5CXP59+mG0fz5A2RyinFJ9/HHOrRg6q4a5FWx9GWFDO0RYXfOtDatCFJJ/
JHlx8nDQfhib107uevOAesqSlkmOchc9MTjG6M/0EZrMz/qPJXC/2GkZK/xWEETwNvjtDFFaNBYe
v8f8kY08ZpemcZPY+YUp+QhphcMXckJDK0ac+atnt+LeeAj/g/GbmtGCpfs+ZrMkbg83HeZdmsYT
ZwMmq1WpSpgMF0B1Q7Fv2kra5spKs6Kayd/EjgOeNdAT7nRWRAKs7l1hQqesXxCDRNkUEwGUH2kq
9Fb8jBGNZG7WvgjVZR6grgmegTH5UlDjam+P07wTPIZs1vICdsq+vEk8AsoShHZoBz1LCHj1icjJ
ylCTonOg3+l51nmohyT008wSusyzyZHdtLGKk22NLT2lJiyYw+IqZ6zXi6D8v2aPbZW7k8UrPQLW
A8gte95w0gl2yWkA1wjWcupYU12sMJ5MQ44STGdxkjJNIuYhGlbIpV8sFp42wmA070XUU5HSgjmc
bzt9d0VNiQcv8sPo3KKu41TyG3w/I9uuG5m9UxUjIrmnl5syVdghQ1NimfL8ZeA5dFChkkO9O1bs
zTrr8VV5MV0/Tlpo9JHEscb/EaZ4Mfc93dIaapcHAWZk2lMulloqIaZeOEbCNgZrz1J4KXwBVT1p
bBEmPNDrqVhSzJ+RrSdQprZjpDMIq4eF203OACpovzuUlDJbhQWtn8KJaxRbxoeUS7RJ94LzWJkB
zp3lYaC97y/Rwb6flxax83NS7R+KkTRzVb9rhIuYjXC5kKVWZJaiuWFBH4BPwiOKX8TTKWy8Ad4V
rdeMV1FtCYHTg4gVey0YKXu6lHG8SLmoAwreiLXh2xj6aGUuMspINLDoYM9NdQOGsquTh94LruHe
RRFVJj8sHCuO1KZhGXP+lLcjHNlifWSpotSY53mdTpMFvO0aL7muNzKsGDsr/OeFWrQI+bhBgt2Z
1gErdKBZdlKqG/4K2rG+vPB65/CfSvuRyky3OlvnnFMDFp3t5erimUOTTlLK06+1IPrRmt8ZENKN
nTuSh/hHS0hPEOEwdctBdDx/GWQqzpjoJiStGhG0PnP5ERMabt5NFrQ8xSe6zUQ0ELH4U0Keh9Zb
HZFiQgUgBqFf8WnDRKWro4bNUUN7KEf2v7kZ6zy25uAZvb9FS5NppbYqPksxi8fp1Lkz0jLHkFz2
Bg4fEGQH3YWMCXac8JO1pE6xVjvrWCNEHUK5C1XStSoHjpmNhQn7Zt7K3Hf9AOvNnLLglmWBHgzH
IfqeMRNzLBEkCmVExkATfT6ZDyd7UeDdfIvEqGMlYPhBqvFTKUvSWhMkfTTAbpHZ/7vI07r5W/m3
yXsE5/6sdYHpHCkyGfSpGQOBfRzXLYKz9HsdTYK5mlGctB8/iQ7xwtbTSeZxramcIMWJeM8OIgJS
edAkInKErgHOtZ14/Q9aYTv3t90ae6MHpNPB9BcFdsdl+pHg87EAWXSob9mZ8MVFG6qinUwHpqIa
UHJnWNvy6ztVNczJK+8rPkW3cxkl6YtnhtYnhFJFzw3lLbKIGx+CHdEKu2t+Z8K5BaqpxKgfQE7L
qOlK03piH7LTUdp9EiZApHrtEzT/nh1idYgyYZ64NPY2hq+vdkVj54GNpnCoxFtv+VWK/Y9JXXS0
Y24cFEXLfvcB6KHentMwzGi+DgwmsZbxyxCfmh46yCPxnosYFzZX0Hy1Sdl/M5t/PccnnfRZQjDK
aaRuAX6R60SQWUWBfBFN3NDiNwVyG+mErapogmXa143A5rbY7u4RmMNXqyA44CWSF7G79ToNPrO/
I67mFCnqzzyaz+zXrx/caVGmHJ+m2GntWhyNYXrs/bB30w5jA9B3+9IpOBF3hVT6hs0FuUx/l7tV
qGzaHdFq77d4Ifi1P5/jQzXzDWmaqLwS977ClgDhUcnzx2LIcWeJABiFWHs2F655BGZ0JSaH3/Y+
bplI3tOYEhC3729Sx1nK67c2in+3fl4YjE3kzfBwFcp28l2ysin7a9ZaISKM1nYU0UmQAvp0lCrc
H0rWEVALAPJQVAdrJOtN/19j5PCj58CzE4QL07fdDlyYWHc91XCNe+oe0x7aG747CiKQYNR2yrpp
ln2sH69A3M7vQzijv/GyBU57YPud5/rmEgsNgs2nxxcekgkpfzLABoiwntCPDWD7IHSAvxG9pE4v
uHcCU6vqNWuVkYAzXLwJOBO5zHrx26ZzppAcpy8nl4GJGmE1z7XipONefI15dvduQ79TrGB0dW5b
4f/GwoYYHFkmOdMW3aLlBpfG5RyzD0JE/hIgCOsROsjugkt9gUltF+Bn2swboEbmNDgbhXvj9VKa
2FO+C9EGoMVEUHaWZwOD9IwYEGRyZYQu52j9begU82P1/lQkOJ6EgRL3SWUwDwmOqMlDIqLK0izE
YS1dlV68FFLuEW0XTkSnwPLMe9IZj5sVKPMt34sPNtEmkbc1WzdXYs4Kx98NA8gBtXRPrt0S8Tzv
S0W1qRxCfSOFMEeAqhF2D2ow5YhtdK3P1nNmpyQuaeA942noFwpEG3E2kAeB/1DXYPWd6y5YU3En
RaE0sHRo/noQRg6P3DBce7OsOzwOpN7uOIv492bXDYF9N2FOk4y/rxz16f6aJTOcW5WOZMjNE223
j1qKxXXdZHOlC2ka7ma+M0i+ddoJ5KY0YD32ULH7AqihqdVKZj9LsI+7paPTXT577r9eGDfXfzc9
e1Y20v3SHbaVq/9+1UBUtqS1GgS43dNiNK0NykvS9Y0JfhBNPszqyVAVSRCauc6EUAFNe+E6BpgL
fSBkwUazjhY4h9nTu/1RfJkbZ9Qxgjz3IXSQLBGGo/Gtmi4HmkuUzdjPmBPkO2c/VPIuQpZ9IrtA
MzO2jSMlLLaJAvKGhnmc7/yEfJasODMvt+NyOo2lqr2C0/MGjg326y0P4DKd7+6Ig4sRaZSmTzqy
qqWV/WwbRhPs+/TUxDIaISJcK8SkdzGqMLHhnVhawNR0WqTe3FbXGrgFpjFitfDSzHhUoJs1pH2Z
ISPucThIo3ZBkh2mOLAAptKG3Z2eLtYLDlsyZc4WRf+r+ABnANZLQCZ8yRNZXzA0yvETMLFjt1eG
MHBEpqIMSNFbw/ghAV1V1jMGMcP2YsWifXarzTJS6mLVaSJY/L0F6BEYImnYpzrPxsX6lRNuEIhF
96a/LiIuG7vFIhPJP7PKA7NpgExo1KIiUP/URqTyfI0rP+Jv8sdGhG0P+24dx18JrbsvpFoZ8ZML
89xM3LHLK3Cg2qi7pgoVik3GIRqSEuLOdVvOaaPqZEYJTLzcHHMab9dITICLqHraAH6mr+qa3HdE
pqLQyTHjQ7dDeYPuXroM0lv+181CtUGdws6O7/jrLv+W8AnLKVtZZsIgead36Flm0snDwUWsf1yz
LqdxlkMOkAWIr7r435tqPw5D0eH3GJd0ng7kvMTUKHTWfm+qS6Sj6j81jIAnl6sFqJe1tFJa0/ny
fQD161mTRs+rsUFK022KjKRZjfm7/IIVp9it43Nczz0vzWb3LgB1UQ+23+puW4WG602XyWcNUdx+
UmnFnj9riJFKYpbfhcCzXB7KNAY50f8LKYTuw1X0Mf3QZNXUrjynqp3IVh3GNqn6LjuADzTMogqA
YlyGQzk+3IZXXSb7bnTGC/C+O4vj0BLrTzDk4fmzPZh93NN2HMbuf1/1KIir7paPowX7gk0mNDKq
CTb1dIepwLD3bhx4arkHtHDRmrRBrmxu+2wwso6ez+hYOqwTm2jUTNkPTR+ka8HFwdoRolQmF+oR
OAXIlN1bIHrfncPMTmtNcngnMEKyZ+4hGLkscqKYt2GMvvO62G/nhYEg53cDLeOsjhHlxjLyI4Tn
lwbcEERKzzBtb/+KjhuYHHbiXa5eW2lDdvIP4NuYaq4kMHb0fA22dt7ROTtGRCRTEEyC2fLEAxtJ
6PWq8pF/T3TXYa+U167k1qK5Z2TKm7lNHP/JikBLYxLTa+gBqtyehuwkwsr6kMnV69Wgo1BsDGnT
j5i07DUc0e5b7oKTq6tYPBiK7qJb6oY3FfjtkCci3UIKWprWX+H4WF+Svfr3n3U+ZLjQeq3BDy9e
kODQePZnHzNv3+bXJaq4KKLpDSxHdBg8DPc/24wtDKm5iVjv2L32SS99/UgmrWXFZ9WDFDbr3eGR
+qU7j/fqOkrecYFtC76NrK6lbijaa0SVP/kUK6Oh30hfWHBxXG3avyhNyeS2Vk1+6brLFlt8MmCt
cG8BpO0Y5xJdZBWadiaz34ObdEhxSqKM6S91pj2wL5qFzvEbiUWgF8854WP4wFUM81NQ7elkJk88
6pKjTT/mfAAZ09TpGCyjThyb/hhkjOFR2novll68eFwGqKhjHkDrqhgh6PpMuBU4YThKA53yQ9Hr
Me1XqSr0y8eGVDDwKreCcdte6ZEJJjgEBrf2ZjnglLsZ+9Ee8NAb24urUxyGEHwIQP6Kqk/AE3t7
Pf7HlfHe2w63QbDWIwWxi9JtsyxCActRt/YpfWQQRaq7ZOliy18aACnxfzIdaazSgopMA8GjxxvG
1VA/oBF2wFnnzpABtCeIP8kElnhvNpcpYaYI3fXt+KeDJWVdIRnhnZTUWSj0Fku4tmPx9UGeVH6P
v4ElE9z2m6NJkJG+NwZbRqkHgfYIDBao4oVzPObv+fYgX/2Oi3BUpH5h3LVLwrHq9yJUKRzxi7fW
tITTOivGrPw1WVBN6TSfMnfIxbuDwAjSgRCMAiqqpjYcl8tzTrVrUqqJZZsc4bsY5rMmRJcKhYrM
siyW7YUVtH856YtwJaFL1aPN1SQh5LNT4FdRcnGjpXc+c8RsKvlnWAk5MPzpQrAmsY1SRjNZVCOL
6fxoUsVPKqU45/4CxaYViOqu3wizlAIwukbUjxfbzlYfggOIjanW2ZOpTW4fborCe5wbpbdr0sgj
LTAKq47lY+RMIoZEeQInB8IqGGchVAzpoSqPUM9bwkjNNQ4RvjT9zVAoIUPTY49kFIaqkptuaSN1
J4AweyHoHcLNpWoP0+QHMq8mLBXPdRMiu8Ff50EaF1JWpadAgrmO+NCyWSBvineSo+gxpFlrUZMk
rlofvQkyHm5ToHy+nJjQHLh3/AbBQAgSHxPeNxITVLTfMx0hZdd4Bpg762D0Oh80r26jOqSqh3vm
YsPtHCAQzwtIrL5ElrxJt8vL88AegokEE7mwVtQad4qLvx+iT48HhG+tPqEFHCSomG6CvZouqhUy
AnJY4PXiR1LtxFG78GQ63qBMTAqwzClag3HJ5dwwb5JFZh4Ep+dh0gdvVfBbLgKPI30qr1cMdjHL
gPiHtdCOM62L0TguBvEE2pINu6CNdQBt4baASh4akP2sXPDR8wjJn1iXq0MJcpua0uU+ONoi/rI2
Kk8gKOq6baaW6inLwoGz4SW3nWHqeUwCEK4fAzbvKqPekv+c/bmSeKnP+33EF5k94wqfsMO/D4hz
xv7KH9JixHYSEYuCCpsjz+HpNCf9VQRhzIQcXzFNUawa+nHv4Khq23JrL2uXNAXbNJ0XPTx5OO+4
90Rjyn8PBQzkUI1vEksf2llqaHriRCw9TaBnFgpGOmcLyY/J/qZHLF8ssB7LcLDASsS+HehHzJrS
q56n5yGk6Jxvx+qfeSOrBTC6OtoHE61B6BD0GbrW3E03uon7ExGz38J6VRFe01kLhd1B1XfPlk8I
2k6dCHMp6QhgKhcrAcWD2goetd4IDrraBjlzEjTw+12ZRXBFXqxC0TsPMe4r5lA8nxVs+STCTn/1
AoVnm/yTYTU1yqAyW7o7f1mHMIjukf2f6P99684ZsIgEM4XyCGSQJkU+T7LdW75hnYP3F9YQWuD/
CqGr2odV6qEv27hLyk39IjFrVgdLjJBRg2hIo1FiV8hUUYc2C/lbKLczfuu3NM4GcsS+n42JKmG2
I0DMMV5Kj62SlptKHJVUnUT0+5EIWWtHMeonBz8wRUlZwJs3hgc7rOhCkGcGSzQtLO4lpRVqxEKm
JXQXB+u591mbBE2Fj1/Oz9JX29qi8gCvGbxKan9v6GkhWIY0jE030QURBtmVYO/rA09fxTUDud4u
eFxbBjbVJ8CcpOKkyouZcUYFXM9366ykU50m/TeteAWV2Y2xGCPygGCEMwLVzfJwtPrGF+GYJTsG
5/Cf3dYqoeJPNw8wKksdHvnGlwMt7NDcfR7Vt/oSO7hLwhRwIUhK/sH2WUgM0oNdwbvh1ztpX4Gs
X+OXVsWJ/3afjxwnqDACAPhuxE1rATlq35OmfvWmjTSzHCAjQM8F+aIWBrQcwpu+CCV2K+DoI5wn
RUrb6jygCzD3FaDGivBKI8s1Imzt8+m6rqK/qDQyITDRwhxofy1ZqKD1miX8YI+p6QgwJ+WfFt7V
y9gP5x2MMp1sbNL6lktEnAbGuqa+lY9r21CgBKouE6le7CKEdOVz2TLtRbV7CK7sVEf3LOlkPSXP
mQLAYvCoWuOn5D5qKz5RNawVrDWnHqdobCbOZJjqt/yxoAv0uF02At+qndVfPkH6Lk1ToGucWn6L
ODL/ujtydrKp19J2iOnfn5xmPCM8zLJ8KFUpStRGTMT1QgN+WlZXq4AVPWEN9xkKxWBkpwhUhBlo
rKfq6+kxu4S3SbVj6e4Mwlz67e1FvFEVHTKYG9RHjtUY8pWWOiULUw205SOa2GLw73sm5kEbJ9Ty
jDWRjepfawsaOX/t2pXRjo2RVwGQMba1XV98ShVDQVRLuGuf/igts2RSTSAZ8ra3nvx7R1cYbjmJ
K8B+SH1FLpdZxiV5wILJR8W9sZYazhiDQkLz7QSrNltqx0ZlaG4d4OPIFn9DkVoM6vX/8N8/esSG
t0mYkj8Zjo0D4gJn9ETi+Lf8whPtw+YV/NdnyfzR2A7qql1LMgVwgHs3Rq9JEJbzT24IWtIUtpyT
QoEcZGNSCBUsp+Lvsq9W6NI5AhnnOe8UNlACNfWoIld/0Z4U/xsnnFIUFKy4WdrkRVbjN97agTN7
VyNqIy2awkkKaBbTkl78Rom1LAcaxsScYCIQWDeX4lnmnBapv/qY+Fq16oC5IyvVjzyEqN4ZXzPY
gSa/WIVAiYUpZYTrB0ND0j+DUBUP9h9unh/96mrrsweWxTegZ+ZYbArH5EcWnqjUfeIDo2jYDjRg
NtpcGmpR5kF/TqMt+AqVUYK8MBiWbFSJLRMOGsG5BOFDBBmDIVwUVrV+oq6kxDRo5WAdRruRjDiA
Xf5ftDzA1aJNWfSiNTD6eAXYqiO446WjCa82GtIMcS4yk+icylWmvMMqY+8wbiT4vHbE/sOJrw07
XIXhFECRIvi5QvFsHFezhE4ou3Yj9BEzXttqvDUcy/xanjISexN9im4bdohM0ahOOBYUPhJu3hsA
l1W9Ulu6/3MNCC8YLYBvRLMkFXAIDnbXudE0dyDF9OuMqjvO4CkBpqS2kmOG6RdHKnbdgzfvNLwr
uLDSc8IOciWq1KXhnRyCaMNS78WS4n933vFl74Trd7SV+/DwFCb2cxUYgtKccWXHWiJKx6mrc9nX
40JUOvob/SFinY0/b/dFLYOCovX+k7qHHMTG/Dv4I8YFs8tNr9Vub3tR8fkvOF4WohJTy6iDzvpD
p74eX22J5jAXbgiey9HvKxtzcCNPSSy/dAR3D8uW8hgs0FcNCP+Pzw23dPXdY0JR06JuexX5oKBa
zbjitEOe4M9BUe7A2YK4O412Nxi5wfwFcOktfleA514wfLOY2oHscsMrUY6pCFz+Iqym0WLe433S
82MszLKqACpYJT6iBoVwHA2D9w/q+yExG7kDsLPb3z70W6ab5Agp6HmKwlztDpUF2aj1uFSOO8FD
rUFkVXm7aX9O6/nBEseV5T24p0cf6yg5s6+jlfNnuSlbwFxLXHfSP82oBgmIIvqdm1XO0WNcXQCc
V3xm7hujZj/z6XzhjSt4Tt9+dibyXThvxmlFEPnHc+fa8auZPfc1LccO6AqrgkvJZf6WTMkMiJ4W
p011cBB0kG5zc7oP7VrUyy6Ho1MSOAd5uWM22KmR//8TKlfW6xl+dsh9/eh5sZ38pyI5M3GuhVLH
1qDmsv8ySfj9B+m9Zmjcibq3XGpJGilBA3TgoSrUR7qUz4nKGOUCxIJLRtO31/AF4obC1aYghJBF
CoVU+iGPdSxsZ5ILsQNn01WkjqQ/gvX4i8dsl8R6DFHHllJi0l3exzMFBnXdyyE/Wn7/sbwP+SkE
7qDYDJpn0OPmqc/GjOrpFBLNcxvGczubsFs7q90IGEWk6tJ7KTTfiiuz7Kl+LV9SCOFfiB24h8tO
tDezeaeL5isbIFiJWX/fOvAJGeS1AjX2oiu+48rIhfeyAXdXGyTukPy60kLwC89g6mFbUM5zKhcY
RljpWlHHriFdGZk5kn86Tv+Z6TChIm8th74EWysvZfR/F3tSxLYrDP346OClqyTnw7b2drnQAMnV
mKunUaPlY/LZKMWH18QW0z9qZ+Cf5cp+JIiUSUP1SWjjSDJ3yQLAp+PuImwSW/oLxSM6ueoapaZN
U7BnGP5HRpDNroWctneGIGTUEZt5qcTCVyeQjqZSGW8YEUJ7qI4Y4EZmulg8MBuUP9+TK4kBjRqw
IlYpFBt6Xc7Mde60Mgv7WHWLj8Q3EWoxSqQfbBrMVb8ru+z+YnxczLN1GT9qawrl3nkDEhbmt3kz
3n3wIXuXszbRTwJwPFgGrHb2HFnplZI9RJyyZp7A6ipcgFF5HKgeNXCxC6Wndz7bquCX863vxV9h
XbB0dVEZeYK/1Z1J7vogOx1l0IlEAf3OtcQge896BvkRMQwQj2Q/cXgbgw7P7EfXC+Zd4COZJRLJ
49xCmoIovmMqwv4rku+S/qE8UtVUfY6Fu/kNuOAehFPHM/+2x1cOSt5tYiEGqGcYKRVweTRLRBXL
Qg9owIDXeu56nx+vUliXSH0/NsNund55R1j/gkD3vj6D0fAVpShNE6sh2w+eI2fUh23HO6yrSmZV
WrQEU7+KBBWuhcdPdVJIAoynwrHzP+z6CxKeDW8X/gKBdBvLzunqegyqhbfRJ55VGUoYAdaCiwOf
4N414i79pdT9Xk1Cefa8okLrubgLrMjWxVxb+169Oykhd68hALB9HCP/uOL0/wj5lg8HvR74N1N5
j/K54FqnVCnd6iODLA3cjXLTE58RKEautT9iCHdBxEqzAQvy/tMJ/8n1YqEuVZlJcF89fsEVJsXR
cXnoIf5MOFvQQVrA8yH3wn7MUbRxRh3cGd0/nA2SYlO7lQ4tISw8llFPxDMbEctwCS0ojskxT5pb
TfzAYNlf8JVB6WpcxbK2hSL2lkNALuxEobKBPPNCUn+jew7/U/s2lqPJWL/yc0YzhE3fjAXnIWp+
vVkPE0wAiEeqOMZbwDAS2pSjC6YugngA4t0A0i6PQ7U9Ahd283knsAcRPAjnDqGqI05DEeSwaJPM
zFIDdn7KQq5R489GIxzFHOal/mhnT042V0fzjp2VqYXjezQfHh0tFAWRQR4UKDPRdlNYi9Ck6fuY
0428uicAOHBToj3izIJdDODQPEHBvsYKSUA+gPTFD6qgtjemDFD+M0m35cwokwIfW04zW4pIYWK7
0ucqSGPMr/r7/rgmoi2R1Y7f2OB8bix2zEKwFabm1Kv4Vhwr7enATHSEd1OFlZPXQQcyPZ4jmOxH
ryyVdB+z8gSy0BOF/bPG+Of69LOp16ZThdXefiieCtvARioJhVPfWQnhUZB8gw/JSZaPCa7APFAp
p5sWGs2SoRjPRy9K1gxJDTPtR9BeKZ+niQ26u5mYpzU+kE43oYURM081xuEoQr8QAdLdHx6BGwvg
SitT19K6777p0QMsH+Xuxmmskp/CqB0iHBOlszzPPswArKUVLXVepcPjX12RPWX4ikLrdhWMpzBF
akzN5ditqJ7ocA6bSznunTP2oG+oPSqDYTr/B3FRuo151HvMNTbQAY2NBQf7ytSKn4BksDKdJeRT
F7amwx4/Rk6AakFebpY/4wDyy24734hyn1avRbBGK62h6KQ0xyRxeMun4dLe1jLzZ6zUOetjYDeC
ZQEm2z8sVFyTcGojcZcRrLksI7Nu6cHn7/CqhK/pijgT7iUUFCR4P6SDLVH7gzdYbgHjqLv34Qo3
KkH5Q1+RKjv2mU3IUBrKCCDH6tmELXXu9fUOKmrgPk3KpnLSkj4VU0Lv/0cV8J6Qr6ohpVjcGCtc
OohyJL2cmvdhSDLgWjLNH1PhDYnJ33bK9S/qfiAcmgQN15nUZ2TAiKwFSAuqxQDshSdu5+GaWmS4
uUIeJNvFrNA5wBYiNlZUuXkoOkStx5aiCLGN8HSP2VP9ko9R8HSqrjnPChEQyqutdk3UT1ZOrGqM
U98dqwGPtBnHalz5/C63tNepWrGSn08wDE5UEUpRKpc2Uy+WwQLIHSmP9d1mzpBxQmaDRoeSVy33
ToIPmKuRKi3wJOr3jGTAO38mM+XVGfNA4EXhMHpsAAxdq752/pIVL8yKiqyeqYahXkK7V49ikG95
pCPlK/f5Cl7vq+r3Lk5YTra7fBQ25zcWwaXOxHP4VxiWAWYY1oqUytycHxshzgpfYemormxjPZr0
amDNkPWa9QORNRnbOy4q2EimUEaEfg53v3CJJEgN9UkcRAmacEYtF8L2SbwdOg2U8fp+URut7fAJ
hWSiGlqCANfX0M+c/qsbq5IIc/R2CnZDAZw5hKaapyWM8Zk9vCxDGc0C/0tlZGC5tY94K0iU8kS0
wSFcDJrP1RLDl37Cy0urnAIbvq6e8KY+/ZVSDVAsQAkpLfF1BnxK1FNoNSusIuaePhUl8zGbCXw0
uj6Nqq8yAJRv2+FF3c/VkWCyPGA9qkP5ClhpETghotyxrp9KDYkp5gEB9I8kDrqXMWHkZE9yYt6o
fh2ExWnPfqW0fCUkHURuFB9tdi+8EysZ5G4/nLdsqgkzA5pu1W0kdWBvstBcIfZAAYI5BZbaUcWs
BJutIKeff87Gxq5W6Y422WIhLXpVBh27kYVjSTJYaO21X7kWgAAJgmBbWgfMU7Oqs2L8/kO7HD2c
NVBPV2D5fzObhFo2+9I4GPPDY+OOtYIuWUy/IzqrCP695mJdWWPFEja5LP4Y8FuZE6eb3S7CPmPN
4XXnFPIF2rxhfizJsR+tnudi0ipjs16Vzd7GG6CHwqnLaWVGhVT2r0CvwUIqGnMaC0WnBMqXH4hx
clfA22j97aJJYEpeBMlYG9yn1/ulyJvpFgcxFKbl29GkaGmnUGP5uIiAhCDXtWWr4k2wDpVUNkyQ
s96AYprDscn3b66L8YC2gZmN1JMoo+emQbiT8dQpRlZZQGllM5yL57kxt3lJks/f42aTqRZLgUPe
OeWfazAnziuG/4xNpbvkoq6dwQ4px/vfG32Lx95ZeNd5jrGbNHZTHpeohXDwPGP5lsYAV3SK2GxX
Ul8oYZHU8MsZBdADb5JfmVaVF4+wx/Mcb/ZwZM7alpXs4GdWTnXi6oTkNRjpvDeY2JNC1D/MPk6+
2a02qA5JFtbPuqNnJL/jRaoNfR6ZWerbUc8jIZCsFct/0nlP7g6+Lc0JkgsaNYZqf5SBMDUDekmB
ZROnU4KIqLGSGcx34Cyqwm8E11D7U7d+wT8OAEUzjWBHmLmYwDUbXLti2RTzDUvjWT0f7GaN/VyA
JJqRGVXyMvfbe0S+7R9E5AkVn6CcCLZnPDQFHGrSBWvD9ME8Lmwkl0Bg7iAcThnedO4q8bM49YDF
CpqHJqx46D4rocai4MrBKSjFZemPSlJ6Df8SHtZLuqA8SL7YgMU5F04CbjznvextRtO8iSnzWBkI
ORiZMJ/c+FrcT09nF4InyjdC51Lo+6MKzGSstyY/ZgaZ96fn8nuGaaLxUMxpBHIsSFL/rj/TFPGB
gYNj64wTZ5jb+bySA9n+HogYf6yU/QLStCR0QMpSfF+kM3qDZd7OksgJrsJ0PZxBwZ2nBdpEYeBH
kXVkGV29tgIIK932tUmKL09tvoLyiKiwSQiUDanadgTuqVDk4mABseiDYLPFiWlsU4+EQlMwaeob
sXDIpGRHCJi7TXPl03HAlskIys9V61kHD4M/09tdnQOQGKJdyaz4I6upX2ST0IfzwAUoMKGigLOn
XoCMFugDEibQHfl3DINELDRqr97WKj3MiNgHw+4zywIHbdougLMGpK55o25RBw7bgVyj306b+hqE
eHRfBdljGEZzJ9SbgzaolL+t5Ogb4j13naAu4Th5EiVh/7aRl1totIassMOowLWIdU92pp8GjPJc
rlZYI+v+jblQILywSFkTv6ceRsFsiQDM9TEIM3NBJ+wY53Rntl/EAzqUzGOUOpuT2EEGbM3plhCV
/d38cdQr4rAkrQejsJW6eqpY/CFouCOhkKVlkG6a9jqoIs/YBnAVo1M8gk39tDTfj14ohDHKccuO
YHmprUcDvw1lZ9ARmj0UbY7Mke0C2MF0D2VSfjb812w49ZZIf7tDH4wfg93i9LejfzEpjirn4xT+
tWPK2UeH9ZSfL6AONb3lzQh7y5aaso97gLwUTpvO/rz4ZLPkokIxqzVOWL6kvWFzasFIox+9q/iU
5Et5gydXSbMG6JVL3SGiSYSDaFVYgpynOjBEgWQi/m1/HfNy05vM/pn7U968rtXFR7xcJ4ABxyOE
5FP82/YJo9lP+BLAkqhQgHqSFuQI2Eg7qaY3wjkoPtEuLiDjk6cuKyzNJcQblZYb0+0Fd6OZ2dXm
6hC0OEPcbruWx94qLBbxhX/Sd3E88gOYq4DKvjG3DQ/sQ1lnQwMtDvihokW2wp0ALfPqBn9LPH0r
1ka6Oh3YgWKspMQraQbaIZUly+oe+q2tJmKZ6kg+RRngZljZncAGb0tyN4pTjA4WefXjhzC5biiW
n145nnhGtlygZE5JEDPX/mueMeRFNoQxktQfEnxVdXOTc3GnE3udFSqLiW6Qe2F0VcGLPmt7MZiA
1PvNNCODMOBxDAifTL99nQZTa3BXJPNBfnAZLR4NxdSQCfCWUEwWAwiIlsYWJDh3kInEqnPWAJ6m
aV5Isyhlh/iiNN0QojyOe0dThwaqRYfhDmqn7ftMv/gEmgLto7aBA0ZeVt01KzykuWH6FWSeHlWF
Zvpm5kkF9d73YFeYXefw2PI9kOa2Jn/swk0xFTtlu9hYavUfIrdvE0dtQPYUHDPMhu5Tjxbf9mBp
yXsi0wv8M3bIQUXlnaVXbHv/EU02gygrLbmi2ivrD0N19oTDXihGJswM/nzj5QPA4C/i/43i8EDm
Tx2s+TFJ1YebYWr2ev3lZcXW6WzyVl6SRctR+rbpGiZ7H5K3Et0qAiZUdw1ieUc7YtgiJ440ZzIg
7PzGQdbjeNOCubP05SRqKoD2C5FvGpRS8XtG9yIhcWlk17ZnseLH1hjx7RdCoKFbopMacNjtbadM
VHjqH1Pfrn6yOKDJgCpU3i0p5VjYPfLn2jOs8p/X/owKJHg6eaaQdKeClW669rhUvh0iP1qqaUPd
NppbO3p2WyWpctAMQ7NCwqAuCXDkQse7r+epd3VIx2pycvxa08k7YmXRc+c9r9OK5HLQnlnCGin9
REs1Hd9pYfblMlgQxtP4CkPTGrBrZHMjb6zmsFooYJtOxb/98iEf9XT5+BkxYjmDyUJbNTUU2mbc
rRaPsleDafK8NNR0NljHK42nB9mNAbSnk9aDa9TIgPeE71BVWsHixbYnpzDgKjF+Fed4YjjQ2DwB
MmazkNJL7EeHneS9ic+Qg+Nt0QkQKUVX9FlWgBLV/meMgJyv7xgzAj4rWSn2ExfNju3T6Hu6dqpD
hbPyRr0t7GfydkUQh6cEO9vkf81COv/XUl7yVbwQGS6Q4VyIUwchawqFYNsEDIiEaZilLJPEIKN/
Eto4FWG3pWJ9WtS1Y8kkSr151rHAt6vY/rZwDOHSF5Y8oDW3L6fV3NNeNp/HpOBc86FHOX1XTrd6
lIkaBmP8ETRNnyMmSiOQ7I+eYVFl2sWCX5g46aZdT/EG237AfWHLMLcwjsJ9JlO7MFB8bgP5gsXR
zViPFAgnBfyQm5Lbgv54LGzAVH3bbGv/R8O3XRNO9Bcoiak9Ifg3F8D+vBN3KwfyfxI9fgZEfgNl
xQ8xMQqajiO6vz0w7PM+EJv2DuGPrizubflfmGCX+c/MgmXhmWFD1hXKZNCNaP+vPK8MsuWhOWvV
Zz/JE7tbIm3HZQH5vRVwYQ3HNP4LpSe5dm4BeItSrfbEEfLi8KzKlnJkD9OD2FQCedsJKetcdUdp
zEVIbAdWYrUrN7xfutdjan7+yNmKz66hgR40ibzlAj5XMtyWE3m8xIZc7/coMXvKbbR9oOnALFJ1
u5z/StE3leeUtdhsryAnEfPV3iJrRglL+a6Fvs5IS5vL6awsCPbmpxaIptu9ANHcTelRnucWNAy5
PXR8zIl+dgwLNFIajFTC5COqGKbbF9CuDnDoUJbkh/yN5fpFCyOnW7rr4J7P071omE3I3zeYr8zx
u9F186STFRA90aEbn3vQ2vUgx+yUbmLvYOT/dFrINoZH5X6dmqMWmGHFWUaj7R1kJGhct0srh4S0
Ecf4ysYNIp+oGVrzsYTOjxRO3H2B8RbCdbkb9eINqzHuBM2NwEKCDbDvKYTax2xwRApm99day+H0
2uET6r3Gs96NI6EqzdAVNhdUk8upvApc0kITzLqAQDF7NCcFAp5j65tn8EQP4GR3tmI/M/SeiHCB
yT/9vaeAd6yqwAvxPsrTdN+IUDETJperOvCTe1CfU5Ib/fGNsyzBE2iWVH2B5U90tjNF88JLtFwF
OdXUlcaoNn3hexQVE+16Di3iUFPSE0oSVlJWslk6NUg6CNbhgfjXi20o+j787vKyA/XQg55pvodD
rjV40wm3xS7R30fukdQQJ64P2YOhJk0ddS22WAph5yWwapUhkDigR2z4mG75Slw5lytILm+7gGXQ
bhWGbjR4GH98hMqLcX9h3SAqjx21bTtqmsBc+wf3kBFSWgceVFuR/avnwXy/c+NC2rAOkswOVjlI
9PnmrMJ8H9S6wpigmkENJMR4RhPtU9mdUdYPEJFnf0G7zx4GVRZH4TiCCHY9+92qQALYoeu1HLxr
YrJrTqEKnffM1BaXzpa6ewmpn7OUlbWyKEv1A0bl9NCPJDl3lbmszRZdDdfQ+7jnLsF0gY548U/L
NFPdTqkc+VS96zOUqac15l3e2pb25PUsDbQ9VadxlZ2WW9GBgefyrJeDcnRS0HyUehcPj2TzLvHI
F1r/Vlms+DIHD3fuVtLTDUbjmi149hP5ibnESF40kb4U8FFZYSDK2paCf1pba4hH5MQ0/QcbiFR8
4r37OT149E+WxyPb68yoxu+9/soBdaqgvgCyAlg0c/zrGDqNXDvzm6N5JpFzb7hnxNx5lV6r3m3D
kt+wh803bHXJk96TzC6UV8mFuBtW8d0AldLRG0CJmyznS4vlni8mZhQUZHICF84qziDzoP94wIEu
0P57cditNvnH9fEavcSboJ2DcpVTJZDKSH7+c97WapnAFONpIjRaaxAl0ZHTBmjQC4X6ElkkFo5s
ewc4vlUaw/ipw7zFtd60lb9nuAegbI8tM+t2McWxLh9zc2IKs8GTHUGfzJPcY9LblovZYZLMnxXi
CeDWqebl3tkA/vkSJA0SrXd+A1QHunIDUsuhpwQZBAmlyiexMAWns58/v0Hmw9zZeKSrAqpeTi/q
HFdtPAifVC7O3091odRCCPTpL2TZtdsAve409OYUMrwwlUf8svBdKI9hJbYnMkBe2IB+YrLVko8j
HVloJYY8QfbqIG5CdjBr7juC+XnowxFuhkJYD04cn2GvrVLSGH90poZ6jyWp56my48Ou4cMqssI0
MyKc60WQNoiw2oAyE2MWjEb+wvYyAESWEluzFqrSYfM/AzL7P9PQUBn0rgSywBMM3OmGzT4xO0gr
qNBZYeSi5w0DU+TU7yUjd2LOIijK607GPRtmgYrIbD0TeflWbWaocpSHx//a/6uvwC7WVJA38nJb
jbGGcQDlHmCZNugX59XNqZNXRtDYT8yTUrkYvLMMnGGfitn2juqk1uWPTnV/kIPkj4zPfCephliZ
W2LlgfNMDLEotttwRRyW9YcS9nHH+3ZnUWH79OtsUNcVcjLjSJEx6eSuh2sbvWKJEniMnt+Wxvcc
ZuL3G80EDGAWp/JpnsBYj1oAqiCh0CzFmxNKiuJ9u6dYlxZRJlP/rM32CHj8601qCmutc3FA/MuK
bA7S0KPbzzlDzrzupEmJGFxUONwj9vnCiaZHcexOwUIKTrLC/QIKWJtAuMECLFnbmmBYhE0/HrJw
PgpoeM5yzy5Ou27UwyXBlRtBlcUEevHkvLQokKP534vS3jMjAHMntw4F+b8J91i9X3bqEm7tECy/
Gtu69tJMLeVwnAWoVczsCkpIf4aWfpXGM8b0MJPyvnFUToCR1tOVJ+LThslo/EP50nw5MnRytRDN
fwr2pLQ3YNcFYb1X8i+jvGb6BcuSRGu/9f39lcxATIkXWgi/9mEkeTTD0E31xeMiK/bAwPBtmkL1
NYFjTF/aVe0uLowVXVTkyX2oQPWgJbb9UfE1sasuergos9mUcFXKnIGyYaJlP+j5mTs2CXXRG+mU
CqJl8HkbVZTfFFhyE5nyQ20DI1sGUJbVlm5P87JVT5KPTW2t5cnKYMrulGCV1rNrxY0bhOtKgeS5
7MeOfDOcruySP3SXvSoQAgT5XstA319dHXfNhSAoxFEoW/Qs4La2V0IR6YbpfepxsxjTzjhPRVkH
0xDDj3//6Mem6heFItEkiq/eFA+tK9C57tlIsWpgv6Hlk1CoD2MJiDuYukaSY/pT8m1YfwFAdnKl
ZzY3B30HC+B3f6V+dQ2Kbe0BnToYMYa3xXH/h04/hANlkvvt5BrxOelVysS+fkJfTtCsNErh4E5V
VapJInkaqPF2TN4DanPPTSFSLGAMGHcMrARh0bBw1Lly3wgY80ocuLvQjyN1OGJr66xM5lgQL+E+
1QTIH6NDpXKs17cDpdHZBPDUFbH/OuekUo+bEbT0xAujVY4NFH/s0/sOvG0mds3sUAnXU6QfBN4V
rX/5Z5krzztcuX9b8X3MNpFicVnEniwhmdRec6F6zSU66BpcAn6d8O4Fye8wOx4v6yfH2W+H/udc
sbBPfOzTXXN2Kjlwec0nQg/wE5ziCTQ1IGvrPEcFkM+UhX+cExN/r9aMEnKR4q/GgOdzeAY4CWLR
W+lJ5M67t8QvmqSUwo6BgzveG2XGb7gahFQ/05QsjespuW78KOtizvx1jX+WoUGtTaHZBTL3LyZv
AXDFL3g1CHXq9mx9RbStl/+9jTY2z267e93S6VixvK4ATU3h7TUJ3Ht9t5AiyrNggkB/b0TUzQT5
fB6OfLevru3T0XHVLINxYQ6XDETIA5lkkRmw7/WkM9LR7ZokQlZXbUN9pXxDEWOvqtYV4QHJLQlx
QNYqxC3z77LGCzfgT5brRvAhlQdp27SGF4Ts2PxkyrcjcwY3Phv0HrcjMPPkT0lRE9DA3PO8pi+a
MRf1PqIXZscacckvl5MhTH3NSSlwQucOq6BuIEYFkoybrmrgrOaRGhzthJvI/1EdYky243HMkwQO
snTsdNFR3chiHcFyf+s32vrCX3J3Fy+tAAm0anj3nPF6rC5lOYPKIX37KObFEnm2DMP9VD+AOmAQ
z2XIBwbFlSWGCVOSlXpZGcL82ftFoHgeZWVXEfYgyFrs8Tn4x3WoacxZKRk6rw94Jzn8bUyMbXsI
Xhr7GRxqlqc0F+PL1MbGiSujIBAKFMQeVbzIOQSj3rckFPDR60e9NJNEM51g0azwzBsyV/pAAeEp
1HyIkf6/jDqV266mB931IqgzsZNBvlXZarzm4hv2H59Gk15H70oZq8uJZw/vmBlc1gyVz5wJJ/an
BPoQ0gTRnNM4YsOtSyrvca7aQJBVcUidk3qHcqTGki7Z0o19ICNO3TgXwD3ZR4uChUYNkCxE2kY2
5TG4KqS0OkNdNcyck5Ci4HKN/supq3YklEl6YVanttob0ChOJDJ7xvXnqdwUnmzhihKDH6/cVJV9
TOJHCZ8ezfEKrZh5cfwTdgmeUhy2RQTyKtK4AZ8wgc4dYCee+kHSIJQOf0FzluYv/rxZC6UbvZBh
dNYWXXdI86k4KGpbjZEZm17sc9KFUEEdnfkLf0VWtieVoQy6oM0sRpxiTXOQgoZnva+bT7+Abdyr
TjpDGVtv3bmclW6V81r7WUZmOfAlFTtw8mvOsraBNg/ENnpjpKwx+gsaRECmrqIswED19LCo+t/y
yR+tbeGaWQUm4ruTWVi0Glp9a6syTIupmp/KJuKG2WbhjifRMJOAvJuKYhycZEQppF4RrGOSezCy
5hy/ZPeFnc3N3pV7onvyYvCKEfZk3ZjiTVpfgSGXdIuppgeQhLAwnpje3zU+EtQ6Dah/qgLMCt9K
AqySQ2PEbNOWfooMxz99oCn4HuhL6n6uSozwm85XEtINZVaFpxFMwRmjpStfhkqXT87zcY/ALsCZ
4nBTQXcLNQiR0oM1nzVVNVDLi2lEZP2laYmW7cde+EDs8Ezwm5lPJI8t3DP/MEsgJWaDZakDo2BP
/UmE9oc/M6SnO4kQmYFDcl98Ze8W1uL6YwIG68GYzTPFw/hxPaLywwYqace3qnBdeOVgLsE6L/FJ
35KZmLiUPDWksDwlaKpAWhjZI+ZcPBMyDaKfbJMeIdSAiKZDU4m7BP0svNoHikWyWv770kphxW15
ftzWO0p7fSCb2RkTSwljkGc/UWPnsN8KOiHjo/TQw9HfxqsjRqypIudd14LMUIwkj5ts1r8FGGFe
Yf61StNwFvHX3p4BgHVMtZu/gZ/ZFmUp+UFlsb0aC5+tc3mQJiv/uiceGzBGHFerCCQSJEBSMDlZ
8OZOkbZNjeXM/i1hdl+A0AvUSUVefXnEHLH053jG82mfXXIzjF4xEDUN2utiNgqlYLZ3oDNkdi8e
IFQyfIju4fuCYXGT9Tjn40pjGn4YTHkhi0OgylKvJNTh9ckCFAo7+o/X24vVDJv9X4fUaiSPh0al
eFRUQ4d1hRE8Pe2RUXxU708pCdnBa5n64sUvsPpcIf2dQMa3mc+w90yUY6oD+mY2nIYXNgccrne4
B+K06krcGZVYIp9DLF/P/Gv+AxZc/gNmQpb9/7ClNWD07Z8A8n9dCYoH38x0jpWqrcO/8F4vZqMW
pZVDAlhAvIV3Icm50cVfmeCc6vWyKkWhz499IaHgszPooD62CsNI2jIXREprYblx66nwCRNQ+XZ2
9fF/EHJTITcgMNCvKo1D/jR86qE3d7fbBinZyuwRxsDNGh9hm9LO2TS/P9egewgTjdKrexYmeEA7
TFP3hYUQ3ZSXP1cpX3vzusdfz4gXZPJLvrUm70hN/inDRhScdcJLewVFbQ7zI/a605RUAAcHGbXk
xZli+elPhmh+dwjj9MD6Hg2jH5RYvKQ6T4h3AbSjPld3d9/NDPrkURNOxZvW4xd1TT7u1yRaSnfw
ZUsO5/t3uqDNgyP5CszPnvLkh2t4m3CMDUQO4VkHS0UngeoG66wanZgSWrVPw2zjazPvbgJWIVCN
a1Nxw3iWfdeO2lZyDlHk9FIWvad6IE1dcVR/t6BwNHmqrFdmx8eDOmGGezxh/7yUp0bL1Yx2M247
bJ8DDBxrpXjDDeTsCnBoaVR4fnBBeTtOTk0f/HKGm1seig4IQpM5XC2KFlB6Md4Nc4rQ9aECSIKQ
O6Irn6kS6Gp2lUz5KUGjE6dNaGC2eAxROlnC9OyW7PWOZS80qwLKbuA+Wy4QTn0sVKXD3cNiUWG2
uPsls+3OKP9OVn3gkpTo49SrzyQNzjgjtUOzlsqesNrftz/ALgNw0uULt/kmteiPSfIwufH+eglt
lNf6UpGjsQ+eAXZsLyJ4A0hSQg63DMvKWwtVYkHcxRZs+JtWVImBpMUvXoNu7TA1WnYX7UX9/wjO
SoubGVrUM5c4ShCFyEYteKnAVza3C0LFyFivx1VOR+fC6qfDooeZhVQv5xXZD6WSXyMXECARnr5k
xzEnhwRz4+ILQYWdCCaSzix9LiZ8qZ7Dj+6MMS05YLB2T9hn/Lwqx0/+yW+cY3DoKQhkTRBt/GHR
eUtZc0UXipDhOP+DlWuTNGQ/glg8xOCo6hNFEeegQdMR06WzDiTKoH7nH4HtcDm5SXye7y6LQj57
Eq91ZnkX35MZxwvKZJcB/eb/ZReBqSMdqmRXAldwXRCAKt9kMCFApFCPQtU72Q1aHyz3ALT4p+Jp
OSUYEUFjds7msGUKpmHYX7vV3PSGHPTvOcoNE+1Z7gseXrgdM1igHeMPV4jDw4n/yHaTjY+oCCGd
RDmnuNSeSlnQs23KDXYH3IwgelY/ySyF2w8GkYiHCs1TUduze1p8yZuucnxMthlHvTec8QdAc22Q
nnUHGBlbpru8ZhgWHNwnw9gjzGR59BCRW1F7+DGM7FjIJ/kBZ24VRz1lGnEW9XSULTBP9s1glChE
enLGL4krz7wcdGjEqF5ffGwej6N/aNGXJ2+hchbqw5EcG3WjKmhhhrABsbv8P7hy9UG2jvLb3/fu
N3e2e4gdew9GrU8x/k42WwOpRkVph3+3ArY5QEKNjSRoyj+yxep+vB0i5RZCT3RzPuwS5PNTzSA/
U9MakROdlc+BenJf98CfgSKCtnIy5R3hAagefT0sfRQMRphfk5gW3F9B+dohaDXaECr0wD6+ydwg
ZE4QNMGq0UFvmv3yjCMJ7oUyyaZQuh0wna1hAaNerZgez8KfXUBddC5vqByCJ9Po+qAYzMeRpIkE
cn9TE2QI3g+rXcMJ+L848O24bi7qI5U3t9L5XV1kKZISUHgrU+nOG4OedICVJnr7GUinPZH/BbJF
8yzxT4h3aodI3qJA9RM4bRllV9ZIkpQd3Vf5PE5+1hYXV0dSB24hzcChCLsKpMHdiIO6g71jG5hJ
BggQ0T8a3sjxUMK4tFQyuu2j9a6O6CKiWV/QxFQCTI0TE7B8qE6itrL72WGmV9om8efWZGl/ukDb
k3ouO6b8RmE35HZG0DZT4eKLo0ZYBnFUlzxDTvRwvcFsDtWGpIvaHONPSDDC57F+260VC10Pv+Nf
k79m1V1EjIs1Ka2dKBh+4fmEl2PhPQN/jzq+IdbmiCH2XdtKFMogEBW/GYe2CbIFOrernB1Y1vCG
ShbItIzicRe4U4x6Xeoz1Dfb+T6LV5whAl01twheqr2k8zVZQcpzHFA06aSR0yCIQ97npDhnPQq+
0FdEeKvmil+0v6WvNMzYDkmc7SJyheLYL5LQDG5m383QhxYZpfNuPkwIl/DYyEkjRkb7PvxdurWJ
zl70rT7PGgoJN1+NmztJK9EKSMPEFUJMw/sqlmN7dLj+IE63Jvwl7TelGWFQY+BbbAkssQoUfN8B
YQ0LsdJDY+mLsPMlEVBfFykoWtm79Sx1j55Yadqq6HIsO3jvArR2wKMh0Jy/z8VYUPty4J0iq7iW
cyqECnmrtqr5UitsJrBJHNMPUMUljxht/1N5KJ2VtHf4GaynKUg0awcRU93Mf1kPuCtF2TIV/fKz
Ew5EfJLWudYnKr0ckXgj2ipTNUOCXKsQ2Q1LCuiofMQH9scb3R6P4vI+IT2BqBZPj25Su45X7tG0
QxwIZVo91FEALrOyabwUIBA53fyHXcNYjxMFlNgnMRsyYoCKnJhrl0BT/e9NFByWdkyVasRrQ9jS
bjAUJ2xE4c8eUHCLdd4hLtFs9NXs8MPzNJK186xr1mxoDnmZYdsDehSWspkdJaZ3vWAweQDsseOu
MtKjehQRk6NPwpOFDrsaoTdTJi2QbvbCZE0GG096U8ZX6wHOTha4ovZwM0+sddymN1c3/SNDjNGM
6h5ZN5vz86xgRgM9bX0WscPkHPkHqfbXWY/voh2ihdDxcWj2hNMUvOFp23DjzxsSqpvYatEkXprz
cmhzah60tFypkP1+KZPQBEt5ZTd7B/L7WPkv59FfIw0GZaEP3bpq5qH7nEIbfJ6o+T/sa634Xzpq
VrubSzyUeIfuzkUSxiy87xuzPJzseLWBdgQL0x400dazWC8MVLWgYRr9Wr6Dnftg3czEfoGBwy49
/CXkBmvP9qE4SH7vP7zQOR9qK6VZY7ZkIEMtiT3pSkZvpJ4tR4YftcXIGlLDjCkmBzEaE+L7mLP/
QcC3v2NqmsaPMJbP/PcQYeBR3BxMvI3IuCC4fK4ut6SkduLnNBwJaIkm4K2HOgVoErlIZ5Q/OXuO
NC3Vq+G+twnFeZAEWgY3QE+BXDvy/8m+WXGceXEcYUDExMxHRcHty5x9BZC2SD30pgJvVPwRcoya
PeH9ng/RV2FmdDQ3u44/FJVnB9VhPykfYiHZyc0JAlNj0uh1QoawnHwk6EE+I34gFlR21+Zvh/OF
kL+a03FVCF7KWv2COQ2oGorZtmA0xHDiyZmbpIj+TUgmXLKKnBpZtNniWkKIwuykLVVeUXhCHHYp
dhEom6i2D7YN59bOupZd3jxNkip5iAR36Jr0wXH1RHEEGWxWGF8WSaVIohoiTDt7vMenAf+sMgkZ
rj2P/81B5C89n2McXM90SuydgfVjFMYBUj66qd/ChEX/0wus6tPF2L41OmBVsd9WPJqcu0/OQhRe
JVQVHS8Tty/ugeE3afRQgrc0w0Rc/iZhcm7o+q2xtsdb7aiONzqdewdvRpuNV1f2Ygy6u5zGbL4g
+F03NGYqdpJ54JHsoiC23R+ai6+5ZqL+Ehhmwjlw4tp7704MfLOADHdT1Unz1Nq8fNGdhqr/TExU
wIps02aeWnYAgWvvknBfBQPpMMPCn3Stcxx3+rChlDZ9aTGMMcNqUiDvOiRHrLq5L5M2zZZt6s33
a42OudPm5x7dvFF+8nRroyqfAcafBv9lOja4FtVNTmFcIMwsZNeAoqiAsOA5kUPvbm8QZwO7ZTnD
EjlfJJP/mOx5GyaqpREEHwH4NGdu0bgqtKgTMAcpapW17bJResapnYJpIthWqyPgeQ5Yr0uwOI6q
NV2rjkHnNJo9rcCfu7G2bMoqvEF/Mq3/62zhChQmtnFha58BiQvh5bZexaLtCZabIeovEf7rFNG3
/BSQ6c9GdcyCw4X8554BreGN3+2/BI/I60mCPmZQXyPm5Lo2wvOg7gEHLzq0/1WPxNRQ/4xL1pRN
eYz5cV7XxxRXV+0PP2TrlxV5EgiAIJ/kM7+gKy72jsM5RiVRS9k3fdBEgszYBkTDfCy+FQ0eR4uI
NYKoP5jQp54uhSGFIBe7ruMIKwy69PEXG1dg8LBA9g25rmBR3AKXpJprMRJ7Z/HYo22+odsdcwC7
jbcqh+gkN9tzGO60talGRro51d+n7YJoK2YZXEoKxm60IZlipgniGLGkiJN+A9Lb8gVZi6O9UFsX
kWImOEBoY0E1x9p+Fi7AAblhypLxtx9YXQ9zzjJ0F2BqciE/LCOmamQdKcW2hPXCToz3DdywJuEr
5dDu78eAgzdloO7pjwhw8BUtHBOPGRLSEqmJcKlJyVpTHC1hDZhaQGWqsap05iya8TwrlYfnu4I1
COyORR55tbXtXL0juqAKvap5InYPlyNbvEUNC4z9g26d7ehLOfQ1wi01ERD1HoUnk1wyWOIfr1b3
H2MShWmeI31k0HZEMJeBsQp4LAngBTykrP1dpznoW6VMHPxzKUBSQ4Gen/5s0s9GUm2QrecOxJHr
IBDPPmpGw/P8e5yoX6xm/yHG2VqFcyHB6EG552LGUSGfKVzU4nkkiUJoUBWGcldVPe0IrO8DAUHR
5YqkBOrstKYLstUdN7FAr9r7CUuHk416nM8WigdGhnChz4tCRX8Tvor2NNRR2cI78XbrfZAYNxul
7PIO/sph2AHQLur+uJMDehP5TyyyxNXnO1YseEQ1dukr2oU8rmB74omzp0XugG5aHs/IKnlaciri
60dSBoqw2mJpci1Cox+VwB//rI1Fg1YJ9wGMuGm5QWwwxPnl7x50Jm5LlE8ZIdjxhwruSV4mDuc6
3/gkwP+yvcqlRrHX6/owbJofO+im9Z7Jg13iTqc2t/F/yh6wMlHS2WpeGXqzBrQsjWqqtlCV+isU
x89wzu9PzM3p8Q2glUxnGD5I0rU9Scw9fUniEEjlhJo83W1vyUCHukJK4Dxfy7UEttOdV8iLeqBj
3tU1tVt2cZcAHNOV2nWI6KmfmYjPHyl64znotZqzDbSKGhAvX189fD6oibruqIVB9nuEp3aFXvh7
O580CuuEH8z4qh2z5j0aLPxTvP6/pyfK2CWJTnCMXy1QO2+xcd+VERMzkCVpS57i++W2IpeOuLqX
pl/iWeW5x7Baqth6vVGbFhwLuXHCgOdgUsLxrbWTMA3kV3SJwxzlieNIPD64MAZ4L4KDylt7zq5r
MT6FDtH4FL85KZOG2THv8hzPEkdUP86K6tNAZEkuth+rpXBZp7+KQHCkLbR7MbyYm2M1YQ9mhdZS
4LEEecprQtDqr39bxnaOMfvBwNOT+ppJmo1sa2wCQVLBwmtYC8/k2N7nYbr9j1A/DJ8e8DSrgIOQ
NUgqEL32VXgO7ga1Qiz1vWnVlYYhAjjrXiJ2yRnxhFJ2wHeCwC4efM1WEUMeyTjbHOdN63Qgaglq
IBACzwD39gqIf+6fnSr2o0XwJnH0Dsbl6U75bcqLo1bYuKNbifZ/uoliJjdy3NH1xa1Ozky+UfiM
GDpCC9DmFJACCUU8kuxhywe/Z4QLF+ATH/4ZBJOyTdzOxLstggGa8lbopDO5D8LE+WaRfpfuHtm3
4wFQRFnI5DEtuiqvpRywpdozt8hOLDbKYCERNqeUudBrxgfSO9XS8W/AQL26jXNmdFgJiiO4jB+n
fBwY12RRfCZQU3QBBkI/znZSJvZjvkR0SbSCYZHNpqmJkSpN7iXHK3FY/ciFAoQYvgdv9/Cy544D
rPBQS7hHZwAqWUf37GNkhscebP1jt+rbEcHnMSrtk8CZrxW9K/Kro+tRSHxutyNaVnONg5RRJPAL
4eRHD/zM9IZr4+QkM2UjfFLbaInEKmn0ofZUB9yOiMtfHoLFNCg1xBIcqTcrrNfQST7aIHGzQIuI
xjgWf+Yht19qGyyL6qR0ssGatjwAqRtLA2ERzo2mYEgNy0d7ysVBWRLcIgkcC9FqVr/5VOC2kRR6
iPvFzGxAf9rIiUNeLj/Omn8KSF8CcQ65HIHw0MovbcDD/AP6BAjYEjaYRPUx4p/7SRfCeXJWnulT
4JorQf9lyXJywYu3+mE1IawRj6CTtFpyRyFnODLAkFnGEuL7FhQxgmDqHJsoZKWXvjzeI6pazU1P
ayoARyYx2icZUWG0zjhixiggAyxxPNUqFKjnLuR8Yk/ZK859ckLDHmV7xxkKEfxuuI5aqSZul8qL
KP7iZRFWzlMLByhDR39Wc8+QVFHBbo9RZ8+77hvmLKzTTG/QQqLBduuBPLSWhrj6EUWBwHK9opqe
pi/jyKyCXlbYqlnRPElxh5w1ukE+tAFRodbYNXIGlUjWOZRAKr18+I+Nwl4yPiATqGnGzwDoRr+U
qb/wegjikuwJOjWdaUbtcZ4b/DWPB9mdcppnMTCfOJXFcyUfNWQmdHmBCtQT4884WJAkOeGSyaY+
w0eW3EMfuK6P8rZ5oZ+4P+sWSqsHrfWURooW3iQg9ucW6d6FzWRYqlK20Ok6JDFgS7yXi4P6j6f/
Kq9PYVa32M3unt3gGQ9yIvJuvnNAgm5SZp0aom3+6S2S72Py3iQ/PJi6XMVNgqluvdQv3uxg7iUi
9anwXMhqktYMPSiPtaDVarsC6sOGYh4KTsYJ+uRHNTbzkrnLta3/3HHHniTFWaV2uVcDjCyEEkru
x27vyDHvN6vjaumyB2XLHfMAPnFiIhFayWXILMgHpQHOpV2nRa0ezVEb6+19iZ872PhqvMdB30wW
faSLJX2+bzC2rnNAt19a/mEgImLVj/QsVTMJJaVypYP0U2K7VO/v+0JpBQ22Qp+O0Kh4hpn9RHl1
92qAVF4mZYs582y/kblrsxys90NJOtr3AFQNVg5vMJrNMGJvHOYWq8Hllj8pjb1iZSyQBo50Ng/i
+9bEYNjvAKJoyJKJBlIF8nprAshjpdGYf8kZYw9URsj9hIqdkZIflPW/FuXxHZWISW89rr4WyGms
zqXWenRalbiwzAExJ40J9fer7cuxSLMxgXI4xNZBGX9emiLNJ4b9NLI7qDSXD1QBrNb4olu/cvRW
9jA55UprhK0012OP2uO1cH/DjqDxaaujS2Gzk099zOcS0COqaLMCFDN0udgVSrElzyGa5P6sVT/P
zkpxZEesfnEjem5aepoBKaO/ZqfBO8iFuRYsPHHZTjDpwjRlLPq4/CjMkUTcHyx0uGa6uPUiLFJO
1s8XhGAtOLlyUurTA4QLMgbi5hkm0Ju5juJ+sM3tSVwi/FfMhujoOdT4m79v/fbAnemOA4HEuhTr
mvbMTPzIjHM6bqdNYdQPFu72uEIJ9Rne3bl7D0H2cbF9AXBUzIMPWINUC80F7rVhmDpMsOHxR3Hm
b2WplvDQz+2yPUkE1zaJuk0z+AguNmBqxlJsd1Tp8jibMrV5FthCSLGOdXxarQXNhZh+DpVR1TEz
/1h0JXyl36NRk4kGQd+UpMsslF2gZECWVr/Nzw05z9vBHiESMvw7/DbBLvezjC4hmUPBNhrMvMgf
OhGAGFMPmARqxsaeH5+ZY1vkBLFWkmeVv+sbzeKx8wt7ATGo/i/weK0XgTyV8mV6lZeEwXwkr5Tf
7Ulmqj0M8I4wiEC49P22niPNhgprtm6fKzF73/En+buZHpx+Lv9+suEh9rsIwY7bMrvEtItp82Mm
RqyM4rnHeMRoAP0Corawj+wY/19taRaqnCsb3ZReLYaIf+K2lfY85t2p2PoZPUsHBdtKX6IBaRjx
PJeyUfrs9Ht1r7ZAdGWiCjLvMcaxrY9ez6hvwbxCIs5qqG6ue0Qmj/kzTNRy6NCWj6Q0P3z7tiJx
3ptBkmOSmrWcNW9rP6fL6WEG5HkGs/Bt/p5woSygkgWuBdoigPbBNrgyBQ7Z2mqovKBwS8/tJapG
KmfNqtuWYqIoWO8XG17jHJrk4806iGkiI+nEsb2uw+NxBF5k+44sTBCKe7izBb9TVv6m1Fm1Gaho
Ai2LP0ahOCVeHyYj/InLmmDozWpwL4glcXveCcYjN8kqtwwx93iclP3ynA2Lx1ofGPmhgVPOOWg7
YutmhN7528UW+wEwhCT138pw3zMrnscSq2irPvmFe0YMJT9a2rJw4/4Y5z1A96nXhbaUfOpIycT1
pKH5bnz+0C9zNfAFEdy4rXB4HYA+JjPD1iRHA65ko+cKVbTmWKAkp3RDv83KYtWpHPHhTczAzhDr
yI68WzExTLuoXYPksURJnLlauKz48SqoXHdQJ2NcQq3hIMRQHdRsp4ITHdvGHiN5nSyUCJFQk3L8
84m0VP5qxkg0PAmXEJRRHv8Gpg6JVOhHVPSKASYUU17LQusdMdxsz57q861kTgjg6r1ItDg19JX+
Pw5EHAYckWwT7FwjZ0VtkeB95AEI1vMz8WlqPqIrMzx8ptzYIyxN5m3nRDqIBGI9sqGhsxpdnI+M
u4T6lfqq7jjhS3byaJV6IgKy64gu1GQFh0dKU62pRE4d1V+rdbzffMabuVszQ9hJC4L73zYgmggO
yPJGqG/X3YtXxEAw2BhtnSD+DM2fBDFdW+YurQxXdhS+6LP6cS06kXph81DZEPyUw8780kxipjOf
Qe4z18+C6s2GIaelWkhB0ozItl8tZEQ8vdv1IGZ/FY05UmT4/clMyNMzvjxie4kr/5e39X19Odk3
v18JeMUAwUsJ3TchSjVu0wYVm4Hv6PvANi1sweJGYfGO1dzLQrpFYeFAx5hxT5dz0PMa5tGVJfFY
vh/0e79Z8rAVGZlHL4tNA+kAAx/oCzrBXb7ZExcLlhEne8BBBxVjGxj/4L/DvEC3lwiJcycMRNS/
20b/S0VEJt1FhQK9DQPmNObhALtR2t53QbSibAR8sN8Hx/n2uBBVULqc79q0m+EhYw+NtQDC0sFa
YKY2Dzn+r2Mlte6CFPbfivI2c3qgZWHGIO7OXbqCHXxa/7cgAxiGnTe4Z4bNsg+bxiUUKnJPG9eP
0pnZcY2nuO+L36VzJCjoL39ohFtFRuGIH08scOTv0y8Uux/UK0u5adZjr+TRlT64SEzbCecC0HGB
Y/ESpUKd3Ukl3rP4zD2fNxyGT+Ad8cil2UIuhIItEB7hjPNTvpgrqSYwUtbtzLAQPYiJAKpZ4/yu
t3Ki3h1pLNs6Bs4z6yWBCM4UmCNoDb6ddorMH3yIrbbQZxY9vgy/TwZPf3NH+RaohxlJnQffXdx5
zyK6SZswMNB+Sv+RC127yhsY2tfKeORhKIrVyRyzEuzWBjjgPE9Fja2cAxboTzhvbEVEaXjxXzxM
+BLnx9OdydF9B+W4V7xLZ2pCaGYTNHvRpWV1nOcJZsHP0+r/EWSH1nxlX6Q0lbLh5XAoDe1gspoc
FKVmcgNWJB9VdBTDlhLqRWpOHrwd5np3WSAaJfPmSaZkvCMSztC9PNSNwrVWbQY5etkO5w15boKU
8nSveWoPgbNpnqTI/TO8YSoNfqyIGgDRPkd+zU65dIs2c12d34C0nBJiazgyIDLgWogikKWqVDSt
FyTKdehENJF5F8rVcnhvIJxoElg2wkENmXLK8BZeE7nAily0yMire5AEZCukmz0AdKbptrvssnhF
oUtakCQ9HXKon8y2vfe869OraVNKk8f8Uj6CefM85xWdjq5qkw2eqGn2ToFM7seod+Kdodfi9qu4
JRDD4GjrHGT0jg5UCi1KGaRUGzoLM9Rd65z7DZr0/P+9olMUlXorehqeiZVI7Sm0E0+kmXa1Opf6
FR4jNb3n1dQ+ifgVZipvODgs3RswsqstCtteGi4x6Y4pAG8Kw0pf8JWIebBb1nKZ38XEWwI5h1eZ
9/d1At4REVkejN38BnYJLaIQEHmtfe7oNjsDai60rxsUdRCoKqaxYUkajF9ZD8P9bA7MOZnMZPwy
0o3clNF2AqB00jf5ORRe2lbRsLM3+Z7tweEkszkqjLsHjf1vnBNXUh9NUoZT5s96CBaK01B8BIaM
l64C83T2uXoGGu9T3r/DFUeJ6pWEO0GnAQJJbY4/9hpSEeDszv76Zfq0zGwc7Jg9onsj3zFyn+HL
w4pKQDc+4d9J7knBgpkASb08Z2JrNgllbbxqoUnjjSGrV5WzSjxraLLGBAibKe/VGwrTB4Tx2S0o
whSGVn4rSMd4KNpMTwgxx8eA7nG8cTvXFkajqEzoQNmlSeou3y4qqPst3N6/zQSjR7hk6DSBlm9N
ZCYSDTSmpW41y6UDBPe0VN8YyyuoEUMX0K1JRjFwPRyzIedluFZVSjpoF6z9RDQir4Gk2pHYWLaF
LJqv43HpwbooTeRG1pPVFwxldpd4bdQAY5O+GeAy8oiY6TTaKyR1Ru+igzK/y9lztu3rZxtA8YYb
cPz9PJqM2OyhI5fmq+oc7/wp/FBUjP1u6pyuSCAQz2n5vouLtc9C6y5Jqa4UkG2sBfVp1ck4e7/p
KiznfcIodvdOLSXSJ+pVHyLjOYfn4+oMi1b8OST1aEtYEGPgLCCoXNADeoaaVMYLr7zS2JUwDRps
nHkiAbXXoDNbRF7GjBbqvx/B8a3YSYAtjRxK4wIiOkj57uC2eTjxbNgdKtFJ7RUVWVRa1agG4z0l
p+xNY7CGMQ6dlmhOh04HH0DeKTHQAqNgpajqKH6UsYaP+Pmjr/VC1K3UHSMAvBWC2LKm+vIwjU0w
c0nubfjfvFaHRyqf3R1BLulU6PUB4mVkEZMXkzQYM/FJ6t8EgLknbmgruBUfk9Gbw7meEqj1DLs3
6/yogKOau5YD/E/rhc3HBqo+apMfwkWBEh0yDNW4dQG9Wm+e7Db6wqRny0EKmVoX6xQ9yrTwOwNr
CAwnrQok1OJFG+8WsfUtCpErUO7ufwpJl2gP4pGbO/c/i6sN4R0rampg7382yt4Ued54LbuouuL3
WhyuO6oqVbd1sG8siv4yRxmRFqeyHzWEMe8B1ZotK58YlEZnefBh5GA3Hio7yI1/LqLomrvA95G+
ctdGGbVgDn0I8RD0yeBIFZgMae7O9xa7B3hterBT9fQtpKNi8k+6yOVeQkmxBexZyoyNel1D+xAk
vxQcJckkP2fTO3ndvGCDRtiqmwZcW0wUZAXleQIfhkikePuM4y1gObd+IRNCvqj6icaHsGr4AqGF
CWOgCrnb7tX9gB+gUjBieU2LC1ZSwwf0vBH8hrHMJBtOTHMjnZrBap2z3s+MuBh5D4jpfP93V+6g
7DwMQciHGLfAcpCQP83YrukRzNS9TjBLQxA7sgwUxc5tZnzeo3VCWG5thoyhM5DVyzvcIIqkgeZR
V1vjMRPV8lVT/lRWoEmOhRLq0M3GSlqZE562SCLQBB90eihzCLfeYb5VAySVWJbIJObjT5asxx6n
PCe5+MzQ+g2UTDhxSb7VDMNK5XbBFTUbgP2KVvMbMZLsNr9ZkRbaUCYO2jS4+e66gwJzk4BUJbMB
jj7Fj13YrxUhJLtbUk7/IWKoqmbzMYd3W/trPxYijZIdUdRYfiI7ZbcKGX5ucfofYJW9qeaXx8Qs
YKUlzIVxj1bQtxzPKqdtva2ZnsleNm+fiP/ooAbQNrKj9o3fVHpWbcep6gUkf4ZYsPhzpIcYHeed
ChSjQbF7xTin/7m25Ww329mshlaJOWLxT3nfcKASmTp8z4GpG9yA1PJEXXMsRsQ8DARU/MRwP1Qd
0Tv98hVgkcTGh2P3Ieeu/jqX1zVEyLsHQtJB3zNVx9NAHlCmDE8HYg7obptz6fEN6HFfUoEYRPqO
z+XAdpGw/UjuEk4PM8/gEHdbG9myHC/nqQC3Ao8MLl/lksruTf1OTBtwLX4s7jFFBsrE1eVG5dHH
/evgduUxZX32ka7ig3qCle2AHN/FT8gesa9k2AgztFAxfdCoaiknyvKFnD2R3z3a6utdc2IG35Dc
F7sH3NqSETJz+Jt+LcpmdSw74HtVp0I9aMeBQRwdrBx1E8r8gnrtZAZDf0KajtUW0kZphQEpWI/J
un0WxAVAy2MiIa+0B6OoRGl6hKqtHTpv+G0OrAQ6unwLqg9gTT0XoRL8wo4O/ebvyM7rvz55yXnH
8kg+rbepve0u8ZleXdMfmjhND4pjnMV/stQOWMf5zce7JI63NkZFEEibCE5YWQZDyQjzDhTMFnrs
HCqzNWM+LgKwWGOmJTBBaYWOFwg39hrb/7fbOs5pNH5aEcf915tMsPjrjF8pjpVM1vi5TNqiyn1J
N1wXKCfahNs3h9+H8hv+MAeZJMgP0RyiLWLCZJMl7zn6xjrIFQxxcBF0Mo07RbJgVUJ4E6/ZbtS3
eHDX1Jk5K55VuqZgaHT5tedZShuIf/e8naExmk35Q+EIXCFXBhC83jy1RvxT5PHx53a1wkRa6uMS
1AYvXt2aYMBVkHHO8uulpqo8DNmfW6OBlploiGnbUVZCWUUx1JORAwbd65+0FsVpEQcNLRKUsY2l
U+Azc0me9QkJUxJOqllLK2MXFvXDCgraRLf1n7GeSO7omCSx4P0OT26kjetTdxrxbd4+ABCmoTAh
QDF0NP0E473kC7z30zCsc6wmoFbu5SLt5LB5TDUbQtVQAaBKukOZO8G8sx+s3T5QD7NFsPFSlxkI
T8UyvOtvT88TxnYnn66w9zoDA/gh8cRTeBMsAz6WD2OWQaY2py54YBtkyCwl9Zf9aMJ9v2WjM58c
XLoLVmztKPCJgYD2YCMFcEZ1IqaBTGqWlhA/ivacoQUfMMrTfs5+9tYEW9fYMKAkEewNQgV6Xz9I
QzIDl9hNNGll1E1Rh2ijQd1YGDmeQjcgM2KcfX+TeGbeJ97Xp7hH8pYnctkhJApZYe9s8YgqWkea
aDjtE2RbgOdbsoniATcVjPhLDCn75oMOFp3U8HjiNpHjrglJaBjDKazZoDYcqnbAhP7wxmkoaDOJ
CpWRJWsqFBF53kp0eFfKvPBJZpY9Fv1TO49A4GhB9abtXQi7U1vbaj9Us3MmhnZZZIlioAPgvvZZ
G/HQtUyyXdXHwnpX+lqsNzq/GKeQtW0Rn0L27ur3OMaLv6PaAmBoMWd5ErzBkrZ0p4AvVGwTBd+N
y8YZquz4KniYylblubr7OI5Kwz0OOdY6RNiGjbFStyL4ZD8iJg36S6Weyf9IjaZbhPYYy3TA0VeX
flyEMBjM0x5BxsDH0lVGabDDBFWLP15arYXjLlPUfooGcJ9oeYGDvGNTn0O7WrQGcSAo8T3SqMKS
aImdaa9VL5DTGKQmCek8aXZirplKLgToQrAZELYaViHCeUmUGPfD4U8WaBw/uEQDbw5XLCxm/03f
T7RlS+mTuW72jbOM12jcYjBCnV7+Cf+FbqxoSiovkqUwCPsF2abRAXibNo5R9wZJfxNOYqwJh6wd
qMC2cwRO6yCpXCxVlFDNBioNS5Q+C1u54pKe5Z8OXjARLlLzUQmlGIvtHZTFU18Kw6nHcA0I8YKm
yej9eGDVqmX9IoUkleIQ5IrDyS/4qyKIhJFFzE0jUjkkx7eL5vi2A5l7ZFrmE+f5Kwq3aINXVQ/X
oe8/QVedNfPB/9OcShu27rrstosAcI1WNxFJ4mEfGcSLXhtwkFjyHFY8KIvcIvKNg1Hlg0hQvLhm
o+NJjyTXAwWg5tTLTzjWPqVQop9XB+wZF1WZ0K9Vq4NTb6zrluyrfRmjLtxMvxdh3AWDSK3DG8iC
tTVRTbV4iO5GJ/rKCQf/i4kHVFTSOZwuqnb8MRXhNW4EOiR61y1UZsvOKkJKzR3fuH/9Oaws+ffT
5VxGBxCfFr6tqozqtqO1+5iOgq70sshNGWB23BwNXNW2usV40B6UknjvmQJzzzPxrBMDVjlb+wjG
z/Rqm4AHy/vlN//rs6vAgwvyTL6pWombOuK5GdNr2PTJ8T2LefN3HG4E0+M0sv52E6y6F7MDyVIh
29PTLpexcENU7a27QPBwkZeqformdjVZk+ElXY2TXBJ10NgOBibzbDTKuBLhS9JxOVEU/QCwTR/F
zDVV58Ye+8aCe/Z4l3wBkwgXWAZFQiw7FdV1oRlNFk1rOm2owoCpjIjJK4blxtb9INVHeHdBmUid
K9RFQJMnRa6ZbTzlZYsufq2OvisTlevIVECJns/rldyt9LwNzEKR0u+Dq3aQIFyDcd8B0NUuPQTC
AW66kEKqo7AK6bEZO0BJnJEEPfuJKaqdNYAFhx3UTGkI+ATBdV0kfK3MQ0H6xbspTgUJvBOTMPv3
zVOzwN1iMb4Q//0xCPd46Y2dEPbLiIQpvwsJYtxg6setxxiNmrtvvVGziKC6blxWk/UBBiSDRWP9
Gs+uhWEGT4zmFPQ/F0P0GbDe74/kZ92YB/JqDMSTKfbJcF4aegCBAO2+zoSquqJ8hDlLgerBB0HA
X7rWK2vLE15c8A7bIwIdgCD4cMjrBq6rcxzSwA2QsjByfEjxr5saLOFYWpFIQxQdaDCB5oobeGT0
jCY0gS59DTSNOFCS1Q3g9Q5PQxv/1m2oekVitSzS6vaFYv1KN/+110Ch3Cy6fSTNbMyLNksm+1J5
MwBqn01jjNC4n+1aiOSKLpQEJzQmRWuwGZH2YzK2OR6QEmim8dNdBlmUMe33f9q2LOQ6DdAwEOk+
+uJvajLfQVgsHrlomWn1F6kzbYIxFrqJ67A4N0YRet/207gQrIyl3zEKaO5dxA51GY+PB0vjWrjq
Hag+uJTxJ23NtUICVI0BmEWpe+ZO+UAjaT60rpxbK3Ec0qbgeBGX3DVzqglvJmQO85UpCeqO1r7l
isZKZJP1IjF2tqhM4KLyhoB/YR7JgQ+CyI8RQExRDq3Bvy4MFiolCEB7QA8vErUmbcMtjM2IFivh
l55Bo4EOEPkJfgYKurlj32ZA9d8Qx+/Y6JVS1nV/MYCVY2/SwLvKRFLkKFhKQDZESlCBCQduvUPs
Bn/ND8BbEoB1jcsinIG65Dtcp+5m33E1SgvW3eCnBAgFwkE4iYp6w2sXwH7YZj9N8RH1HD+5ArNI
rhLOw5KWVH/fiL5+nGlQCgjghCbT/2tufndU9vv4IWw7QPMO7ec8lk4cX84XmZSApVltMuKMTdQk
nSvsb8/zScSpQBZf43zRwRpgnEgFS7jg5r/xFk24Tc8m45DJpaAmMATy6fgVQdYSGdmtUcPwKFv6
GTFsQE2dQjrVCXJI2f5RVG9Biqqm5IKxr9w6S5w+qC21jWWTA1UR0Zk0p9uLTDPnSY9NdHO+ws1T
EnOiLbF1SZaArgdmUPPokMPQ7D4ceWSCzKbHSHEYT0vA/SGcalokrKmXRkVH8d0UPIPKSBMH4cRQ
PPbCHxkpLcKZd07K4++/toziMPffrA7ZWEcdRzXKVC8RQaXkjT/9O6JcqOxgKNJ6dXkEeNab/Pw8
TOsckcDoFPnAvE92fXOuo4iKjlLkqB2kq7TIR8JccE2yoKeBXc7bO/HtWoQ3PTECNa/lY5iUmdRs
Ag47nF2fQq9bDpsQhRtbBOsk13BfJhGHPwjTJVkr4qKVgGvY6P730ChVnTxMaPXhturvyOhR84Ft
b6A2lvTj4zymhFxWXE/BWvCOP2zVygKj7QxjNcbM4IB437PmaeFSQuyThXl1OBJGpjYLi+OTJrWM
0Yt4KMArAnHnKn7pFGis0KJc3Z+g+J4RjcnxYJfMH2YFJpBcHM8ie1mF17VbCbhIel6Spp5wLWKS
+HjVuzwLdV+v9yXX5zf5wwqwAMlPtIySHinxf8vK0vl0/q1ATRMm15u0K0iNpTQ52A+mId+0PHUX
1kHewex8KO8BuKnjRcARpj7ItnTy5JDcI4z5kbWYoaV2nlfpaXlR2tyPBUmBXN650JeSPdR6NOPe
YG3OKudgy4xOh/IfnkF/tKq5HJydDRiwdqRFNzT8z7oaBApqcVKd/FI8Pd9CJ75/7qQjS3vabxqj
USQElOpi7E2HLIvK7sl0A2XOE1LEMHLrM3DFWUYEnmaRwFfxMEfn5MIrxaYPLnBHdC/iIl4Dpiq2
dlTp0RvmsqLHjQEojZTIQaOxdav8V4O3r7clG7wPDhzzvbQy/vpBeXBu5Gp+yc2mKFFNJ1BH02+d
975ry788+at65lRah9MNIhkIH+iNJGnDEDKqxC/iiEDIgf12X7hZSdQYbIZo3j+9HNa7zWyX1P/8
ADl21AULGwSURtySSpkpJX6OrCqclyZnl4xGWuPj915bz0uVUcPLXHoyeruim1W5Hc4NiqQFO9Oc
HjVIaEg1uwwxMenYjiWwGmeN8XIfPs/kVdJQx6EywdkDkU+YZv8RaOms+UcaG/BfEi3uJcTi4u/6
zx3RRDkCEusIBsbjuudfBsKEK0JFCnA7WDzwrnS7P56782J3WgO0/ufxg8k4PfuOd+utvCAgYJZT
YNBQjtHR64lgqjshEMQMeEKBMVsMOFDiOkSJ+x4roc8+K5xZ9qnsSzUV4CiqTryiZauyqy1ROPMQ
jiOtKbFTMIz9cFBmC5hd5X/PjiChxnwgXyk7f8WHukoCV6IQcVQOFgMd+CPNw+lTLAXNiopBUTy+
xxGwW+2jHjsr7hzOWmCBrEcjJsnRGIxidm1vqGIeSuBc+6he3zVlmBRK4/z3xyUUiVP53elAi/Ao
RlFm0mkEFGqI7NeRy8V1T1qUox+a58m7SORYLJsi+AmwwaUIJLKUZE4a24N72rUt2RDR6JiWsYcw
/IXyDTN4ZLmoBk3PtQZJ+4MIh/qs8RFHFtn8cKiST3nBUrvSXJHlVIIN6ZRIwRuosYtb/Za1dgHl
JRMiEQvDysDIm76ciZtRBsB7Vsnew40NdKsXurJknwbwvIkb1eDpU8qW3vu5fnIvqo0I4T+EkD+6
qirNjShd4mwPErQj45UWBOSrsBNMtc7tRXvCBM4eaK4GgkAsuRi81de5CpuulE0qylOytnOwYkz3
8X7yichdXZsnpBU9jvk9JttUWicT/i/w2Xan0aMYco3SwaLDTrou57rXvW6s08tZp23vpFnP9vDL
sPlo6hrXT/l8++kPtpvCWkd51AXRhHIt/r6qHCpxP7SiLzjvhwEzgRAWZFzo3GscQ3WTUn1joPRO
eFBz0WmuL4zvUiz2NJ5cV98DQgZ1BZIqQZpwzWXIMLO9zNPB+Xl/cyS4LEREb16PuFCo15cajnAB
F7OYUZYMT2N85fPqEH2tLlXXzPC+OcX68yvVkNfpO3j7aG0htgGnoNbHZTlVbQJ84pNbRzMulgeq
ej06tPxACfkJ2YMZh4Yzpf7CU8mknkgyVGBQlRWfuaP04AmJ1xtvpzxYPJ1FHHlpkXSNvyi0uZcB
wuvdAhe5J5y4NBDjr1cUJBVqW3063ZcKWGgc7G7ntIupI9bRFpjta7yWbPu3G406O0m8v/nuacoE
HVTACLc5HnotSU/AWjiOlr3NSUtkmDa2rqsudayoJXGYkSmIMqAC5Xkdv6qIhdzFHCjVVoPe+PdB
bqTC4zxk3kJ723mLW4ATmPlZkLfqUzC58F+k09FQCKnnYbLZR4Gii4AikUZ1556URLijBh3HYGm2
aLr8gUxSwDzDaCyI3vJ1wZUpUIh0Ao6BMwG+EkS47S51wpMAo70rjMkpwPvJOUnd3FdYNCDB3fDq
P+Xm1qeTBlkE7Rqb7V53tXCnYk8G6omsmIX98K/SY7KC8Uoo25P4ZyoK/v0LnfESjqk070kIVpi8
YIqCfgUcB/bLxYW/ugdhUxrrA08AFvBtGxeITCdi6XL36Cckb2ZiNKmYZsqHaW2SILYYOD1/R33M
r8eK8yfZFLxKcb0FChnxFH3nreutGoFISu8W0W/9YHO8ujpXTf6dTqBVt0jwWDn4TrjXLI1HRREW
5afU7+M0iDeYN9Z4F/HKv0ZNhXxp3bBYUQ8h8SOGaD7C9wXAJWDTs2a7nCN4sktgMSSNb1jnybSD
CCez0IxZjSz/e9v7lVDJV1SWEEzvd278LLTp1cvBfTlZBry9PikguFaCST7VE+msXaSK9//fJ6Qo
zlr8EkUuo0edDExnx9Pj5Klus1utEfJ1fAzSdGbxtvJbvWbcLEE4O/pMwrTgW45dsPpe9w2aMY+y
pWbTqgu9vOFtqtLU2SIQdGKhCdevLQZdb7QUPz005vdsRyt3AYNhwU7foXZnNaWOFwednygyH6hy
v4uxaLm0SvkJlwi30lPvOOLvggGg2WbKvCtJHRTqpX6qSU5NLq2901qaVCGWbe7fI63lgSztpZSz
itxUkgZ8AlUaENmPN+xOkGeCKJiV75Kj/l/ZMA/zjxG6X/0/X+BO4CwA5HKhUVrm65jfwvXVsU3M
0+srvnMTcEnOtOBMkv5MLSlv1EtZuQiolj/BlXWffAJ1bEkUh+WLWdmpr+/VTXONkj95vat41PEz
vBvR5PwgLQvT1Lb0jTgaL5jqmLSau6MRJ6pVTB+KZkbssoQXMMhFS01fjhB5TeZqpEkikSYAP1B/
2bAuKceEoNpnwKaQgYiveCnS/Mg1NcmNWkq0O3eLgvipvSx06LKLNW8/8zYttBNmIWDbHjnsRSqY
KAQB37lI1B6qWaYz8gqDYgy+Gyld3kw8CfANziiAclyhVR6hX/PIEZRBvp0bYBNzEiXmxS2tl3u5
xuf/IUq6MFHyUlu2xsE09edd1sMbpToZ66I27jpRRC+vblRAYO5mbpQ8v5gY+hXJA9oAvstfGruL
Lgvf7X0swnGAtYw6FJQGVj8d5Xwf7WIXPpbT1k6it9rzjTLWFlx5y0rb2oGK6AhEzv2sxnFr31/q
7Oezrp6dHIu7cnE5DUHNLiLX6p2V/RfIA/Z6cIaJzQCYZ4/LzNwbErtoDncqclrcfQXhtdwtFdWx
RTZDQSDeMM7cXNYBHObePZqPuAJcqKyMWcrrFe/Ys9orTq2X+RXcp8IQ/6arpbkCjMPx2cxIbev0
RFaD1yX9/+fZm/PoOaPXLfJdrNmRCwih6tLrY7dHRcsGRxb6ZSG1/Re8vb7kGfyuYgzUB/6DeRSI
18m07tYxCdNlGEp3pKZiHUKenqupFLsy9PWjRL6eZAYJU/1keTkPi80It4FnKnJ0Lmi2renwroVr
nrp4mJb1ghKxGHw8Bdppdur+KiiMW24l+Iwj3zW28NkaKAoWEE5YpXI4nb6DrRCd3rXKOtuKRQCK
JCeTj7CihSwQMq5GxWdQCFcPrmsYpJwAGSipCfdpD6g4i/gS0JmICxYwmVehhoh0/6vRfrPBmhyh
5amri2QzK/LKo93KLWBx8d8lqiYJDKwpNGgHPd7+VyUBLqtdQxncHHsT9lIvedDQVtOd/Txr79+6
M/LdeZPB/8J+p/xlAm43nypjXeBQ9TbFXNirFTGjV+n+x0zH4uDpnZvny36bfnKOlnAMOj+M0Al2
Z+W70ng8fQXxt85ZbdYNlqk2FXU/rVzN/xK/hnWIUvCZz63/JQX9jHCCOh7VtQkbinPB/SQAQMsa
FKYCgRBaltbB8iz9OB2hV3Q/FMyQMdxqYjdcQzQFyzk9XskexPLsXGLl1j2f3eDGqbg6EGW+8y94
0O8e7aNzJD5olMsrFawdRtiWTHgIbADklJuzxAUE9PXQa9Ux1fpnUkY3NoZIM2nh0qSzBRirAkha
LhqkTy9CfpNls5x8qA8oi6HqxVYCJdNs/K4RR1HxcjH7snY1ZUHrtdvr+pwYm7MT/3waDz9Y55d6
0niVThT8Uz1vkjBRaNZb6TZz+I8FboYdh0dOubYQPvUfvyWr+l5SR6ohkNEoQtDK/39pgcErgVpW
1+PDT7atb8eyVRjGF6gL0W7HuB3xSeLcpYc3r1si7vM05BF1CRRq+ZZ0p3m1yrqV5oB7cYnZdY8G
L+Pn+mSA+CUAZXfi9u7i2Q6zF7HvwAjCxWJamlP5MgyEWsDSpEd2yCPln7H/t8JgFgdKmEuz44ss
kRBRTcvAimRy7D6t8hqtSuWon71WVVk21OjfcM7sHpyClQ2Ije5EP0PY0kDmOIRE8aDI2X52H3ti
cx6xGyEb7rGYPFAHJ9EAo9g3Ac1maiMVxFk4IerCKasO2gHSHO/g5ILcj2Ct9jShm3/RKD+sjJj9
MRSiCQNkQa7RyZnjEQqImoBHGHNW45PoYxjyn9ORJtAEZB6c1DZzNU8WD8EMq9TUh/6ybXx5HDOf
xLRNKZiJw3wd2IJZBbXTOovN4kMJlS2shyRz+CiwIzo8xyf5MbXNopwtJ3KTOpUmd2mUjjYcQZmY
MSnrAikrgi6k5fa2N3xFrHc8hFbCPKK8l5iUcKYg61zpcNu9+KWqK1A+x5/ONG8yzuc2TWk2ULrN
71NuKpCbyLBmqs444m3x0m/5DqE/Lk1mpv07u1immrFa+LwVjhMyoJ0OB8j+wc6zsVE55zp64Abc
8osNDXvlThutyJP16W5IzEtRcOJkzX4rzGqh8+WwbfmQHldx9uVcGTPpykHuxnMplPj2VpcaUiiO
zqYkYhhjgSfiJGH6PUCkvzfX7AgUSIUGClngmr9uIR75WLAueQmsQcP7p3n4rrSmEthT4Z2DtQ0i
v4/KTh1tq6rBKhVluWQLQzyKWIVjCqjgi5Mp4tnkq6hdiJVlmJCVhT3n7Sp7hPBDSJJE/6Mhfv/K
p/jG7UyWjAwBsZqPOULKYPsFDzG/RBnxNSSdsyYx93p/Sd47vSWeAM9mGBcqnHDTdFeAn7vq2YQk
ugVy0GPMuBO+LtRbXhOgVKSlxFoiLwYnaGRddnlyAFcvfFlbKaZ+KFKKqdUBs0aJM0eyQfFnddpp
fQCA9lnl5R0mjFHez92VsFaTfrPUZfCYv7obgE0/JPtKrth25e+q5eIStW8TNMVI18fcqr0dOflf
+oosmJP1+prwWFnmxgbtgsPB4Hzt7O7dk5s4PQXqbEa2PHhQ+Gu7l54peVTdteAApRi9qunrbff/
cn9JZ7dCPnwmp1A2bR2yZFnUClT7XPQ5f7KUKTqaFtd/rlLOAEMkpnBeiybLdvPN7BmfeAusfRBB
4zhgUz2BjjlvT6+NciNihqU+mY9T8/VO7y5BkQEX1oOgr5rgY/cGwqeuJ604wVnVCvZVv4XgnYju
HleoqRnmJ50cwiDKM6JiL6vbq/nyA0k4338hDn1XWn4z22XS0ZzUVyvY8eDSwwlnsuJNgd9ZN9jQ
bvKRDUwqyTkxP/PXncAocyUjXL9wIun2SvaFzYzA0vJv61TFEHHTYj6/lJKgR6QXoP0pONgxuOhm
m2uO3sg42njuiH8XkpriY/MJD15wMZJ/2tMB03m39t1E7DpVCjkxwhRQh4AMl+Bi3e+cXvGSiUGe
6msgO8P4ZQz7+fh5nAfjRat9ru1a/pBNo+sqUorLqpLIP/sgn1Yw0BBC2TF/izzENk21w+n0Tcks
wKuFqTeafQIIwCajYQ+7YBzIe1GBYYDGOtyeY4dn9L8IEATZSJT2unyTzBJjGg84BG4tGCA+sina
IcjomaEF7jLiislMu4NgwAlE5Xv/n94RXFdy0hhQLW8zNen4f1srmJLpCvMwKL0+LCOF5BEzFQof
Y3pB7984YGKgM3wyx0dJSrmcDr+DO5lkO2PvVX/ns+Iy8QLQ4bSYEbqsgyWHEV7c5Pe9DdO01BPn
R4wF5cmjIpckA/mKEABotxMgfZ8W9DRh7Mssb7LWUYnablv+h26ta7QTYfirxuzcvHPuxOzzWBy0
GASjGW1Pm5MAkRH58VS6JLU69rpL3bJEDDOyncMI6NCUd5slu+pzw2RkfS4G0o4HiBIn/49Oe1aL
yMRorE07z9rpWlKqbJwvhN2gYGQFi6N1tABk1dvIMAi338/PhnxIWD0UJqMI5RskjgpQQXsoz2cO
Nog4Pq7cCbeDHZRy/4KLpfJmi79tK61ucgGlgdf/OldWDuUmK7g3Ix1bZXOb+A7FiqVPf4Fyj3O2
dI+UobY/MsH70C3egcKGCLpjh23RGOM5p0aLgKnDGGKfPLq/N3BLvrGz+K86FfAmWIA86ZVQdT7r
4QH5ip1HXRYSExezwIBvv60JoVDiJEhVyIc6t/z1bHcGLAjtOFxzwdRIJh0tF+sfxG/ptLUOn/YE
b7hVs+pUk0y026Y8qUdjHEBdOnhtjYoQWU5vsNE6apY/3QI5DnY4UnKag2vWKLE2DDFM/OqkOhtY
uf/paqi9WLzmUjsGj2z3eBY37KH8lwlJq4x6YaWotDIyOX1/wqspEOifRp49Fo+9AeXLosII5a0A
BtidEf0roHPBhrN364J3/kdfmgKYbEUXQt7s9EAa29VLOfg/pwuo/SKGXA4K2jZfzbZMo/rKnkh/
IAj2LGQQdb3/JZ9c8pfIGCKpgmkIwHkPXuiLQESziOEyDahlD4ve8LrXc6SjGYK9rcqZp98U3kVP
OX9kwy42Wk08PPqUYdLGv360hgg5cHUIOBRyvvKfFVUo2CGcnNCB4ZT0ejwMwRFy916lPhI+ZStI
xWi8gABUMFrXaPizv3+TTKnq/d5FRhSzLuTFLZ7LuwYD+gJuDEuJGl4IL4SD2bOMTWCGFZykRQqX
ktVbKG8J0BVehzmONCD1sO5eDVj2qPbtKhwQlmyAWkHm5g8sE3giosfBZsfMYtNTqvLpKs/OrHjI
R1UD/FBcw/BmcNKZrP7rKf1a/5JREujXYslqouv5xErwg9+bVgcAFx0U1pNdNUIfKcHJIGBGzm9I
dDk0FAhAV2kebSntZVSVsXpPAtDyisZyix5/8WV+kbeAYQZRLX/nJMhCmXDb6Bsg+sHOftxj+XA7
6vmOtzAWlRb86yJM6kSAtQpHqxsT6lHIgORdQMZ/4UfaWV1DVuPNi9zkAnFDupmsXz6hnQvdtStE
zR0y/ipVntVmJXL4bTJ/ax+z65kfpc/S9BfAVX/XpMnTO38vghBEZVEFnOc/BM99cGcQGA3EUYNY
wba257iHc8Bnmd2klQ0KtnQ7NAzVVoqP77TYDbzK4C1COO2sCVNcLZSVVAlWpwJkCj2QGJJhCi5C
FO+dg0xMxqRe0zm+/WVcjC6JYJ9+v13kkwHIvZtAMoUrL0n+0IRose5W+wmrdogaR3Yr+M0v2elQ
URhE2NzzN5zkTXz3XhZdAyVaLrCAaVuy4No94mSerVKwYX6yCvOV7/vnY9hHbPCT8+Zl8xliIwAP
lZDbdz4jNqXbgn+2+Bj7Z1T76NkoOM6norsNpnkrzdqWWrvJx34U4x7GMC7erOgS6W6sL9HC2d9g
HRY/8ONX++oU9Bqfpi+nz+C1XiW5NNZ6QyA8UCTK5Bo16VmayoEIQNdP7sSh1qFznFfQZyahEx8y
wQcNTRQMyrz3JgxdQuCKzDKlBT4vWKYgdvVTsVYNAHsenbY+l00baYSRkUU3Zg8jdkvB76DQ3wH8
UBFvxKpEe+ReQd5OJmp3W6OP1s4L7LmzqdvIitOvvlbbjZCFFDbSkomd8u8Pz097lshyqVq2de2U
0AzCw0hQYkl0Eb96N2tXFEcOMi9xSZqFhKuAtzndDDWIY9WLnLZfAvzKkTpaVe9f6n0BB04kT7ly
anJD/eX5ffjaE5wBrJ5MFsFrVMWk4+kUNGTIyzIhQzzk2ql+4chpj41c7yySI0kp9lVaTqfkXz/V
ArDphfzGAXDADS/Emt2SmQ6GUbFA1BS/256og4EDsdkGpbv1R9NMwjWaaJbovZ9gSxZLgs8tGKXa
8GixOQT6gTSzVwdWOdl3P1ZJPICoAgqM3nXguiM3aYbmAoSIQYGZ9UB6B44Jata5BEangvijEVZY
wtSVpFpYikGTX+z7rc6GkBr8c5GsJf5gZ0MYjffhNdA5dZoJFrjk0K9dafxO53n30dRuUCpBwzER
yBEn08UmxvEUI2jgzVrwxO7aEPR/4qVGSLR8mEL5z7B7on1Fj1cmMXnEm1ktMJ6k/Ox/GeDP+4A3
x2NZmRmg8tZUcIaWUzSeP/JlxCOYmYGQCsoJ1cR+gFhcZ5IcjXzWDcvaayK+ReRhZsFGqg9OV194
nKPnx6QA0vh1DP2NwEfz8osK61P8AwxZrfAcJcejzcrXyRDpximY0xek5AKrnoGf1E45kgqti/8q
R0Z5Zwt3oyySq65r/89GJjDTtbcJY/7SoDejhjOCDnphyRmSnqyVx4b6mk4EBhM2bqbh/9gpeDKM
in2QUF3JSkJvCNb72QVCE4qeFVXBqqGEaK2SWMWNe4qAgE9GK2+PNELyKRC9zTRtfNCXeUvS3jEb
Cqqn3kW+u0hOZ9qeIkD1PGtRZm+jkKTEm0jQugO+PYF81J4xePttepkNalFJ9dY8kdm2vpnMZ/FE
H5abbrMntQBdkgzLEBJNpznlutJUYlmX/LqAqYGTLPNPlIuclUZVx8+L6f+OSE82yEtisZMto3mP
pcbSWHA4C9o4+lVn24MiycUHkzA9EwaRD/LxnC4fORc+OmCgnWUZ3a1s4qfAw6sVY4hQqQDqcFbj
H1U+Z1XS6AoshA1nwd7I6k8Krhk4exhbWsHjAuhKVcdnMxbueR+hmIToPQt5qMBy/BFBMarX8l/k
foatmqhdnJ9/IHUZDDNS3HgvkLcMfhgD1S88Ps4DRsJdCjFHtU/xD3b9AfjaNJyxyjWH6b+J7XCU
5NJpW26W5L5Ow1yV62I9ZSrvMqKq9xnjLBsnkLRbF9bvKVjTKPiSjNPB9U280PZamRiAAcJvPqMi
KnbSEsXYBI+qHtDTPLG3zlabD4dzTwk29v3vkW4Jb81hkRvcwY7ZgywKjHYsROhLt5hZouzP7aFG
axhh/qu0hGzMbHda/QnvGJiBkv9yS9f3llrYkXksM+dALP2As2KEXT3Hy1plnmJrUy/xgsK9+xdx
2ehqpJJn9m9vsbZpt97cdqM25LX5Zb4tgdcZJxGdng3ItrNnmnup7cJSqdi8ns5pby++wPOUGe4Q
kQT2AYzQxZtW3ZajVxk/W2mHcz/T7EYpbVieaSU5C/79k59JktM5siKUBKqx7VH8FFxHjmnZYkKd
8l3jQMG5d27ulzZRGwIsXK0GuQj0zT3cvbl9ujsK4M6OZ1YHKKwlYDJYy8USrViiaQ38pGGg9gcd
i4rA4V52r9+6ZbjE8fQN41GGJwO2KQwf7eXoGSnS49k5Pli3jm+Cf1m4XCSC9brtfG+H592Ejdlv
Z8YglEnM9eIbtkuLqz9sGxVc8+acVh/m8osUDm1DDC0ECLSpJUozfQ2Bhh3JKFO0BL1+jO9PH/Dc
Ku0FHBAhj5wiHgES7kqYZ5f/mMq5eTkfXqRGE9vH/Gd00OpvL0nBkSd5dXvVWnmKtVSG5U0SfhGf
Szj1qbNdvekyqzU0A845XgUthrSl8yWsQPDgNDKxxlvOzP6myWJ5kvSkOlHxlOqgrcMGrKqNk9H6
mZXB0dJdmQXz6a3oDtIIJcHM73TKxg1Sx37ARoGqNd/l0PRgQt8ZeK0Euu7lvhmwN0+37QuLzM//
ytW9+NhqA2xGFG6FdNLlFp21H28m7cnI+x2v77M5GW9ukCEFp/sEH1NoMtYuutONNnRQ/+XOd7vI
03zEtTNb4uJiM/cOcn4GhUIi26+oP0Ur3RJ2hEzW9zFrKU3tb8w4fgWJ9ts1DAeZWRBGW0DliZcM
ambnk5Gj4PhIMO3IQArCcDQHtHHXbUsFH5XGwEbgnatdIz2UxzrW7fTTl2Grl8Z5OqdyaIMPcm9U
YjCYEUDUev7rCjV+ahrr3jyov1qh61nps2s4YOVOKYBs6d6N7xlOZQCIxB0yVOM4T20fgKZRrYBW
8YK1isrQStw1EIedvhYEb2OB3mG044A8MT8X6XXqyxgVWmNWlgo9Pd7gABFUiTGn5tF3n+pTUEO/
mfEiHLbP/2Idzno7F3RoDfR08Fqj2oVCOEgS3znNVdNCWzjOq0sSJEgn6LrdXnFAk+r4FRHHkhmT
zaSQViwEWJwI49xgCk2KbVRm1petvyON1uVC5soZaoxtarirCWKdyYoRWxGPSFWX2/f1avgphpxM
yENydk4/snuMHxnwBeQczELnxphuMpaFlCMhtkICkKsRiiSUQZyfCJdoQ8Ojrv7y2XtdpH33Rz0L
mH+FslaC3O7+fwEkSeHR9P1C3r5qc18eDCd07uuIfivBc/3ePmVlIYMgjCXiiSvs979T312naU5N
Tn+JgaqtlitWAiadgpB/gmvLdEKyGdG/b4bLxyEa13a9i62SzFayToF21YCmRDR9pHfJ9j/WG9XI
VLR0WR11mGuET3QcRW4dJ7jaxVgjcYCnDrTAjQdxTMWZadYQEM3MjpDH+f3yqHoJtYLJ/+RU9f/K
+CkydAl1me26Fqy+sesP9rQlFmlK2/NiwJfCC7DHjeOR+cuU6uhHLwTh0Qa5UXJRdWHTw2YtmE3+
b9UuHWM5OMst7HwVkS0Uqkz8kS6P+pIx87LlBUG5AyMpoLOToLFfqxL/R/ANstWfNECq9uhvsw7L
0f1lfhoTFJeHaIT+SDFFYIsbUeKIO4qmqXubG5CCRq81i9aB+Fek4WW4OItQrG9Y7pvYyD/FnaR8
YFMJ/dm7p/spduV187oei5mX3cy08/pSUfq7ijJkQEnVmQg4Vk3ddeibpIvTbZolp0Jwa8dYt/I2
+3n9fFOC58K+2XGRPXa4hvUbJVXgCziugN8ROjJG3HiWXYN5U2fnxlEgFliDyvQu3MYoI+oALXZ4
B0euGY5bMzOzn23R+rVP/nBVdQMlSkbzx2FIVmfa71t1aMPM/5VXr9+yYlbTCNGRTPJTtyRvjgTn
XbQ48ti0qJwfv4YNxnepovT/CiWD1SgKBgQjBuDVj5nzS7siOMuo5drYA1uA6sf/3KAYsJdQX7fn
JsdgcbldjvhKHp9naRrXI0LtdALKJ3Uy3BVi+WglS7XXmIIp2djaRvnzhnPpp7pIzyMNwxQP3zZd
S0qsA6MgtNYkmeCfhWWcSw9/KCfcyPDvO0OzKmlBU2qr7E8PnWT3OnapmVxrjPT8mcph+uN4bTf0
/RhsZ5oiQP5vbM+KJlwZijQuOeRQCxN+FrNgxk8ykClU+equnrcZwDg1HjN1XdkiaDY7vZGQ/ART
j9T3o48RTzSW2Zl7c3ObUqWAVFm+LIHJg0kCiGo2v3vgJJeXEyHnjO/bcBfKpLZw028WH8lZZg2J
QNh6XL4AUDnnzQBZsgO1XSKgWvjfK8fjgGoYSZn+5n1YzxsX4/zkEEdBkUeMpRAq4esyV7wmgMBh
wZVV0q5CkLTx5pKtT++JjHj3Y5jI7zt4or0jN5OXOXUF/i9PixRwfxGseTyCXYV2CAHCRMJgCktY
Yd+wLmwkQI5rvSNGTM9pUcmRU0hFNFdbYgn16qGP2trYJPKt5t/iJeEhj7VuH2baSgMZs2yWdZmt
+8AYskQ/FNpGJd/4U6o8WO5L4MYXYJlcvDTWSrX9qheN8VE6MbuoEkdgy1mcgPsMBxlKYug82Vfc
tRT4tHYndbCbuj98wTRNnbQzbqNA5ydbdYbflJAG2Gztcx8zM9v09SdOlmy9v4G9YukGH3ljT9wy
HHzyRdeLYNS5Ph0S7jrFrqp34AVaYh0Xg8JyXgvmk/VmVwtmyovlNXko9ba6zdv1qg3o7s6KH2mA
OxmPu/kq99cZBPWn7eFaghTKlmaiDW63wCFHINme/t3+eUErokQjC1TRsi0yYv60BnSO3DkDpzGW
CBbuQTsQnGOFUtpt8Y8pf1Lhi9kFRYtYytpw5YnEzXM2+1CbQiAf8db3OtWN7bUm2Z/rIM6k1Z8J
GaFTDV0fiE9duZawsaLgbhejYl+NQQdvvTC6Qgp70JWG0rR7UZIjQJR7759iJ+3Fhf9HilkbveL3
RVg4GfedeS9oD2RupSvnf02o9rFuX4hj3ZxAj29T5H6odt4z0isTSPUqc1tE7g5TSqLHL1FUqcwB
mpUgDR4xIwFDjanHTpok7ItNGPrgkcld92cI/UAJoVyH6VCw9kmmkbIAE74VksE5+VTwEtJKo0PR
Mhyw+1P8eU0nV/c8cUrVxWkMhOD8qN9K+uryLibNBrCzqFoPuPTmvq1lfr+f1R6Fk8MKcRD9oymu
+rBy1moMQRFqqo7ila9NDy91ex0jhSfNpD2v3C691qQYjzi2udrS1Ycw0qgoyONHOuMHL5dZ7SIz
ydPPrFxQ1DQf6BL+1a3cl4j4DJjTzXh7m3934RY4IRaUNJF53VR8yoz3ZJw5Ri6Q13j8VHuVLDuc
qPMwtmc9X1RroAzwjqpeRy+mvIcGuGSUyqZpKhdoGQ/CWNyf99YmQn/XTw0BRyk55KVbatsssob3
fVsLgjBqd74zjeuwvTuDftaRjU36rtCEXShqIWzv94n3WBKjK49OH8U22hKHgUUqRxjTLUR0rzI3
f9k2b4+tqBZn9ffA8sg19IOQHYXi4sWRraH/mfZ9+luewSNkPDwMTC20wIyviKKU7+aJ0uL9cvQK
JlQooGUsYXjzRhmYUz23/wMFpgM2QpZ0/DgbRdkgT6+q0cTwO4g9Unpu9XDCJWcUJPP8rOhuZ9u1
94FI7ltqE8YKAgA3omvoCYE170pLCYZnzF25HdY48ukqFmjXJZYL9pZV3X+wKk45gp89iicS0zII
/fE3pfB+JF5zjvvElewMqVexM5boDi5D6FQxDlu4XvF0x60iZdgfSvPt2ZasQstA8zid6gZvXur+
wm28GE0gDjK5np/k66epBCnz7IEoAdbZo3YOYrv/nA6SAe+UHVQAWLJTGG2OImXPCsmR4h9t4YEG
qsH7+m3ebN+9LQmpmbdxmBz2ct8BjPpL2qmGGU7Per8LR2OEFd1Ie9TxaYoON9vCHw5er+k7Ygu3
i0lzQ0hzNGlzOVu6QNR3JJNElUUCJqoEM9//T9Y4fK+2tUtFJDmy2idseacDvrU7riq+6XPL8LpI
yQRbtHW1BiDs23Jh0LVtySB5uFbwTaMOD5DBR0cFaUbXIDDvL83QBVQMLrrto8F3zsihf6HU+kLm
FT+RSSQBOygDbeEm5e1BLJHhIMc+BGVEceaqWrQLqzdA2e3/cAmffVIDNfO81aliCeHB7fAf6iqR
3FDp8JAp7uA1lUv3sq9h/VEUHRFanB96DSenrs2wMx30QGC53MZ9jtlplejYeHC9dR+Zr4ihLqd9
hhrcijU1aGE+YlapriMrmeshe+2mm/wZQ7ZMtcpN78aK0eA5nmPaOENknnRrMEOxLxiB8EUP1U+B
k8CS7URBiRiqn7SPfpwGhnwi+IBTGdHqAW8P4Bo8YmZ9yno3Ueo1o0wBB2ugNeQqZP0Vouwl9jJv
Y8X9Onlw+ao5qZKEhhdKJmpdxmXMdksIz5667Hh99BvabQFqa2YayzhV5vIgm0pTi6J06oGs5c7B
LjMlBXw0DJcxjJ15EPYU82zBNOkX1X7MvNBbChibkt7yK6S3CAEde0maA21FCVgJWVMAAyrKzWDr
idGo+v2yyVvzBhJK8+0HvioS3rCOS5hHBlDZLEjXaB3+6rRmw+JKTdXOUHI5dVur5l3i3I0jNJ4t
ttclL8uNDdVrs2xnJrjAwaIxV3SZu8JBSHB+kcBec2RGDFsYArDJtQHq8h0M8Km8bEx8GXS3XoL0
g+O1tEW93cKskZoMtjStHe2KqBLpGio+UF6591nhzi1zdlZr9x+AjJbEUtJ4xszZ91LTnriIlCIB
f8FCi7o9C1YvhGQEp8siCJUW1dS9TUyYA1NgEzY12V7SW2v0EuScRf8K2SqRvL1rOzn9phKdyNmg
DcDD/YuoWUDEfFMaUCh152MoEULb4vYLuJjoYdErZV/h3irmmrMP+RGKoUNA5lR8LzE9OLrY/Zv9
cgGxlzO7fLIiYyPYtkpZfcAhKSSJZR7DFO2JKPl/1DrB6A2dzvql1VDWuAceonXIbrFH7L4HTO9o
fPW7Cop4J22ju7dWTBPSXpQ3iQ4XYUfDXTtwjqKOr2/HqGOz26B2/ABLtWW9QVUMF9KWfjfCUhz6
M1dh6Ljpc8bm3z3L0FHvTROfVmpw9yKKvI58FgoNMURbb/XiQQ9G7qQHDJ0vwwyEe0HDi9wzUUZ5
vaNEZzWic0H13jaN0TrgEewytnDd6JaxrVuDJsnl++c0l9MF3Bm463k1nXQanQea+UZT8kZwgC75
fY/qisi931DBFx3O0W+9HTQ3ZHg+yozkCiShUP5w3brjgR/aPA1RVBVleu6ztLwtHD8k+ta6+rdd
1Ak+Tr+XYjEvn9sL937mlfxoyDB72uW+uam/aMqvjjO4Fvf8xNFw6tXlHOwYXTqQJlpIqiLtTDTs
l0w+JwIwMWP7C9HFNfgLTJZ9+uUWJ4hv9h5KvNUlf4w2mgeWoh237uKh4l7LAmoH0lAWJeje5f1n
LxmS5JIShXVyBRLWPgLDsMh9Rzt2Vec0d/DEFKJ1znGyTtpTrzT8WqeMHVSAUPJ2fzz6FDrqNDdP
VGAj52hq4hvuYZiV//Q8AX5PtEHdBvxLDK3nsZOJigPG8Ano1EKz4wF5HAfq2X2ib8wr8TM2FN+F
UTkADddSBdh23Subbg1fnHlAXkFxVf+0g2qeVgKjwJ9hxgA4R99vw3CsQCi9KCXOolbxOVl+EuOm
7Z5/Sh807jgwUNEOABy+OMG8fxPJGjSW9eD9hj8PpwIvEXB2TmWVpBzVutCWLIJHW8C8TGY1ba6u
qAJ0qU6XsRf2ulAzN1gAypX6OesuM2WtuxAyPVcAZKY0Wj/2CGau57xW7y2OR2HtkLUxjTaHRhU+
1Ux6FI2OJuXnQSHxeKr1PNi2lIv3ri9mEOhL2g53cBjsfV++/EZ0qGwULX9UkgmGVmgbLDPWWujK
ZIATtbqgsLYrxQ5BjyKgd8VOeaz3dWZJcBUHd36duH8kfqkWrbH0jTafiIgmuRTOXbMrKQ9ehFTE
YmCCNFuUmw1sseWlTxn3DiZ1FKsbEv1ZYG+7+edgpyXRqFVpb6a9JT2f2V25gdI2TWXwot2BQ6e2
/tF2xUKP8/tJYeKd+CxjfB/ApWeR70N9DFDEKuA/Z6p1cFZj9DESlyOMWzAVi6vqRPJrxr7IR6Me
hrRM73pRr6Np09pERkvUaOAbo2ZjNvN+FaEWXcr34cDq/iEAIv5LjfEpA6/dxdjEArobTDxEIIxC
peD6RKOj9xO1YsQrp1GFKdFQhQE2XDaL3xlME99+rBLfptziAY66CrIPD/ThcQ52olLhxYF6mHrG
I8G3+c1rzmQlH3U9195Ajw7h1YGn9JBTgtuQyBwRmONu0Q0qwomELrSASLxLHs4jvxmmIW2uR3CP
pl4nUOQ0NBymY+j4uY46ZjFcltlQQX691qNWit0/aqKqRldcYINJYlyMdqmbMTH9Jow/oBiZARC+
pGf5gCNmHrbFj3AWhpueidHX3fP9SzntpzOwcCKqDs61wGcyJWD0KrKQQoh7xhwugHmS5BZ6ZYFI
Oo22fx2MT4cUYHQvbvz6onw8p558XYyn6XdBZ0jsTz9uhMaHdH9MN0gJxfray+D6vuSdP3Z42cRO
qR5OVYNyQBdd/xqwjtWQ4/0szKoZyRF8ms9a/rGIpeuNDXMI4HmpiQ37GhbZr0dnMqxzWEr0qxt5
9PGxhcK3F/rDl5cuc43grUesDUqb7UnHALi3gYSS7I18Kfp5uNTmjXCTmierHaU+M8UueSW9ZkAp
K572xRbxqKMVhQbQmZ4RAsKI0KdAITwD2EiWgkzyCGkP812sq+PPRn7hMlU0KMiRFMXMOmBh5suc
o3gIaXL1wp/ro9xz/OOiisa+wyvLj5tPYd6xtoOrIoDdrfkYpDTRrvkwIUQRFAnP5dJK8NfDvzhi
6scid8Aba2Va3Di3KrefOd3v12RAZ5VegePcrXOuBgpeiJdY8HwCaK3J+dMrB7oaESsxAyXMIy4n
xvkj/TBiBlSw40rw1sDcG7F0TAqJ0fVQgLVUtshxveTWf0Lgt/nRroCUVE7D+gZqN2DT4nMija/t
OxZvNDbxJl7+mTSJtXb2dXEE2StGchUXnEoyPGRYUU9dSaAIFW6u95BOFgKIhxi5+N5VfmNoglHW
D2cqLQno9DyaVLRSS+7BFgTL0AQ4eDEpjgKJgoEhOle62HaFvUU4a8knfkY8yTsRSmBFx+auQxbE
txyu31FZd5MglUJNW5qjeCHhkhkufvTErrencOqg7forSCYvHn6VZwpnVE+qrKfvXwF06+wBlEJ0
24cydaz/xO5yvDJO44JEmk3zbjQmKcS9hjBnjxNaUOeNK5V5UGqAHhJEZwCcJeMnty7BeRSU3azD
j7BdIVpt3E/DoK8nJYPXO5yeVZD4aQnzjKL0yoX4vQ9++L+GOkMA5ZKaEUM9++ab73JJlL4QG1l5
8tsCe/IAlMCeQsbm7HgyFzTjSNyLc1J81tlLs1B6GAKADCNtpZ7xCRt/lvvKRiahkJ8IAF6+SfdX
yKmh638UgNy2G+9PraNtI+dTSeVL7LYN1/xlRfeYgR0J1PDC2q0PsizSttZmgDieIuuqOUpQDVtY
PZ+gH8ZinYUx7k7HXSven10VokqycQZCVWcCpgPDfu0Lc/0uZ8Pao4uUwykprjJ2qoHuwHuBhO00
5wFExP+cMh+e190A89Oyh2ksxJlKbZro0obxmInjhVuhY/6uL8C9ancDzRjdHXxxrLwAReYA9WNX
Tcz1wQ6lMXSnhQMZkrW37I5yRrC5e2XUQ8Z2Ac2abfQIfuYLZ9iuGUJxWzrciiPBLfqMEGCwRoRU
N3JG/9MEqvTlOuV3jo6AmMSY5YZaribuD4ExNm5W2/XxM3TGNYg7aemW5/4if2yRruXOXKWFrkIV
fPE1BzKYXsXxWvEpioYU+5OA8q2BTCu2Ng5fdfHYmI48a89KioRwKF4jD/7+jYY5Q1oHSrFvEZwQ
2LSUVanJJzwa/QOzvY4/yW1yNfMs7/VctaDoB2bqMLRABDBN3ByqyRKmRcHKROw7kwF/ExorQQZY
URn/SWchkZGOtIjO5PyzRF6UbEUJd5mXsa5pHN4/nyHq8KMzc774OF7XYNpMu16Xk3mlzJm9kTW3
IajGRzvS6JMykHIRJqYOSDcjZM59nDMOdKdaLd1Y1F5pD7h2TpfBSNfiwEsbAujfg/ea8PkhKW+D
T8HLQSUsXEaJz3UcW7i4tm/eOeYv0BrOHtgUOEs3foQhBGJ54N4UGLDBDp9IhzjA+/Tb9NIpE26a
IMs8X7cNpGlkC7C+Z5SYEv3QeoQbsVYhrVwdNnEZYCjUj4Yw5cURbznj85p/C1faX0cpud9uUqRz
YifY8CCVvqJ9QYXyrYlS1IZEfPzhPMPBmWbGyGaqeuaLB8c82tK3XC9UECODSbQAIlb0fMQAntQR
Tv/DLExyLtAjyP+ygo22BeDjnOCIQc4t8q7WWJgAHXlSgIQ3Hl8qZmOlbaz63xm6FYHY2wktUjE1
1zDoZofSbQaGm7i4Ss9bqS/21Edn9Oc0Kjr++DZQytVlBE60JR5xjQOqL/oaKjUuCTmNdNTuAHdS
VfAzZNkrvv/iq+MSKKIFanTFqJuRuXCeXrn/IP746ro9X8X3p6JNW4dLBGMzlwhzMlFruCHvNJv4
lvateXTYkp+If/eH2dwWNTjf/P0tF8re68Xqd/aMF0aadGE1A/KwqVJfrqiSEVo9mOSWo7B0Z5py
gViTiSreDgb9TnNtGFEQThcy5BFcLCkvRCR9KbFzyqRtYrJVJCLqRamx8B+vh500jeFrV2+E5O3M
ksBQmMI9oh/Rqa313H2vHVGzp7iyX7ZRd1YPQMylz5SWYZCBzgWz+HiYy7UQq7zzsANBk7cxzdcO
zGJA4WMcwWy/q1mScjKdSZALksDzqKrY+jT/nLoUNs7BZ4tcUNW8Pk1exmkQwX1AfWt4z9M7u04b
xXQI75Yex9E44Mf3RXHjShEcSYLKd+UoU6RjjtLH4V4uislfnkz44YA0r9RW0OiY+FMUU+MDJ3LL
0TBoGObJqQZFh/W0AXEi4o52jlrFViU2V1SdaOUvfATkzggUnHYsKevqZpWN99jwQlYb1g3JV3nU
+hhf9VDunbpLZ73cjGCpQLdIZF9FKqSxKM7oJco0NlWb9TFzAWOwlmAVkFhgp3ysU3oNMPDQgp7P
mCzxSkwdISfmnkcUoVyoLoXfDtLttNZ4Fow3LQBeH9Cw7CWtVtPdRraGZAXpj07xiytatWSO2mWu
r+g1HrVGuXobUQcNsEN7UcNssPyPl7vA8DYaFgMx/0hBRLpZ58AAGkKsFgkwnGXGpR7nSl3lPYtj
Pu+vkqx+kabS+Z84sx4pJg6LBy+2Sxx4LuSw52w5aIQuNZFenTlGhzvIAvuIlcRq0pClO5ec57bK
F4AxPBmYj9F6fUGCUUaWhobAZpVsFxxV515yHbQbWQIbBxjM631o55P32qob8Cbs2t6zUxhzCZ0F
Jm0W1fM08QOoxmThRrTCOdxRxbAlCybv/wXu7Pq4iblOObgqRsblWiWdYqcgVi7DqgdOEIUrsoY0
tyMZNwXfZ34VA8gET4WYDlMfimWv/lm0mGTrjTgPB5yBaxCHhCY1yn1u/wwSTNsd0oZSCaYoL+xQ
JKX2FR+1w7zdyUvEek+RxaYZH2S6DhJeBTXHa0OJkfodSIu15ZJWYg5RS+0z1vCaSSNTx5Y8CnGR
CG2X9vaxBFz8qabN1VDCWL7A8Bcb6ZrMr239vsD4BgipZsDp4zF5jwkVkDwRGGV6K4sOaq+TqSnZ
Tx4A8JpOb3zleOAhFTFJJrTFsrSHWNAMr+KBeaNrBiFyipCRKkUgeld4ZiMQ8XF4ss38wuPbGR5p
injlyt2awImXx6Pj6tz9KFbNIuvgEu0c/GYb9p30r9QOvnfc4BrLiow+D5te7kPCGztpg6cT7OGt
KVY4RdSOLAlLzKbNv6TAGoJIuo9jirrbbX1WRQdbZwhzLnjNGU0ZwqzpoA+7UdzugIhXkWt59VTp
vmYr8rPRhzQyPvxvpoUFNOFLyjm/MU4MPnVK8tqtY5podvBEHAu4o4rsdWXIUMmUJXsLHNZpBIV7
CgMFtcVT6xO18Rs0qqGm1gEYqGeXFSmg/zMugOB0vXx6oF4b6gwhtdSbvkE1fC8bUheCgGDw7CL4
fedRIxzX179xFzPGNr/P8pRG2Lyhl6ngB251yYeZ8yPoAaxouCylXdFWuNG9p9o8p3o4vqMh5NMH
TDxSkSfc0LUXeyBmPf9p95s4+CLz4vEels3aZM8ub88PS7XZC+iBm8AZbCA3n7k7pFUSE6Tk9mKi
Nwo2zv5Q6kQhAl97ucpMtdDcrPQ5YtWCREj+qUnYSMNHdQhcdaDAty2uRdTMWlf6A2rTyNVUuENZ
GzGTmQCcmwnWBNTdXKQofkz2WeoJDiIxPm7T+dUoG4OfjQhv+90E28S9AsRk6tWq2FQ5615YwKTC
Cjz2k522Qz5rtP5YVhQ6w36hQgdQFNEwgM5b8bQkaLcePi8c5USGtyFEFHvULPqW7LoB9CUJYcKf
O6TAr0CF3ly8ASFH39kKqspv2TFfU4zlQ40K9Rs8Ru630dITJP1NLJKO6kDV+0z2q4aSUEG9XBrx
53xG7qglUFOZ+1kThxm9m8KLgbftthTcuSME/SS/K7q2kTG9tsxyK7K9j3znsZb4VKy1vcvadPNu
liizGHkpuXdt/nFdQcfYNFPI3DiToDNR65rWGuI2h2TonCx6WPGGqf9IJ+OHwruNs+Zt0A9raT4g
KWv4neDR0w1/VIPiNbUwADzmmfQN8BbA/FDw5VCJpmL2yMfWVh/e/SsgBOIltgoAZXSBUf/iucr0
9z9skUvM6kwdorlTDQp9LrMJ19SwKXHJNxSFHsrcgkAzToINS139hYpWFuaC7s18kF7h/YXux50i
2xsB04+/I6us8uiMH66nGPGTiGPl/44UDOlaCtMtax54CwiFLsc7CRUbbAYkivaJ8VILcspIG7An
7rQzNmdbr3BY+1nRLNAUOv/WMFjqtLBrw5JUNbp99Dwc8ozYcJawJE6dCmRQLmEzZdJH37Sv0LSG
bFbSZeahaLO9rbsnMjh6NMRiVQSKxO3I/j7SO4Nym9lyB9jkE8ZGIeNK/VqM5PHik8feNLqEj7X2
cFQVwKtH8Nbx3SR+PedwMZTIo2rZaET2JwYHvPvVHcpLGOvSfYfx+5GKKjq71siaETWKomjeuAYw
BkIe2HPzQgjGbBSKgmqLWrAHCgWH8FT1WQ60dxtb5pfsg81Ml6zQMwELyyt7W1wylcNlEjY36yb9
nB1ItC6SQl408CxnkHWPq3k7Cu1NfYWle4DgCX3S95OOiHz80BOOVxNS3sQRM8siAB6chU2ubgHS
QC6v4paBUbkykjCCe5Sa9Qr1zQS6ZIh1wSfY0gBbSzCc0KlOhKjZTVDZ3xDbIsLaLMD6dURt4gs2
5l53T5fVHKcXS4ZGljEC5vpan2lMKqpd3m5OMgZyZrq9Hc13DWr559FOi9uCOyOgvxcUwF9I81ka
TGHr3kJuNCfCGJ823UNfyk/xUvVUfNsRfQrvojke1p8woSGxDRIZg2EaEtENlSkAL+Y5clh38x1w
BZqTz+skeM2dKbacIGHMH/0BaJE/0AZSAyr+dM78CBAy5i25xDs3kBdMPvui7j9nRGmdCsdqcEsa
J/tBDPy+tertOnR9FKf7g4q44qQCUdUdncbbkeit7OHnUFEE6OU/5hlNioeFxx6mSd87v9pU0j1x
BO2+PY41oHxR7v/iUz/HuxbJnLmk39pooMjeRQbHnq3XeVJCtA6JKR3lkQQKtPpvZa6I6i2+Xk1I
pTUE7sl9dZtKxUgFlilGQGQn4xtgHhw2PijF1pSTky0J7PbHcZtRQ3ALCkoadMlQtgYWNrxYUzth
eBwp/+IkSFL/Ue1NtFPMaNrKt5+fUeC5nu2LcvaAV2Z4yUcfErbtmpcTKUsNcynIBrvF2+IeMmuS
7woFOv8pNloLg71lWjvE9U6CUi6kNvOrkxMl2MYdTtw/cNZ1hHMgj1JRIIzxAxRVrF6B7uue+G5Z
3vW1y0x7wXdOPn7h1HR4DZxfGOT+ExYPHSpcitrHTMDxjgM4+puth6+KFFn5IU6QcQPhYY5gNKpD
7b4ieC8AITkTPGA3rY6mIXYdEhq0AOZUXvKpvlcZMHdISgK6mjFKrjOvi1sEuD523szH86JyNShI
/Sj/YV5YVYH0r28nQHeFGPKvxYq7l9m9ntgYRz0C+nEmvgC5v6og5CqaQijo+qwo9AAvsrodSYrx
7ZhZf0jXvZoO9hH0BFwe6a3WbGC4k3lwkKOuEMwZn9paIkoDM1aJsvZ6UHGtKa5RVF9iTqKFx7yN
ZMQEtuSo1Lmyf3s1ZCM4YFuLHEmStT7IiOThUIKxuebgEL2xpXt+DCFhCuTdJpSM7ikcV83TdA5T
eVqmFDJYLPgNRbVikVwOxbJAUxtdyWWQe4FBMLq/c3Qu1kVx7nRH51zaUm9f2bV2Jb5m1bbLHkPw
lsV5yzhB15FhANwhxAoc4GmExL8RWVtqVMbP9KAD9dXsn6Y7xk0Y+AFTZiY+VB4/x74OwypWRUwG
/nEOGugl49k8Xis8VXdFQw8oxDpoHJSVBEkRy2uYZfw24vmhK2YXBhP2sAGOeXHH3mP9Mi2Ekk8O
n62LK4Qvl0IgtQxosUk/IQeAIba85hZBtwV/H/QGHkczAdlwpnLJGBVzr423HZQDx+ICOV0LlQ9g
O43GkVhypX8Y2xJCaRlWYCPUhXTPAFpMZN4oGgD167r7/jiyUlOdnVdVbKDHETCS/m4v7Yi/LjSR
zs6m4Adza26vrFuGir45CYJusuBl1Fqg0HfIoM69kdGS4/wfJGMtDpkwsUuFssTZ+IuPCnSfeQTC
DZcg/OEcT14jZxEogv7cfk48aWvADhCJEgqg4HdRZs4n4CWe996YZyvOfosq/cK+awOmcJ57bzy7
mYZLd9rk4yX2nxCECU942DZ7ERCk2XWOcJjqDWnY3SUGDZ9gNf+nsqMXG0zx5QVaosbMFlEMZ7eU
WJkXL9L27FN20e8wLt2kZwQ2a+th3isbp2DBESS2ma6iFeiOlQICBGKRkiiCgF6OlRfNI4kLrQPk
5Z1mlzEp/6x4ktWcuRCSxzJ2Kz/8CSEockUpXvn7sbx+/gx4CtZ3X6KQLhGl5+sW5u7gc2NSB7RX
RihZ4KV9VyatxYexKqvPjMHdmALnwdtoesZYS2yKjh7+YTeMCKZIdt1mSpzaZ6vTa3PwSGdP+wqg
GjKMCxKe0+KGLNdWrEUP7JtBld4BDl79VHh8W6Jdz13gyuBRcje1mY4/5Rc9c/duy3cozvA8hC4f
RE0qmgyyhPurrHfnAg170vn+WSrQIHip6uxo71zqe+yBzGXt6yJ3XubtZa6rhMU0hhga4/SG4edg
p58GziNPnepLtcMJCQvWoddVzi3yO2mc+zotByBU2otwF/bZxotOPEfnKKCXdkEsyitzuATyMBmi
1dnQ3CLncs/qGESreuuGXD9kbB4X97DlR/5L1UvcHvKfSHeEOycL38VP+3AzU4/u7y3Z4LJdCesD
EL8+ENO31CVEjlY3jtAlBD1VHSxNie1G/WBdpCr2jyr5feJYiawxg5twVqxuuzxHL/y7lXxNHgRj
riSYXD9n6oIZGS+P7skvAedF0b3ySeiGXb/B9UEJltDa2ApaViOKdhupIlwpK6Iv50z2AKlmHwua
0IdFof5ZCzMGpaDvvCI6xUDqeulkWIZnFlnISHPcdhJspHLVL58L7en5oV/ZycDihjdYsN8fmNwE
NuglCQ+KsYnR09bO0+RsImjJyOg99q0oHuiZ3nkbaAbu1Hsvg2d7D4XMoOd+sJlL3Fm3CxyyVDSS
xKWRWQgS/suLZc2Pq+0xkBXS1/SYDOyeYFNzYGnPEbt8gzXmIhKu+BKBCjwflr5magzjAVV7Eh8P
b7CmKWWZnjJGcfPQ3dqYSg3CezS0M1Igq8qx3TEUc5junTvm6jxBLRCyE0shKyWrmGaXdyrkwN0O
5ZAlXhfqxumvrM29vE9A2veOyNpr5Rb4UG3NepgQmpczIDDCz+6hQ3fzj/Ns6iEeNArg0HByg3M7
+KIJiTEizJf6QnVD42DuIizzAQclAPXbez7Fqn1cMFjH/PWuMH6b6A3ofq1TCbmlz++ppwFpJnxC
yb1f16tYU4pK4uCQRvm09+TyuDmtizoYVZK6OqapH8vFP+8eiCiqneMiIqps/mhx59loF1W0xfiI
ktQSj9nDUTvD/kePdfoSX/P5UW+3+Es5i4bciZ6be8mZuvS70T2Bnos08sIlRWpgiaIOTx5UGJHn
3u8eJjiK4khue1JhbMJR7uIRldVsoSYia1YCXAS0Hab3vLSOkaVi2OcwiJzgvDybRoaCW1pBGPjB
yo4ThxCM9sW0zFYusaYVJgyXCqz9N3hHmatIJTGomuGCVsoiMjUuDUbqysxiSOCiy78SC567fDOw
TlrmNR00x3c35bAzAzMKJEUhnLs+awxemSK8lIIP/QyBULnPBelmyaZXmVgUvdKNDQSx+NAfqURt
2YRYr4OeNdID3mddj7U00N5pfALjrx/lXSopj+2S2z5aru5HUWcKIBbxJ3BY+xh663CSzZEs65mi
l0+yYhkHpjzQK8wjyjfew+5XKneqXLmbIzY6l7kdJofe/dJIAnrbd6NHr92P9wfir8fgxqZSWBN5
x+EiAssjH/ZI8bdw17mba7FnF5n3FzWrbAatLM6kCCo18ADopArBQIrmqrkHdLTQUlogo48pnqo/
a3I0OUVDlBmMo0AYatJaU4Io/1mHymZ5XWUoh358coUI386/0HEtxG1LSQCzhVdzNcZA1BJurche
hM5ibZe94CkawkubrohUVpITkqvj+dOOLK0L2VtVspMizTQKkddZezRo6YhJHTx3UnRCP67WQTpE
iEmGYuBTUBhf8Xq7IQKrZ+7wwooToKouh63BZVisOjln7iiaa0v4e5hrp9iAI5aPfMewAy8jDKPV
FitDZNFTx3JqXvCuMEwaUCmfHM8W/gtPP6A3Oa8BphMxbcEBd8w7X9ipZbAiqGo+ZBEzJFXErINu
WSRzxsJDyM6xCdvrwD/n3bBnUbJSf9SaDpEV5w85gGasgG5RqMNYVUz0yICxL5vjFrBnPyhHs28c
ioL6Rp/xnxH55pfyupAyux1auabWIm9fNfnXmd1PXf1ffwS1zfjHCsRgM13Mn3JIx0zoz701OHfA
biIahHzg/qWimR/buw11XWvdpscKXnWorhnUMi2kRYesfOQq04XX7QneWVOBulTHhI0gMBByLX+U
lK6lVk5DT+BN0AVpIZq/iYVCgLxqQmENBZeVB/dHPDlVbymgRYqDrLWkVQ5VqPjwDNAvDt3SEYWq
AYLCLZQ0aMPOVfmkC8eCezTm9w6o344xDIxZuHOiTEYZH+Uf0HM5papNEJBORIqV21LKWx+93II2
Y/OQHXhgY3dbyuuMbs4KGjB45UMF3H5CDzxqsFqQMSRB40qI7L1LMZO9/DTW2N4IKgeMzkFZ6k+Q
wcwWfKzZUGq58mWdDRsVqvK+7/jy9f7sqJs4JxFIlu4WrNzFV2qA4caneJAljyv4dTw4ac6+kSp5
GXjxRcFWWD6qssb2/HWpiXABh0slLOs3Mf/9DFpABSZEGWtrUnBGJuf4cppllO5QuNwXxtvJQtEW
/SlZYf9bfty8vHL81WHr+X6ipHNWlz2gaEDtR6LCukjTWikFT2toeX4Yp7ka+mAzpdjQtpGo1qld
S4K/uY3c99D9sekzkE5oec1UFG7aKuZZNsgcPT12kk4BEXQt62J6BJZ9WJTRvOUrpMITmqfJsD4w
MkYmEe0/RkEMF7kS107IZw8d5bPJYUWb5RAUQv+lLEdX+Zpd8XAKm8y9bExEiivEFPovcr+x0jXh
NUzRszON/h28EfzekI27MBGeK3/dreVUBWWrHyhOAHd70qWHzADxXzdabTZMXRX5fpWaBh/LQLx9
HLnkUPWGIhmPOPwYSomK4N64rE8wxue9mZLFEmIXsEjskbdyklADq/08Er2aUsKlBnN/Pxt1hQhH
zt+qzDbQV91OnUrP11lQuVd7qRCJawkzgKHrspTSYmz1aa8uF4So8yB0a4Gbl+jwf/kgy22BVPHt
ECDBWovbS5XsTytc/B+3YiusyQHClNyMDtbsG9awqi1vrnK+6kxiuRwaNR6e6WVYReS4Ck06WG1h
skNweIWlnb0Utiymu28ailweMPD3eF2VYHz7sJHBWK2JEF6b/8iiv1mPzuD/lFzm2Mo1bbtQwRKY
xBemjukmBtdYEStbFA/lOulr0pG340uelAxq6tnFDeerRrAPAj7d5dNXOyEknV33zCcokKTNRi3h
sQZWi74zwbTKG1i9P+Lw6KW9ilG7YaodIKTRjmbV0mHoIImmnBw5smnkPs53gIRJHAn2ghxry3qy
dp+dzWjg+TUGxBCdDKoj8NnK9bN9j/vrcWspa1dOhyJ+PfaVCpPRcwH8x6oAJ1M07/fYjlkHLZf0
YQDuZJvisAuQFDAYu6drpeh1SF6zAbQVmufiGeQb4/2CacI2y05PrArOrtmDPOTPutkSuUKxCtts
/CmyKSNfRPVeOsEbUCJBn0zUCur5ngIsRz1Ddi835jQJ+TOs72iTfEJgXfgZF0XS1wSNjxc1pbIx
+y5rNuEkIWfYih/IOX0mctkmA6AvvoTbF69uc3vAdW0MxwNR2W+sd5i0pWi+f60p+jTueCPgRwQ3
BR7guEfQw74lWNsKOcg4Ls05sktIjwMIK2VfSpCfSdy7BH6VB7PmWRR0VGn6FUHAsMiAZSBvZZCu
Ung6yJgfC4mx1XWnyDMG2lNpsquDeg0ee6WmOCCRne3qzw5IjwGA5BU8D9ImLTOBuZqlei6E5bZe
xZ7f77f/90/HlfAYQPhadraEc/VgZUDBU8f6NQLW3Dg5Vj5UlUXUhqW3NXY68JLuiN4K5DiQgVD7
Kbna0Pie7bB+Cew1b9NohtKxmgPbevx3gOaLrAa1RN5kUW6voX1F/T12/koSmLOIXq2jDkdDAEiR
WHCcH9YCwdkDIqoR+7I/+rgeiC8I/30PSgRqeXYOpQ/wNQpEtx2EtYa5Jy7T2WpBeA+KRClK9V8M
nFUr12MVy/dhTHTf0s93MfyCgWo6cq1aA/fFyvW4WxeHamXgVMnrBlqlC9poAp8qFOgVmtqSyG43
6ieD1q0H6RTzxM+Ae4IqOozqpRIv9vf205oY/XItmtvEvTxdbVD3YNS2BmZPOM4JNeXzP+7rRTCH
9oc6HkIyEf42Z7km6ftD+dN5IC3RxJ2QeEf6p9TYbOmmfRBJ8SX8rJWfomVC9JbFVpuKSt0JF2p0
YiRCdtkVogPyiXhkRr0Du5cQrwFqa+ZUc30DRq71A/1DOpKZy+XlQQNNXEaYC86eaaohyRckP/i8
avwFzj1HTdhGQOd7qAjNSFoThgQ/vKH1auc9WKA4eK9n/M3Mi7EZu8Po8mRMUKZF+lVHU+0QtcEB
Dk6Rvj8HKJj3Qj5H4dB+qVOzC2ZK/T55KL5r5a+ryyE/6Shyrq5u8jLC/2horUwSZS/h3CMbSjIb
WaH2AFFWBhdR4BFhK6n4ix+6vzwlJEaBjGNlOkFgcKOYd0U8meJWbZ2OJkPA6Uy8ubU9REY0DDDw
nE0SiuLeHYK9LNwMmqpEjEqkZo0Jtnnv7D6sPNYx9VWAvA+VCatgORSRyGBkIEKvCyum6QdF3sdE
6yjLb0T+gPQDH28P9ZYXPdN7EC47LrYBk4HVNzR2dnTmzDQjtASwTzTdtZPFgtcJnumCMuqA/FKb
iZNd6ZUvzFOJUubZf5r1+HPInJtzqDaPgzPoCy6UVnS5hqs1DHsVfe4jdtxraLTa+IiHGa5p351t
jRLgOcDD9eV7U9F5Mn+DUaHQEjsPNdexSzuz34HcKGHnaujymWRnno9OW4ux7HgymNM+FYDi00NA
SuPV3gvHDVUAyiAUKhZIxiRJCHdwf+IPNW27v6q/bOVIidk9/o8GEDpLHrX75kmW0P0ssFDY45fn
r+Hd3sWhlHgGWzftbQYerIu9W2y8zSYCFBTDTTg8vKNBC7QVfbTiRnA2sx0pqIiI1uB/FAqaG+XG
HXODjkSz55kTbVZUZQLRgyhF4bKgODSq9EqWQGCNt2wFp5naADHr9+3ryP4yC1v4DWXKzO9jIdL7
6Qgt88GGAhqdRwZFJLLjNt/4FCLxLB5UR83ffGqTebGHDxM7YF/fYrg9d6fcSo2IllfHEJxAzlUu
cs8/ZBWtA8MBg5iLzkaCZPUn4vdEqq4FhnMKfF7gzG9JYixPxZBdSk3qTsJWxZwFPY1gMi3szBKh
iBm6bbHtAMa9yFp1Bu0TC3ipfDwe7BGP9+qBuhRuhaM/LlltScQQaAVWMEy9urBWeh0/7FDao30E
KRSjbCGo23sCviZ+GbgZr5boyEc2OxI7pbeBklwbODNnU2uyKf2qaA0HR1EcZXsbGo8/0mjM9+LF
rdi6OtaTL8Bo5jUM2Cg9nizoU9M4Tz/pLd5I3TrNh7VnMqhoqjSxl+YfgMYtQIyDjm2+ngTgW42e
TOFNwLJChLJGaI5AvxTTD14IXIJPBgsm0BGrVFli9eeTaTRCy4iLTfA4nxA74Bf2AmOJAmGvifpH
C9BpjHgk+qZpLj8LJ08zpF3l592WyIDmJ73ylLxDQ6700mHrQ2xUcWx7C39kWyfAFjL9zvvIJYJn
MmtI4FZTQ6E/SaS0gCrZjH4WXl0pU2ZcdIOYtaUOHKI1gySfriqlXcnj2q4NUn+8FE4fpN018oMp
m56GuHpqkszq401RM5muz1fOYVOwia+4IYribai7Ax11W/0+ZWKqPYcM2kpYc+xz4AMNbSCcmhlq
Hk9y5VXgSRhGPAlC+veDbZOUHvhvhoKbS3bgdGQy3yCaqE9j45mNjFwJCJUuY/jxa9e2ce0Ajfph
foZPL4sgLTGkXqd4t0//I5rsPEuEzuytg79olPH2yu1n3pLqPzJEhfhAOb51EUtcXVn0A2VncgNy
B2AXbvNhRANteq2HjdL44i56oAZWgTZeqZC1/VdWYsCwK0kAnnUc2GoIpcw8hy14l9fy0KJwny9F
ZHQcSWENXZswzEDHHY5oueqcDaaIUUq+x5bJP26MIgy4ktwDvTJjT8sbNVx3FvV94r1r6FwoaKSu
YXtjoxNE4rvMIrtB7lH3WRtbve6Wlrm9Gui0l6Plck2l5fkQ1nOVF5Uw19DgvCz/G03BznnxirF7
6lslWwnIHFrw84wPwjDZA3k+5gulhT3AGfArmq05BKuD3JMPVFi+WC/UmAtthV2OhRH58toM1PVO
HNeXll2Ok3gXfZb3YAdQ2E5OPKTI9chzUSc7I8YOsUT8mZRQriZEf+dEx4A7cxufAX/6XqF2QSZg
+DqTzgzpm4aCkdGtH253BAo6waF5DLMW2ifZ5Btii93cE64GqNjbsQS5yfaskFDXA+ry48epntY0
ZbB9rL4CVh0lvFmqXPRo57z+HuHGQg6xc9fWXhPixkDnZBqP7HuBBjgXUfli/ScH+uKrwaATvnlq
SJ709hrp4bzWnZG/20/sXkHOLUONkMueqfE9p8Ggf+Ki6pNWo/QCUxtZOsvxAIqMcLRV8Xeqn26c
8+2jhQmsYoEQwZxL6hsFeJaJqEbohdygaCJisRpEveDSmpREE1boCoTgYFsBWdcI+zU4OpTLHqGE
6vnhDpyiyOTdfDe9n7d/RgYLAY50EGh8HrJSVsIqFNp7tO/o6pONZRi0r0Moi7HYSJ2g/Zr84mCi
5EQTWfpvBS4+pkp1UkelGotEaHdcY20PpYgPXfTr+7LsIda+6b6382jXDYmwp6qM/SmmHQk4Fgfm
U0d7ZTwB6HSHND+zAoqHNgrjubuk+q68kMsEJ085NIGkUY7woHyoNhNIuEvQHinLCEdSNYv64r2J
A3ZeMS7s/ZVfEUlpB6/D1Fn5U3fL0gx/LOIWaEDNanRD+KDqbpd3aZLh2TcwfSHolyVu/ToMhYe5
avDAmlLFJbJjsMjRUjwF7wsFWpOzKcYajMmUu56NZVQTbeL5YQf5uL+qYGYnQvDcnrkCklb71ji7
RUCVn8uTm4fMyTMWPmQUXFzgBKYid1U4y62yc7pWupcjFDzoZay+uP/KbfbqFoEnTsbCBxWizmkV
aV3DrhSRAPGZj/doVs4+3aGCpeDojWav1kG5wFBRIYYOnirtHjgDD5On/JvkuN/4YUkdiJAHFE14
C1O56FkTnmEy4UCzrYjJT2Ug9gXScN6bjKaBOObI8zk6bwhLKC7Von6VZmiaP2m86XvrC2WWmV9z
V+7e9luPu301VSIqOHQrtT4TP2OQ/UXdudFFWtdC5VOmFUpCvt8qCeZ5IeOm/Siwls9nNtDXLWKH
Na3UrDzTkJJfeye7yfP3QfH+JlsAEJGwOY0qj9nvqnNK6T0Ml/TV4NTE82E76mCZMpD52T2yvMn/
UYAKszEE48JQmrr0srZ9VS+xiyf9cufue91boWhRq+4185fuRhwQs7WxJ4zgJmOHA6gj9kUqKpn6
X2mT+gP5sZuMsqAirPL4iPUmGfj2s+dC2OxSBDXJUbHKsLe0qsd7/li5Dol1+kptqtLz5ZK3Q4uZ
qUK+JIcBCrzT7KQsU429sJUaN2GPeRPey74oNZz7ADrT+hoNb1ltWcgKayCXKNQM5Tkpv5aaJ+Q1
jkNkxcTMjKu8UBSwN4/s7/dIYphGO82oI+HK5iNyuPWuBn90x4phExhsH4J7VQl/XRxZsyepyJ0t
FUUcfOOLy7xWba1jqS6lE8eays6idLtBrLIR4T7b5hFTzpd5y5YG5QHFcKecBsBw7WzjlEhDi8ip
faq30HkxPEKTmn8zOns65Tc1btwOZGzeQhTdeDELd4/abu2EQBVuuAsvbCC0g6Ot0Q5aByIMB3Ey
wyiNU5pJfnOWWRF8zTTJUE0stGjkWEpWMw/gTkS3Oa+7FB/4vd3Nv7kx5RWFz0tMHecf4ZrJkQlM
P+UuQX0eUZI1q4cqEWMmMGwvQqo0YheOM+LwCBLuH2mE1GzaP0m5CVD2mUY1VxfxoSQFclR+BMj0
BModR9haeITtV0RCdSrr6/2jE/D/IBCNutuDxcHGEdExEcmy4BW8WTukyHgaQEy4jbj5pDrGa0fl
bDbOnaBlB35hfU8qLiX5jGTvcq8fQtnOpjFpTKt8fEXJ6ZgZZvGgOQO0TvRQEQvKuhyw4cQflM+R
3XR3TZl7QTuh7/JJAoRK28O9Vn9k6keoAQpi2Glqc0G+urct+l8V0QMLRQYX4YJWzI4eikmNnuYp
DJ+LrsY9WbTlA/c0sTDB6m3vy6W1pFfV4RxMyrD3sVAg/po9o3EcFY+RWgyvkxfuaW1JGBP2HlrH
fis/VwCsGeFKVUbfRAHpi5YoGDkNSWFhOQmVoyd1otat1+dmlygmDj2T+HxA0lP+VknOzg0l+DLI
N3hkbju+RA27XKoeVb0hAhTInWoAQph8F0QpOgO6E7cCWFO/1XE4xdtXhSF4KM06Hd9jPjhHdbfS
6wFa6a5n5Fkv0cZ3ZRCh9f0f6+bdHNlZFBz7uFu5xBqLJejEB4UjBJecq2LwuxEebVU0j2V/70Vb
zdA1lW2+/uzg621To5ysxKtlK++90x/JmDuH00sqImtGF9JrEL0o4ZvijSb45Fv/RYsuT0DSEr0T
lbohRTiLp0pMubI53hwIYSlou9f51I+85HoZvtqTu50KxT5OfNgmDuF+E0SF27NxTsL4ezpoicVg
B30MofXSI75+mOsEtUsqPMsZiZDVF8Le8q7l5okAisEoBHVGoEcRmwXXr7OhG1cQ2+X1ZxFI+f8g
CavYFjlKFSSf3ScAljLhBxgj23yiH/nrOaZtyr1qffFMrtXwuq9UK42bRbQ1HvtrPOGPU5etXNLO
30MTo/zlJJQTNEXAeXdPa7V5S7F1JIrWCG/BZ1C9mktK2nr78yslzG04VaMbFyPxgEsvFH1r7d29
rCg6rYTzTDJjKzdoZiKybqW2vEefI/7Hm3B9Y/EcO0X7sRcQSKDlruzPTf8jDd94pR50XQY9d5O9
XDA1SvI3eWkKrzSfLXN5OIvZFVXaACpP+OoDyZ7HHfN68XoWFoGj91b42fsWFVDZpN919uKWFC2J
JVEZqTGy52TPf1WSdFdtjinaJZB+4f1CTugJ8vA7kI2SAB0DdyTdtDrKubkzoFeFqle/mR+DGAwI
uIxCTODlXk988eu0vRKXzavPPIw5aghqR0vWwB6e01YGvc1L12M7iOPQxFY5HW6qYnr1QBb3t5B4
ian/W3BG9GG+h3j1J6VZ5FjIIjBZdA+EteI8suPlRif14myWHXvPAkpfpL1ipxjVspyOckxhVBaS
5dXKEuXeLo0mYb/GA5zVjMsxaXHYe8V5SxvJTjMRwIDx6zCs20bs7zRP9hNvMKt8b8UgoQvZ1gPa
wWGQQXE1lyXOcf78EkeFDK0dL4TAZI2arYo9CV+2xz4rcqWrbqHgFHtsN0t/2GYLf/BCUd5aIFOO
l65JsOF+rpWnqA3M48EetI8DxJPwgkVBPPvinO0y/wgbu37YNNGUC5xO6+FEoZQgL9xDT40KcFGE
nBdSIl4MsjaD0xZcD/1ZmaDPF+NMFe8G2+bNhIFTjR8yHzzzp85aUQrZ70WZDMJtPSCjxELlmOrG
ktvpBrX3Ztse0Jk9G5iVrRDyi5RJptxBEEjxaBzF0j24jOVCT37rxIU7kwN/1UHNwESod0bi6Mpg
ETo43ux+9A72+0yDg457yriZNdXGfXVMn3Ywvpr+7qS6buPZu4UsHALxkbVSYC8PLgagZV1Sjz6d
j4Qcuw47xTnwg+1sKoD1DqFFlyYIxo9AdLBF8pW95ZbYWo+MSWwZcXDFODV/eOaG/9wf2Remqi6F
W2RqvbwpK1LPVODZ8LsLj64VCt6ABCCvI9FoOWR19UulBVaHDBzCLnnALXeFb7dtDZJ5vzeiJr9W
BRJ+C0PPzqcUDMtMSfR6rRQCcmGkqscsQKZCcN9D6kUzb2HZSrHX6VkSAlGbm4ZBu1hutp+aWW5h
SdXqSSp9xui2sefmM+/vvO60K/J7SNxvYEp1ZWFj5jVZNe5nUuzOAZ+rYt6oLhkHAKoEFRU85mR7
9MLZXvz5fWbGmUGb9c1/bgihDB8QSQfMs5/fb75WV4T2f91funs20fRzrfiFf0La3XQIIEx4dYwH
/Jn/2fl/hCJrhPBUzgpH2/WelpWIi7vU3jxoB+KW1wq8CS3uNvIUX7bDu9Tk7bbXW7ZW3B74pp4/
2a9rm39mudiBxOta39onVGZctQSj+hIS1nzMsQU3JrmQVbWp6rqYbw8EijaBjAVQ1QWYc4pRaOsV
4OnmmEn6ZFoLUVeRDUy600zsYn7ZSZpIXrHAE3pRzFXBAMXE2id9RjZoEcI9EpB1m/mA45zLeyAf
FU334KshPR5TA2ggdptzgsy0fBmsAv3draG9w29kJUErqZdnE+vdQ3F26rP3xdXoWCQjIDed5yaL
lhPBkVve4TKNCcbA1/fZro03Afvrt5K+t1HNnw5laqCTjWLaq6FO7RWsmvOeRuGOW3aVZVCha3yN
weLRvmf1/SxazfT1uFxx29R/uARuwHm6QZxjaX6D7MXGjoDfxK8TaKKs5eSi1zTcVRwdpS4ucNto
M5g3p4EwOToTw1tZXI2ECIq02Ti8oN06kk0YwUyYgzVgDMaJ85gl7GymVTuDmEHoZrofgclf1Riy
tHFhqwqb6R3ef65jX2xEhlvWP7AXpRji0em/9JELud/mQaVLb5w0lV46I3wI0Sk/Y+zwsicnEqRT
0DW/RVvCXq1Apz0DLv+AM7DOvmohX2fInpdq8KTGZTv95w0PXdCwAahkktmPAWu/7d3uOELIXsDq
UyDpjg/Yd+hdmKmM6y2XrvbJkhh4Ky6jv1XVThDsIC8C9YUUfqXaJ1h08bqk5Oteagv9INJMOKSd
IJ1VtEzCJSIFfMbmcrf8WSAEBF0kGdunf9vOPb6meapzIJ4Re58mSR9WQ8nOQT3X1wydmzIanFAx
c1YFsfH5p7vLUCnfUisYnhCzS5AgCn2Y6uoly0/XNRBYAuPoENG7EENgU2apE0+Zc4fIJ5xPSpFz
Hnpd42PoHp1ZbtNRS9yiREddsy6YJr8ukAplT3wJly3WP9vhXZba6KGOoVEo33cbajT2kjGPPlCI
X7NkQAbcAab0VGIjGumoIhqz3gIFmXUwIH3tbwZ8X8Z6PDLvwfSJxrZ90iHQn84UYjkEV0jEBzcx
FhiuM5AZ0Xx3p84yuhQPbVf+yJdi6Qg6l8DLmmTRTxJwGM8BSXpgxWPpe8AvaXnIia1Lo7dvVNYT
mVhyR66FWiZ1MFRIvMaAtVfrKxU+glxSISjr7r4275wTk2bHoLHDeYCegh0vBy1iD0oJpoKszR7K
erOhY5YrC3K8Jes4SoBUHhgfMTLd/rqh3xo8tu9OeGxytZiktXLfJfJ26y2cb/bLYOjImvIVMEAI
c5CJ2/UEiHVhHI9QaHf/QTwqI++Ws0eqc4gS5fHb15XhvYsTpa5SwIiFBko0IVC6Ro8P2T2K/WgE
/TNQspR/VtMzrH0sE4PKAtZ6HRv2dt7KIazhWwqHS/kFQbnpFUhONhVz+VD7Mxo4SVvv5IT95KBv
Gs0krfWi0VRjw0BY8x7tVLGlufop0YPpO+lWGbd3q+gka9MWbx3rcFzc2NvD10yd+yPJvQfxMMep
MDt+ykZN8UAgF+OLpRhldt6HBRy3JlJC4snvBWLLaRX4SDvf3zO5cP6yRofPmxpd8XDyjGA7//OF
fQD4L/vrAzdqYGRouJVpC0YfCU1fJOqPO4fArPjcAqdimLY1TS2TzkXra3wXeR5MyucOjeNxE9fZ
hPAgcbxWFiUtwzcEyg1WmvMJWvduptESbaAB45g0ZHG5yAR543S2iYL8yeYLIod6LdH79JXUMpf4
yVC8PgtIqJeynCnlEzeayHu/hre6W7rwZ5Xnt5g5Q9C4Q4Q6E733m3Cml3sI91lGdom3jCcZS05b
s+zdjT9OygyVlAu+33UdGfudz0YMKLdIqpHYjZNWHPPnsKwHSV59iK+0g/UI219pEVZKtWwI1NxY
rJd23AS3kdbgEiGkLxf2P6x3e8DH7kSURz5lNpsTqXTGoAYK9ZTwbQSn59pa0+lV2nfIwDdG9yMz
whIiiVDlRLyOLc7GSUtz0FoZt9H9sWV4IJXh0j6igSE2KZUZ90992DnI5/TDPyPCJRisgdhGcDvK
S2u/sp7tbJ4MS/oqcd6zg4sZd5+fd+Ixv9sRg4dXs7LB9Loc7cxKTNj0a2GwtHkE04pXnXB2Ihlh
9gkRWIfRFExEwagragfZIQbpdQwJle+nmBsZnXtYOsrdN9kDEE01fNQ9Z34FG0tgCIG/s+sceMxn
TapnR43QzFOOdM0Q/wSnU9tRJNFJYQIGI1qtbgpgS7Cg8AfDWtlqepBxq4ftq4Ju8Aaj3/Q8GN/G
bjSxSkX1N/D0Uagl6KMidN62/j4/4EbtuzvOsGcxTzzEBSvfrNfr3Y31QDWduBUelOCaQkGr2B4t
35Pv8j7lAMOWZxUYI4s5U5tNUG3MkcZ4hLRPk1K9e1Rt6Xs5eQkDg2nl+pYc8XxtuE/1PgbJ+7yE
M6J2K+5Z1FetC/qzEZn95K6q8rZoBJZXghVIMl6WQstcl59rGgfb/jx9hw4x9vhcCSDIgas9W4cG
Z0vHCGj17qvmtzu6384MkVRD7yUAAYzGTM9msoIfw21RuAw2q3Sg9tAgbl+UNSsB/xbDsghE2rsl
I859dOziQCpg/FCdlU0KhTf+ZVkzv99MyAiRnl9TliAfdpffL7r7IWbuyw1DLa6kikdFsWjwEnrP
0K6MA13CBoH69pPkCzCRIQLNpe9gTZWmr5HvwXFH0sFlkRZLJBGYXtZDFP+vWUTtsPTzem4VCFJX
tX6za/QmXp3bETIsHh+UsOWc2YCN8oa/Aduw5O+r3x/T4Cn77E+uu+1N/xUHckL36fMQFby5to7H
rZpddJcbrCpLevgF3XuYdUL+IFD5UuVDIIXfMvX1OIlvoq/QyT2jk0nYUuumL4t1WI9bnnJz4Rer
oUr/ASDWIwopll5vVO3gKddvj5cPvj+3t+Ci5i5jy6ut15Nqi5oX1XFHMv/03hEwh35RQWJtd+YO
F3GRcvISGKLq4WOhiwshgurBPfuZGWdQVbv/OG37H6MG+ugIN9Z1z3+x+oO5hotPrjIE4o0hWi5c
dg+utvijLcOyNmmbgB6QoCTBQ5inuLeFQhkQ7JBZHCaNoi8lktwXvQFzRKYt845YNgMJRS+UbqoH
2P4XZiUQXwlHgHwbILTUNshf+WHpvJEYipRJ3s9vJZATu88y/CfH7WVDICc9b5idU7FUwy683uX9
RZ9WQyFXLUDTRLlMHAANx3HvkIeZXkurEo4n0cHHf4YZWWv/ae7if9a0M0UuzTikbrsWED+MLWC4
7XY5VZjAd2jXIzJtnYLvhLYyRnHQ6srkloiBhcAyIc3UuQuyH8b9APry77ZD+tiY9dzShRFDvvGx
CPqxFmm6gNapWLovLPjU28KU6ueux95+6z+28TsYFsAegCVgnEWpRK1PW3xZa74Yat7dijZqBGBl
Q7ga89BI+uIzMpfrLQ7k/q6oQutvfC893E7ikQ3F/6ONkcLzqYNktN14FTWiiwdR66L23V+gmkB/
rlVEzm8u/U2iNpPhsp506rr6eLehW/iEF3DQf85Fxk9sOdfkg37ltSJPMku+z7IruBACDnV2DOSv
cL7L91llf+yPswgFLf0goiUBephHig8o8/Z+86bN8BlJ3iab3GKHkGeSaw1jqNunAVVjLENXStRN
5/jLCLLfxyAuOkj/dXvmSuougSJ+7QEwBVI4zy4f5nZya2mH6wq4jGu9w0juDq+83bgpC7xnNDr1
jNfIgRAtmU5+Y+ihEfb51waycG7mABFw2IzDsNuidt3toW2Jy4Hv940mARxOtGpZApyUP/e197ve
gWZUI+lIyDJt3aAAzXp51h87xtZR5VaWwcGh4yCorGiQjrUGVvr5mv1y5Mzmycfpz5lDTA8SWkdg
ieguAfflXI2/MBqpZVcexYEAcCWxZPMeGwMDb1TLOmrXIlA5b0jZZba9qMNEHNX9lqXpPEl9Kgxv
51LF1De2e2luKKwmvoV9/JoGe63Uqpcbxd/9P4VDox9Mw3gO21ziekN1WCJyL8J8QUPpYoQ0mC3z
3uYE6BExolg6MwAJjL6gPitW7kah4GUWzUEJ1h1ZCK1+uT2u+wzpLDEI3CvU7cjvT7qi+5y5+wbe
0t9gtalK9xwylgBt8Uv2a9zlOQ5zM40dig976jxi8JoCI36cezsugEVcVE8wrMqNNe79HlAeM5k8
SmkacQnKDXTCJDP76P50cr6n0UINflKB9Rg51rko7GceEkX2wDLASvaALYgov5TsLkl35fZtikak
ep+ImeRY9gpLMTyorouAruRDnGcaw2YAntEiRFcS7tZDOM4AUIlPIhVHuqbw3GuRpG7LReF5F3kC
btBOOLR9T6/SnvoL5YLIqGW0wUcmCmVsRew3qAo6pAR/C6fqYV/sJ0FIyvEPjPmdJVuUoKMBGBMo
CurbPVcZIbnyE0Di7FUeY99tvxnadjfPzi1LJeD6Ok9KeFqyYSHLX8VfCgNFuE34uPe6PTcGlOQA
uacsuUxdoGXLd8rZhwpXbHLZRJ/LsaZ8nkmHQjrrTPJ3mgpkfCgm8/OPcM4Kyna1Clf2EhOsn3e1
O1/1LDSbiOFRi0JWjq3E6202m1Vg9CIrEU4tkXq+uLJDjzu/p4QQ6x1hNhVkccKfAxdzo/tzN5gH
aRmun/Fsizy1rRjhkWujGLE+CHqXHXn/7xPcpdr3TcH+//a48/kgKR0gFE0N8yUFRe9OXs/+LHqL
yp6dK3nO3DJ2Owhbkwy2TwVZ4bphei9iRLkEysePl+zIyUD2XkhpWfhi5LQUpx6PP9Pv54SFFa11
Kdmj9luY152iNf31NjbsYSg8brprls5E8qk/sm5dH4vGfDcTlNOzvmG1jyIyMzX2D3Xy30im+vZV
VAyaz0a3K9+MGLhvscghREP3vdW2vGWlNG7vgBmoVXFGNJ/27QszKaqEV2wGlaacaH05LE76sPJo
cDAuf/DPDzTfD4cwn4ANfgBdY7K21RWN3j3UKpMSK7/U3TVmlk9p/VxyQuL32hCdHdawnMYId8SA
1vHTy+ZNq3qQnlOl7hqjUF2vYkXw0YwBFC/UaxCuEpkHZT4PVDvDACbe4Zyf/l0gHy5Hx1vfaYiv
u1kS2VBTgwey4m95i5Z2aFcELRIAPPfz+32gUWJ0hVKBB2rF266hmVY1224un/F/YGzci3r689Qu
yB4AW5+zp2mQbyM9LPkaniMC644KOE8RherBOZOi1FYxc06Ya3jxVLhwF6NOrRX4++wuNHIrQyVv
KR76EnUG94vS5HFDFWNqyfp8iFpyo5DyyDnGN6jdcB4Rz1LPI4E4KqrHfpoUbK+quNXb1XlcziMa
5JjpANRwVnodHuFEvQ7QqgLpjcl+UIqhm/1AEnCyZQQtjpq+NSieQ3w2wLVxKaIkUL2sel+Q+3Tw
0TNljGO3DP2Qz8JZVYEIM+8/GNkTBWj2j2rjEsoL/5dMZhK2kh8r8rR2SP1wBN84rcOuGrCDntUg
Yl+8iaO1Vou6hCbDnqABC3Z7FqbZrWOGNwjGOyDsn4Rz7T1dvDB7cwnnbR2jPj2NtE2Kgs9VwGuJ
uo3TCmalIxibsMlqvjVkN+4kFjhSkLTYxEbmi4M4JL5+OgupWQwJAGP/sXSgzRTUb5Sv0CluUGor
0MINb5MoD/6aF1c4QVl8NJBryfolLVcjcGtNukjoiAtW1/jluciK8dTGaenNIZDI4kRMwCCNxV6d
3wiS1wKIIyqupo6OyJKNL4Iyn81PJ9cgBMxpzlwI96IJ1a9CYqVZVFQFndpEgVUWqAE+9PwXmOik
OxuBv7u84YdkqGUjQvD2Yn0JcJbC0h9gyP7ixhvlDJjqMilZ4TFWVlG6cUqp3JzU5RFgnwpeUrOv
t9jNe4DJ7P30s8nI59GNmI3NfkKG0yGeSUqnBMSYRdJ5IRIijdgYmI41t0cQehuYm7GepHCOl2MF
qqUeTDos6R7RwCz6fJoJZ+5k5pRSnvJa+y5yJ/XLOj//xyHL26wVE8hTRnpHiMhPFCzl/xu1aJRN
TIGg0oBmSkiXbJHBMeqLmIjPZWBA2zqtBv7mPOa6ec/rskJHZPbaxAr/JpCQB0HS2jjvBoAswDxP
SSUuYwF7vB2UmcLCVnn+E9HhyDLeW/Q6nidKcmwLcvxiJfi6PZ+TUnJkwObUrLZs//DCMql9+P0M
IGiE7LJljWQU6Aj+Ris7/e8ZTZUUQV+QBcv0NPMUdfA/Br23qkUx4ijEfOm40Cx5ySajDHELUaJw
Sgg/j2iUau5xRCtLM5RKnWrlUNSfTTL+u64XIcCl0+1xwR1uDEp9BtUSqTrfideb1seqYsM/aDNq
WMf1V4LkCaSCLtm28lwh0tjKPQ0Gcmx7BNdDiKH2A7j3pW3DUU/OFVfdyZqwWOxskGtbolMDx/Wk
EBlOirEMHQYm9tELOZX+J9Fp2Cp3bseojYPdmDI9p2wUvfhiA2gq/qFY763iYxBintxE/X9TS1V1
lkpxpqgVE5njUZRYHGH7zipu03Ikvj1x5Xa+4Ngrk6SVjus9a4W0/QmOyOPVIfeUGQtI70PImxW4
c5o6mFloN4aC1mWpSNGRsBIuNytxsbhEupkqByd2tPgglAqjBEnhicIcw5ZAs9Gh4ZcMR7OJRe/r
8M9K1RxHCTHs7PYQUo0UBwPAVQIM6r4KgH1Z6xyFpSo6r4OdQawIShzA4Hec8t0SBUgvKr7hSv5B
z1NNeYdDJlXxbIlWYbvZub+YWX0CtdCFSlGTaM7rxcr9JkIdfGOJ3e16ABzaVoQYZdm7zflZwNS9
pTIR/+I2/UazEehf4SbE2v3azf6MzbNjCXNKBXt95nIm+9Y/9oZus4syEz4o3Wqp5epsZ7Ceetlp
GVO7pIS2gAYtKiEtvyvNOvvOMRM4ylTXxSS+AeUWFw7bNOwuq0YlfKdtCJK9kFg44NeTp+K7dtfv
Bwp/kuVmTU/NFch8HIMS2Ay07HBc177S79T0V3R6qND+vjAhLbVZMUr7uRJDy08UmrSOE1xvSsEt
Ciba3G4yA3RF1wen7q2OUl2gESiRteeI/7sGZwGF4d1qrWn5fqzaQGs2UTP193/3suYE3Yr/nzWW
QCpueqi4iy30RjUljHGuZwvMHT+kweQZJtfEtpsK5Km3rm2B+Kov441MpapcGcOZXxM8mcsDwlFv
Ha4tSX1WuA5BcEVznRAUa73apV6wr5Y3cG6dLzFRz4h8JJi1criU/etoDLUYw7lMkHlgP5u05QSN
xtfVOGX8GU/jJqon+iC6OAkbq7+y5TRjktvKirBm/RrsQVhVWovtCwoCQ8nj4kqieMeCHw/YmtEe
VJxvCG4UrI0wmy+07J+cvmvKrx2DEaQP65cclAGtoIRr46JTRrqeDo51Q6adzdVZHptB5FrDaNx/
6CHf5ee2uuv5hqzk5W9dh53o8zt0610vv++SPLhjmGoJlLdS3+eiup2QsUSsH494x0kkbbSsJkAs
jqEWxxMoE6boKAewG4rvdQ7XNRRwj1ZypuQxF5xjkFARszFdt8Kv+/ELy6E+plCoJrGoOk61d+Pb
qKnL4hr7840+X36hJud2WiG2mLrEiCdVvYuriAbwY7EK4O6OGW+UYwX7f5UwDB1UFgygvt4TBFdI
yxB9dvn/HZxbvdFNxKtmH8rQ66PT9Y9b2qXLEm1QH+l3gdZVul8cH/Jv02Ot4Ei2uax99tgkehQl
QQdpeFhG8eMQYEA74Gsd7rgG6TikYutIdKKN4mlK0dtOVOFrtYV4PCUxk7SV2qW1xJ89gVWapsTk
MeuVgFi/GmWSTjgCT2RENGHwZx+HJqAltdrbi5jbBlnFn0DFyR2dE9Sn3Zu/BBgnQnpM/0cTdrCc
4UFZYliXFHLNKiCHKh+flfLtvb8G4ni9QSs8k+f45bODt9gs5eG1QxcZHtZC24ZN8nvUHAe2hVGr
SkaxHsUjk3Q5dGsoPJR1XQQz+un6bG151oo37NlaYMXK3yCs5Umpf/+EnNveQ/rYK8R+rn8RPNEY
XOb0r9ff04xekbhNKMmOQBRlZYPGPpe30ZoM2r9NCDVb0+5PvxKNvP8+Ys2/mls3VnzqEZPOIkIq
Yv3pZZaUzyxudZbLnq5FSme2rz+msNti12Z0t5DaN5ydokpoe/sjiJ5Ar7nJqKky/EjmOEpsxj+n
ZhyRvYb2V1ev/zA8V0YIYkZODzrb3a3y25PQBB5Or47tfw3Fvu8ocD18swwgO/yGnnNkr8sLxVVk
ZtBzMZcC5nHWSHyIlFlm2q3FBaySZl6GN7aOW6QgYbmHV85hfiVqdW4gR+/nUeKTkjVwCndOpcnp
To2b4BMAkVgPDlhj7DtgvYxkcs2BGPeceweoPRttSani7Pddbu8IbIgYwfmVb8BMXSOToJpaW7R3
tq4YmCXVkq3NnIBuWcUGbGQjiXx4fqhZdShXrm5JO0vd/Dui9ZlmUclp8xgrXdl3Efc7JhvCndaQ
Sj3nRIHy4s9CyvB6GFXDdR/HYb+0T2YeF9jX+rWxraSThk8jHSuPD0uB2DkjbLh5jWwcZ3pJcwzV
7pLwTj9snEn/2f8ddJq8wCOCVz0ZROtU4DDIUS/fk8fKrFXSn0HpuncT5nohfLCNT+9u3NxsClzs
lF/IWr+p+HSnn1B5lwz7/mmeV4q5LV/QikMA8KEJXqrvalnktAkC5I+WoEA3283NcD7v7uI+TWMb
52HhWSKlKXlI7r6gvDb5t0REJ4CSMtlC7hxqTW5isHgPixLC45r74WXCiGeccZ/qFrpLWci/vL3O
d2ddjJxm9/bxFGUCNu68YVYvJwZsL2jLn2jWlL94+BANzrWMwLCwChb0EGvmume1uAne8aBRqRdJ
6qXP98X7q4hOP6kSnvla4bTbf9jOeR6y5Me4NfWmlk+gN4WzqQfcU9jJwwzluYHXdesXnvaKzMEA
P5b7RXoAREhPLLDy7B+Rfj117K361BBvNMmz2Zh0O2W0s+yM81jd3sSQ7DO0mtZeQqgiY6JVUMQ6
Tuboj8ecC1wDmVqfuRvWfucOYKdyDG9n9w/2I5uNkEOAAV0CeJFLPVYefKVY4qyNlNkCqJEA+Sk5
uq6x37rBLxSTDRExvXmU+J6xraKTGd7AT0ykwma88YFUOcNr5QfdJtm3xugpdtx+t/MXAdAEecHD
G+sCD2sRbeCyR2KM67RWZep5uFw93R/WjnxU6JdfXLk7WSGtk6Qq1eV6c/jVgHbdHGRDmnfBUEbk
Di4tc0/vDa3KH2q2tcLrD+k9iMGMb+7/EPtFPFIzf7Oo+XPhscBH8NmqDHxy1FtnT3jjZZs3wpaJ
ZFnlqwCOmd72l9U9iup/S/gs8sw4hO/1BIu7lZSnDDzho8Bm3Q+KQcnX2eauvwtvcYGsBB8+TEo8
2W2FaKjkYs2vlpdPzeE6sZ7iz3QTEHuX+cNJ+oe7FnRWnzUChv+oalP8bdD/lpaWiqwAD6P6PWRa
3xFO/gD8Ya8ONoHyppB6s44G1VFDSz+ZlorYZWzX95XRiXrYLF2EQqEUN32L0RIDysNGG5C0qfYG
S/AHZq40LLVpHGb6tTpV9FKhmkkW+DXMKC976lOffOeO41NEw7x5JGy1OyIIMiJHKGdV1Dy5hVpM
9MQui282yFG6EG8Qin6PKCsY+KSvxUKzgbxjTH/k9DGOvxVvaGoOhUz+hOP5wCw3m4WzuarXMD9P
tpw3yTVjgQ3JMU12CNk63kX4AGsAWuWSr14ylojXwZqoNYSIfNB9OnTrzmTOyjHo/t2SkeVkMQ3R
KJvgSmzsRGPpvCz+9LXiwTu9pKQhOaY2jrrhdW4ohC27oAkg6Q5o46INRUe5Y/gbHlGAHQJWRkO+
rnOKVRVqShRZEtZVfmFcmuBaBAOxjBdOkcQbC49LlfA37SYIUe1z4Y5055rttMKGqu2Chny775XG
3nrP1p9h/3bx2RaoXdwpibgdTm2JUk7GXo3jXKPJXnsnarjbL7MdMBX9iGv7OaAvH/g3/MBFTmBz
sqlEEQwVS0HIa4Q6tXlW41MAf8vi6tfJ4+KFE9w8nslhPpUpMc5mMqsfMRvKALSWbkIDRPzNUEzB
s5GkV1lNpCcdcWo++7L56dZiBoi0YE2TWibBhLeYRRYOHofhajb/a6Xsv7jHcUd2J3gM60QTNpuZ
4uXLbFOCU6sP8jDJDx4OTrLncZQAuPTHCtVThOu/wWdEfi3e1limWItf3wpVRXPXWbOmG5U13fW7
ID5HgR/hToxKRSncyH5kqEuMmj64MbBjZSGizlrDGMbN4k2GIDCBk2W56aysDjr9sixsSrv87OE+
DMe5J72i88XcF0a8oenWDbo/YjxzM1cNz1Xf6SHKlCcPwww9K/WFEkqL/ShTUitUyMNfhDWasHX5
Ys+n8FUuGcOC5zZxsYaW4WsEGjauJhYJgvhLzf0BiJqkWLCcb3dvPbla8A/feZ3tDl+OGTrwHMQf
7Uifl+dkdhAz+JPhMJ8cJBSte3VmKeo6Y92LBADaBH7gvN4uvqlz6NhPmPXC7xWjq2KJ6Ukcgw1B
AjziOc+s8wEMqRtq/m5ocRAjxKOr5MDAVWhmN7CXlHDIvutK6H0+VV2fuYO7LQrjEYz7LPgnzb6w
NAH+VAw14mCVTcuoDgpbOX5/JWKLkBfclk83u6oFxmD/zRWADkZETZeWS21vfngOqf/0vmH+j8Z4
IbdK72gEh9Ts2j+gw4uxt4u+VzK6H3NagDqzGe1nj17Z4j0ZZODqSkhNmzAjT6gJDcUX0B9CVR7E
Zy0StlU8tUieWEWMDSUkQ0kxeX7P4uxaYLmnDgAaHAIkCHPgKs/doHKP/+sEg2OFw5OzvcP7+zy2
nqQ78FyBpNsUPAbTbAZTn9X6JS7Kw3Kjdwr99lPV0SvU3+zdCtTI161MDhSfs8iiesn1CVqmfkE9
ODF+LPaz2fHOzdb48ys+v6wcop96XR2DzQuCEkuZ1gIpvqXuQHRMRwb7Wu9DawfccPHBKLA2M541
2LQKGQRVM0Cn+3+SH7ofAWaqGF1QQ8fnXJnJsMhwro2bEu7ZT/3p+3jFp/K3o1N2gV3kYpMItTFQ
eScFD2qClVgoICnNv9+mx0mU1QLDds0tZomzXSVPLGDoUBh6Qh/vUSOps5M3KjTbmY344D6HxCwC
VZPVkSF7AQ0AXhEDzG/rGomXD+BB3wYs/rVeyWvbjvOE+EMG5WpW7L8zmd50zcNezhcN4OwzW+h/
Vb1ykO+6kOtPqyR3Edb9Oi9jR+EETouYa7pVZYrwYAzS0poAuMuToJHu0N58PkQ6ey8XJx6v6RQn
rnZzov4Y+9ncg56OHLTI4W1b2zGe08iVppBR+iBnVJr6b2f/6IEhuuDwDKeEnmmNhaKMeUnAbMpe
DFfBdO6VJymmefkbai10xE02TGoaumWVmjy2hfdrgNKP8XjE0qNKJ1VZ9wjtHyGuN+f5OvpP7M+Z
CQh+hvAB0lcwVx/Uat+tgqR9CHW0CGVvJsIJ6Bi0bG+VaidBKVUB2jtGDKFWsNu2jHoX9HfZBTuH
eSMK6/5ZLIEXViPOL/GWJqM8G6pZfCjue7iQ2aftoMVMSG6Af+Ld9ahJJTkRNbPJibio0pjuV8HU
5MTbIyJ2qfzQZWVvS/7MwstTYJdZxzP3xYc6V+LI1jKlI5FOGfwDPQQFKc+OkhSZ9qCo7NxM2Ueb
HOYz7qhWIxnGfjKCqjz6xe/PnGcweiP0D1O90NA9frNEdN127DWDXstMZglhsfRzU6P6qTriKaYJ
JnTqJRfngs/t6kTpAqKexORjRfV92h0KwhaYnyLH6p/jJflV+Fqsb3eGC2bpKtoOZkXo7aRjewta
/06+Hl8ccVdP/FpSu9ys+kNvt3HpkT57vjnjIpfccXIwVt2dHi5wDjeDmE0UPwk2kOgLzsIOTWy1
F1YhvKxH/IlmnUt8nB8o+1zGznmCTR+rvSlyGGch/kEocvoSRC6OABjta0LdHNGr+KGJVATMhVxo
SMZJQPR9rmkhcHnuQ5i8+VVDmJl3LF63o5VSeIA8E5TISdqmXIUxNpnmkR8TqZr1MExY2J5DkK+B
mQzGh3nhK5/DpKxD68CclIeyoYqjXE4owc1a89jszHDle6G70UdkGlO15WV7B4OmWYr71h0ESC/T
cJEZno4PvgqXSNbOffWYtMVMDLN2Tin4Na/FWIyn0uDseHFtj4l3HW6k4mxRuXnza7YghNNpFHQP
G0vz7jryc4mk3HFFZBWfPwr0fOXfnHqb5qytWwxcj2naX5jzkQOSqx/EwQW/d9vwVnI72984PA8N
a97cVDsRgLR2aVBKU1LOq3/CJuRVVu26chMNOOywN63E9T9/rx3nl20oJ/Gu8whQTV3kwvNmhZBX
KnM+FrjXVh1ULa+Ygxs0q3wqgdGsP5R7p+7dJsdHoBsx7DsvT54wZYxTV1KzwEkohkZCWspkmddd
BoJW8HC6t2Q3qVmkLekDO0VztE+8EVbtaV3BgDcquO0k4moYcBCqd0eB/hffzKWG8a9+SPwD8jt9
aQL0WlaXfwVdNgFnUql3e0HZhUOB+T6TQ7PXH9Bbdss9gSUsteSBcxhVxBbqfdZzmqnHju+ibn3X
m8OxcG4j/SCk4luto2CpX6b8MQ1qlf2YHTiIPZ3aSIpbE7oeRMFZmb3NxEybtTbzWFjmBghPxUFh
fQGEG1Fxfsz4s/p6EYexvR+cz6juHctkvCiLo3QcYa2QMh11/17Ijqjmg36e2W3KtP8Uwvw+ajiF
Z7PdSpbPSnK8VB9egNkIYdFLW2gBSdfjWsAiwv7WkKsIQwMxSE5DYA0Jocn5RjdIZFdboxaoN/AA
KssSxZx4SCh4ED3YZIn+QgBd6PthdhRX6CxrYDwNYjkY8mrL5TNtHx0Wo9byomw+sbtwMCL2mD1n
zKPhUfN+KBzvB2kcAz/BUezmrM5/CB3nqZXyX4bSNKzA4XjRtiXbDu6pz9E+0EQbAvcvAkU9nz1J
q5dMeO4rT1tF9BfcDu+AFUpgVlTjkWUdW7NAg1JyrVQGnGcs5qAWq5TYLBecJ/8UCUd0dozhe0X1
d992hlBvI/1zPs2OjQpPs0hqi8G9n4Fp4GeewyAWIg2u/NNVUsFIIbY4ZtDXeIi0SSveKRtNz5YM
ddleAeyhaMgH1ZvKvJR9xtGBWDv8/ylWBqhNSSjNhXVoy3no3jDHsSLc6xfXkVCtfSI1f6IOXN35
4igY/HxCY3rmeOkjFmGqlfZ/q/kwSfqD1Ybhl0knNpC9nvEvJgUjvSimjSFJG4GnU5vwz6WNPH0j
JxDVu+xiWV+wGOVm7ROkqyqnO7kBFcOjIiW8JIf7Sl4VOW53g8oRb/VtwPCmI0p3sdSBiGAD01ZE
eW+tZlqs+M9aDi8heIfnjXlgxfsiNqqgNN2nQ+iqBLvoSTwYAYXE2dJ/6OzZwyu52lpCdqC9zYZB
MveM8LtwSbHtekw1pdM+K3jWq3ovJefhW7PzK/iAT4tKzAPxz/o2wFnrGsu+lmQ+SlKJA6Yq+c2f
RROwSpMl51tNvgcWDvwdsWssqj/Vjx30VDv/2bT32dKs3tn4wtv1jl3S5oK5dHTRqH2wXeFNYa3/
95fOTE6pLkbyCc/H6IRBZuH5/KJYF/r5oL+c6zMzFUeC48vr1gfUQ7zoZb+tKRLlf0d/A2K1nJHU
8Ok13DN/ys4QG1GF/AJlHcG+3iqnyea+uhz9+76W+wlbdIbjq9YFR2eS3pjGsvdlv6RYek8Isyn/
2weGqlsvpP/MBsiFLNn6zN8T/tZJYI+2maceNM1/A3fb8AKRvsG+lowWWlOqBQ/Xl47BAho+qEUB
1tpkCpqXIyvcpw4VRw0O7uCPQ8qYMynEGAsR8jyw5zWTYQW+/WFhDVCv9Os7PnE4t4QeBhVWaIn0
3MaEcKf/bD7Cmuk87Xg3p6GXpHOoLKMTIge0zP612WtSyAdr7heQjLRUTpMKxEsFZ9O4gObYB78t
qTzGSCRxrMgWhYcrl+WrkysRCbNXcNPWwpjWk8ojgLRlin9Fbi6Xz29ZsgznfVRdjKHDcdPkxtfg
yGPMWY4tQ5eP3BVQlHb3yz92kaMwWKPeays0BkYH0XvgM3P6udUol+wjCAkFI845YD1qd4Ctgk4S
vcAlnvsGSucGueX6CICjKGvfdjibQp937WjNyQu96SCz9wQfoGr7/SrpOaNk0dy3CdYInVUC+RLM
j28vb18Pdn1WJBr4ZoXkPdwBlKi3akzwxyoOGiqGNsprKZfI5fKDS1NbeZzZ13wFbSAXQWsfa9qU
5FxScIOTwyx3em6T5AGHmnau12GmOc/xdcd94RPuDZXP1lDPEKdZmst1UWzHc9KyEtA7ULDX7gSb
V1rWRZRDqU59WI9JmmlGaQLFTH9QBqcl7aRYHOKQDKyfoG7WWD0a50mg/e2+Ir+SA8ht9R7V0K8X
hZWJJ4NuYSKmfnmaUEudC3JpJH0iHwE+Tv2Z/cHJLHci+zrP25bnWo6JGsoIykFSHAYFP+N5U8vV
fBH0ZUYfU7Q6gFecufoH2EPUcY1PajqClIQZZ7n8xFk9I1YX7vDG/Fx3EgPzjlab2Kgk4muu50Iy
BDW3a7n34neYj3J7yp6aRuJx9AQVnq0OR/sxeArRaQ/h/Njrn6zrAuDA2xAyoHAdEt4e1So+wfI6
AXZYTdcfm97PITfdfe36jXeQCfqfz5rgAQYJ4oDnt+dXzSKdcncBu7DG4jbnEQ9n/63gdQsfmwjM
R467SDBdDHdioxxf/2elMF9Fd0JLznaZijDyeYw3tRpmuUKZ2FijMmnvl5CcDsJqywwSwul6HSkF
+Zgdigd/zxncwbcCEjMoyNb3Zv67pw0odAvyiBUfbR0R3ti+Pjtkxi2MFaSMlvnGf7kGmWaU9C+7
hTZepf1h+ljktFxNYehVhcCzdL1UHizsNr+nilFwYLzeRpIVCrJmixC1+ytT0hLKj9cYDQfwmjMN
VmgvN4DBPMbYeAf/0PxzuuvV00Hui5JOZVf2F+TPP1U0GtjXD4RAlczAmKVsEHbFVRBJvWw19xNT
TsyMxxxOt9LlJpDgTmFimw3TffX8O1fiqyb6/0s1n7vchDSSNKocUEkfP7JrhRC6/C1vAUqZbzuB
pCx9bVOGM/iS2Nt3Fa8seLuPviPRQXTdDVnrh/uSS1g1jxOXWB68zWVjMZRWgPTkr4270Jvp/8YC
XReiujppwkau012huI7RzuXunvhD5VGiMJEYtkvw/XypS2l32O4fZbi+n4tmNLDitdxhIQyD8qkb
tDT4/e3wKaBfDt1vH3uRvnUkCF8vhSfIbQOy8CImCYNiGyvbEYPMCJZ28w726LyBF3waYsLah35X
juNfdgyceJlK+6SUzqGFZWDBKvai0ltk9QucWok/SIfkUKqUa0kB+bIFLsoSwrhW0Qr4cOKbuZsP
nMez/LdzsnFYGU1Pi5/AoWnBex2eOh2A+2Z2E+tQcgj2VMLla5iHbw0zpsF+ldtytzmLnkwCKfdR
XPR7zZkUqpf5NsrbbviM7z25X9bcW4hgcZYyQBjwNnJ15EA5NHe1cxMwTq3Yxi6lcvcHpf9REVzk
LVCaz7rZY/9K15SLMrna2EltCFXNzup3gYFPLcj/aiMFqIH9nbqsj/HDIuSifm3/UnlPDYZTKjp4
FI1iI0IF7R97Z1jthqoMt49yn+BLvHaw/7p6oMDAMf5FLGf7kCmwvJ+uo17f7Sey+senwQEvWubd
Rb8bKAqTWQqaKZPDgpID8+7ipId7J/MRw7oBecPDBsp949wy2hggWer+FF6iXHzQI6cLohWQRK0F
xfhwtDTsi5JIYTfPecY610djIJbrNf5oo1aTgLmZkGPINkNqdUQeA9ASmWlKttdV+iwcQmpAGleH
gf7CdT0FbMq+mUtygxfMd37fxn+bGMhr5RfEhbbzrswihUggQK0fFgFmDpX8AaI33/SDeudkbqwq
Q8Jj023AHNmmXiAftr7OCHTLbAr8XDCSLLeSdJ3HKgMQJnW5hFKYrAWNJq/0tp+z7jNy+euoiirG
UQM3MWjX05VrgJWSZzXMhX9FgQDJn6CRR6E9wjITm4XGmjF7bRLGBymc/hHHWp6UKu6Xypl+E3tv
ONSFSYm9HpW+S0WDOy7LZuok8k7nrjuMzXjyzd6WrxRJTMk8sODCRfufW6FO2K0FmB0xCaGRkGFt
JwgocG9Uif0th7WqnG+YcaNgcopKdVBCOD/G7f5BawskE+2Y64GxX2ryt5Z67hpEHEjCPl2qFW3Q
9MAENZmaxAOExtvCrcM0Dtl0cDn9Le2ziF+sTZLuYOeyrusLxwOopsRDKN7hIpAwh5gJGq4GpUrX
iZPd2aLWGaDY7v4uwxlHIOl4LYQ/LzXs8vivzejq4amVizWBbHN6mraCH30LcmTY5QVVlFWkdNdB
HXUgirRGFdFRuFvlIYxM0RBPMD5RHZP4hBrxo5Fz3r8qoYC1DPvwJ46MFTeJexLIkitwZJXWNxUH
5bbfKoCIv2Rz2WVZzINEmAmDz7InLOMX4RKkkbTn+hyO8+IQEUWNyZbpSL938IROflROwIronf/3
QzkjHXr+CLVJrzQtI1exMqzmCpyXVecpXfmwM8ymTF+Qgte4bP0/ajYxUDVnEK2UJVmrCDtlG7NS
WWl4MtQuMc9Lv1g+cV/aMzNZstMGEXaI3nwFCd39xe4rLqpUeM9pg9hFJ+srbZ1iDEix9xkHQbJs
y7P6o5ewzCda+3ZpdmwSwPiMQb2po/4Afyl5ruDSpHuRn29H5aK5tIjduovebYCJPn7pCge+uCZh
kLYruSLJFjDfeJIqHwdWQJmds1gJkmFEH4hvoK7Aonc3W0DWkAWC2GhFNA3/Uy2RXz92GJrg+nij
bk71POTFZZvgaG0iFHug7awX+RttfPVVY+z60B5RYvHdboZpZZoxTC6Gf9IrfvUm+7KtExOIwpfs
x2WDnL+X+hPl8TLogGQ9ONj3J4aT0bQjWNOsxgZfRyM7oVr8XK1tPns7NK4DgXwgrZo2RptlmBqv
1HmYMcEpw0iDOmmDT+/zIXV7jJU9yx3iKRD+jf87NGcXQO7F8ct3WbtRxRbnv8ocSeb6KOhJGd4N
BHYsWd9c/MHhynCXE6S9MsDyf2b2XVB8ou/e/KpdrDfkqDrzvZ7cmLDmiqAspI1v1b4MVDfojk3u
APVLYZsPghGB/hIW04fNuhbQ9sEpWoO5MkZ/GRpPvLGrV2Z1fOCHyz+eODIwOD14OLwQpYFHJfdy
oPsIfAlvty0kMW7BxS903VB8njgj85SEBAMua5MIITCHHEUxQrVfamigj7XFo+kNElu1jVngvTum
LwN3FJ81bit6dtHm7HI8kdUvi52yl6CFTO+1Lk4T2utFeRcVY7jpkrWrtwPmOKbEqp7w26DYh23a
oXlqrG6cHZq3waSVT3aggX4jPb/JS3aNMKdTjv6MJSeYT4rNDe8wMS/8b4R69RRP0gt7fUdZ9nTy
K8X+R348bpctQ88KynqoL/KoiP9ViI8qvyvMPgGV9Gyt0uv19M1PMwxVe9fdnAxMzNU6fTa8bv7f
/FDn+4QdqicD2DLy+Lk+ugYDqeDfBq7fJ4oL/b91BsDViscRMczYBvajKmEJSnXdEIYcLCP9z8Te
VYwInIVcEhWaLgQCbR24GfhaPTc8w0/oL7qPIQhI1I/HG19Yd4RrWhYdSbTMRZuABWcpq4idHwAq
F3pbKfRB1FQNlSy63VnGoq/exuc3dEErfllQIsgfix2aQx9kU3yH00+hFsR86rrRu1si0yZ4cYwO
Hvmll337iX8UDF1ME2fX3T9mtixRiY5anWSqrHHXdAgoVDWI1qdSyWTClRHfe8OXHc8OLysUgVl4
3NmAbPttAcZ6E7tfkLcD4CFxc1YqVM8qkmaGRyaOel+trATj00sfgg1WYzXV579FUjiOurf00v08
rJQ8T3Ea66sjIC4xGLqyH1CxNTpGwhg9Qmn4jfhBV6ggj955NUwBNJfkyrzBOZ+//WvxjFuHsw9g
52LG3uVcrBrVQYEw6LmOQj5eSvmcHM9HJex7LP61iTGz7HXy9cQM24LpN86upOovtrRW4LuyU1Mk
8jGqNRc8Y41Mxes4ieSPjTvXLnG4z7nnhOHVZBPQVapjIKt1ydmHoSQXRwLfXQu7l++BXk86qax2
mpi7EbMYxrroR+rnQeCYnbN0FjUvlY5VLTxWFrKAHeBVAXmzWSCdR9vVUbNgH7gyzqFbK7m10fWf
IF1c7SdSWJClx86kTe/b/tt6wwrGCWwxCfx4se0gyU41deeEsoyG2THGpAw/oyda5nxyRdNhn6/J
q3ONXsCIYYn5G+6YLpw3U/pfQGQjPfNL8rmU2Ofxoz5aWR9qmuaNVMreEon4u/fF+xIcFufDHo0x
ysQK7sadPNiWqgKS7nppp/hZjRfryZTRmVnE3P8mQ+gfH/4je8IJcj5/ShzWAwXT+5ijnLHpJsoQ
KlZkhTuGiXTP/lSyBBiR16iUa42RXi1O0yOb8n4BLExWwOxo7Y8dE3jTnIe4E7sGZ51pKxSsY9ve
us8Nyn95Tqp4l7ZWgx32p4mrhZe1GuOlB8fpye45Yd/kyHXhcjYCJcz3DBndn4D9ulM7K988yXxW
9EA4x1PM0VazNBMI3hV2NmTNSXP13nQFdxokialMt9BAgJxrk5i4lLipEWuvlkiljZ9Vmd/rD2/a
P7alvC/WBWY93O2xyQ/GtF7c7BBrZxSo6DRBQpCqQ6PtloWUAsmRY5vGRZGEY7HlpVKgqSc8pBTg
PFUCW4a5j9MjaMb1YHmbJeEM4/fOa923poIkOKL5ZNWepGlB3xUQi8dbmQGKK0q0hf7cS6cNq/xI
UEOQ6qh7Qi1Wq9oJro+PY+/junnhJK25hXxuX0h1Fwp2BUnwgCf0PuO8oNL+enlu//CHC/plcZpn
6AbP58UhMrTu+ZwzQK4n/KIr/opVQTud7DMyZ1epK9YHG6kVNlAFRClkGxoeXEx9kYeGkpnPLXol
QMHUAdrdhsEtnGEBJI1MjyZSe9q9FuwE3n15Wh3izCw55XxSWJ/nre25XTZRXG9NZwDEExKQ5U5j
r1jZWeJTQ8c+51siMpMWdXvf5WghKWgKZlvHYIdwK4IiTt4GVLpVt93uJqdYXs3vxqbTVCaLV8+L
DWKjbqB0uzm+z1ESktx428rZuRdwJBBMSVJthx/kVD+OD1vJuI3snjKkfpXls0dsFekEa7+kuLJm
s6l9+NoUeXAKoXVEApq3pSJ82nd7b1XPvEUXnf7a4xJys0SwkAFbUyjLouWUWb1TIrdOySfCKzj+
vbVgrGjg4Js/xohkEUtdRBrdZdMY/2TS9Y2/xp4m82Jcw384lRInJuoqMEB6MqwknIaJlmRNy3kR
qSJrPfUuWQaq8U/XoH61DHBUdCqutUGmJ2nOMzwJlRXE0LNQn+t6/Itx0VoriyBGVuFnfiFg6bJv
/CsB/Jh0Atfn1GQAEPHlKyptj/uWnUtvF+9iDwqenw97UpKgU4LD+MedygAYizENoa6KGfSHf/1B
OcTKJlKcGeEGoDjN16AX/vwgV9JJRdnpk/WybJysFuPHooFAMA4Jvxl0liU1v43RH8mq4TOOqrIz
xFaeolmQn5HQkB3Rkd9DyNNbtuBge9K6lygqiWPaGTTmnlmYZPoyOnAC9E9+Idquhqadk0axGdwI
LUS+qU83UGMeyya3NdE38OYAXbc+eeAiE9J3eh1rRdKgseQMbTlpiVT3WxvRkw0y7YLKtGVen3m3
lSeus4kiDHpJRhgXMq2hp/gVSk2Bt4lww0EAYN4qcluvKVEaaVKYJ0TAjLoVE4YC2ZEtJJg1v3zn
s9MzHorKaRdGfmT6qlMIpxuzpuOm3BkuHWcUWhgm2u6sQsN7NfE1MzcJ4ni+3pB4fRy9gtgHIly1
kxhFhB0DeaK/SEt2M+DbFIuH0M1rMSrD1G7N5Zc0pedmmQOfCGWJ480P7Pe4H91Iz18wXg/+Nz3q
oGhi+Dd+zSxsdIomxKIvdYghUlwzEXqyibyuDcq0Xbhda8wFWreOdyR/Ze6Ihtc8sVMyChcwfz+F
52lTkTraBo9tnPEuC2+74bCcXQP0EjLOXNJHt0tqkxRM53xGitxNzohbMJ/O+BEYfmFWSUM6FHkL
08cg5pNLDuHRKY6jy/VjUibIBTdn4e0QeNBLHkACRSnjrQM+pzmPJLKXdT8rFZiyfTnqTU2qLsdf
EGSQkicocYz+iB2LRlq4seOTSkNIaMKHaX0Jc5pRzC9aAlpoMSvJgRhWL3JmPd6PzVgl1PLV6LSj
1vU7CClCmReopteqv95ci/kYFOfi+ViB/2t3udgqnE03zi1ykXwUJbbXxFEpMZOubUGx1Vo2RvQ+
x0FpVeNq3gHpNRwx0q2FonkCkQenVk3c1JnVTpS/FIqvNWDwKm1IhLLGlC99QcXshbDBp87tcy+m
FPlQny/wzwgO5ESg9b9mP/tmhhIMcOC1g8buE900H0oWDWC2y4Tw4GBk/Az9ZDlhgu0DRvVN6kIn
8x3ODdSx8hZ95Byk8SXZvFH5pQ76o3CwKOf3fHo6ZE7ezNPHBWn+e6Cs6I+2wKb3FcxdAOTKVvI3
QHGiLD3oN4ve1IVeMSjYqH0c19UmBr/+A9kno+KM/LnIK9O4TkcH6VixCVu9jhAgj4dM7UisOdyy
jMrPrKLL1GRMqVwdExIKsUK7t82pS3oyet35zoLbUVWMx6Yw2FmfNYdZPJOjgC2bPTOpojUA0OTH
/lwAaKvE8XCIc1LpkXgacZGTspxY1Tg8fVxS7GNSlIpJz/CC5EKqA6UFUOI8oYAq3kh1V4tIxwmD
aWmtJVoeyKL/fLaWHWXqWt2uaFjt3exttdBS0VRIDiRIq1tykg9+7IjgfkHJYC+r7UrJ5c6t+j1K
0i4RlR6T+9URek4yLsKhN9xLUKYXBrs8CC+DapQrvG26C5pfjQWwlpPmipknpjBSdwpV57K2uvZe
f1jTkwluOgJCAZTaodPkUHeeB5Z0LRLgyKOoGB9KKNbNA+mMPD03r4xthYFQ4Q4hDVqJ20IYiqf+
qjke4CUd04JAjLu80d8Gdokvq0wD4x2TQGCoLQCO9ER5Ta0DcOn/toBIyozNZjQRcoJJGa4Z5Bay
48bkzR/431ygCIxSWAssQSLKdvK1o8DskfS/G4WM/v6/Qy8ZGW9yT0fri0+GnlRxqC7slSjcj0Tv
wbCRA+bOEm4ZBuAv7gAlcriQkBh9IuoP0iYWxZU1m0NvQv/IU9WQgiHLVwGIXe2YtCllkmKPchj5
WMcCWraRxS4qtgzPOfDdZjOEChrl2RViDXgAB/ne3vt94tNT6Z2/xJEdtKo2NvQz9TabO/oW4HP1
RWTEj32PXwCYf5F4mxhQn0oK9JrsM625EM8kc2CkIyWsFxG6Kj7Ps29JK8l1lcRGGt4iNHzZrL8b
CaJiRiF5kA+Jmw855Ou3UJxfHpqRwnO9xBfDifzhcDvdRWkO088xrqjf65P7y6rOJu1ujA1NuqMj
dcSIlQvv71yvIQzjGJg9/4WmVsVFgQVwmYjCMAlkoUWzAaw+2H1VESY5XWS6u5lDRjmPiCgkO4Il
dcVugywUNFw0ObQTsb+T0nMFiGlDIPQrxFTJIRaSxQo7u8XrB76/JDMMp57yZ2lsVKd2vGm5t9TX
HYXz9BAvtEV/EVDXszyT+rpAO+NlM5+Y9ykIV3NpUr3IHAtdDU6CGRYiKwjQGVxYQpeSeNhBkjAl
6Ni+cRyMIBqGvph3KTQeA3kefrq7FRLoOQDozadks0aH/e86btcNT+9o6LfO+RYtWBTDMy/ExD3R
wvH/GqCvkMi0mj6U+vKC8JjSvpenmg2dbMeIeYifpkCrWmKzq31PYJS8OBZMS5+6ljEC68K05ohq
UVmgWEIJLMtsMxrHTPikc9s2yyY0DM+r3iYjjEYCl1F+tpdkYecbYth95JhaCtYDbqQIl3WFtEY4
H4CCJ84ny/HLDkzf7pA3Os6NmeBvw2HdrXzXS1HmbWRM1uXiWeuV3zvIhdejQrUG678ZFnrVpR5l
gM+c+3KltxeodSxi+wvfPpYnRjV/qhBwI2vpKl/IF4cIWd7y0n0owOEVdOtvJpK2IFWwh1HU78rs
BDxDNWtKgdbuSRIF/Jg9JoX/oWyAN0SnULyBy0+IUyL1P+az3DWHHRwxVy762w5yLbEm6zi+q11R
IJ5I+frR2b5rJ1886r46aOKU8JS4j+mXPnkyTwFG+XuX4w9NYAy8+2+l9zZCytUtO4OyXXjZv1QX
tomltiv/Nrbdd3BZlKpSmt+3qe8LPjcDpZHbn1PTBsNaaXbvClYwMBj7wXvqHrhH4hUkJxHjk4rw
Eazvo2d75LbHxVeyrJqZmlvKE75sfRD+zQ0uRv9y85yq3VppAiD1xpYsOsD4AjPMSE007cQNVC0/
TwZHB0CT7/o4w7To0MbviQ/sZPeErILNqeQX1835A0LXU0iKA9GrEaQPMVMY18g3BkGQsGDA00M1
HvQQju/VynflSdsrRXYLKYUuz5/S3RLHZCHE5SlOFICH0650SKuUIIAKzpBun3nUewNKY9cDdW06
QPOGp8vZkQyVGX+AOHEkLzldrYRdVl1n05/00wImOzOM1GZrixfK6x01EE6fvA3fmV/n6nXFFtoJ
u/C3mYW/8aQm7DWH75X3vqhOnsyG9gIORae+TtG/Q+rMKqzhzI7RjXTnugDNgqxVa/pRQ9XnzOem
2+4hX3zfily6NGgx8zPsBYPC8ELM0bFL+Ir7GJVkS07KGcOydzMbxZZDl0WtBROoASeDkFv4gHp0
EcQiupouKOtVqE6P/w0ArF/eDmYRNsYsM+Mpe9snqRUZiwhdF9yOr3G2PhPqp4UdC9CBW3F2adMJ
/rx1eyITalot9edax0YuTbdfq6jRpfVqQTI0RlHHN5wQyd/P4t6GoxXTsLsQMD51dKLdbdHJ6MRB
rR13LaAvQRNC/BiKWfdkheE8lHDA6TaqiWt5h8AvAP+CUg9/8tBYH6FP7LyHrknZFn/Omme+MkIk
nzQMxzHf1JjTRDrCHkBKCiH+FzTjTgTpBhJg2tr0w3UkXYGsxu5SgFD1doNXz5Y3JCK1sK9dp2SY
oYUJoWia09OCBMJYsKuFxw4LcTyel2lm7tKumK+ACVKKjY4TsEGDNwz2gy38f4RZa+l2cGcLYOxh
O+mHlPykaI7dlPYCRfV7gsgQrS1Rluahgtu6bzvE3TYw7aMMMy7BaVY6IhWI99ZO6NIywGjpN9mL
qS5l0urtpY7DbXvtUsnEQxFGS0Ptg7u+jr3I9251vMq48GQ09PUy9YgZZ1UFUZ1NKMf4kX5UjD27
xptnI6zR2fMZ20vNCUEucylj8mqj0xYD7udOhKJcI2e4JzHzSaX4B1roR0NZaWz/Ded6r65ofzPw
vcAa8pbUZ1vrUGrCb78hNW0BN1CUTI92uf5/ZGxHLqjDI7pkSbasgTsIAcPTVcEgy6RjWa1/8NRc
o7qKcgH38oEnhpLvVRyURtTO/2rOAdiOSY/y1pJc23B06/FNjyokceLVpms/mD3W1vCe/XCnIcZX
tdEjV7wbVqcsQK/6tAGBWqvrtpoAuz4b6IBpV7b9TNb2wu6rOcfOi39Tf6WZNPBrf/gJDwfBQi5/
T+aJ4MmGNdSR2CGZwSxBkOFpExlmuRahpVOEJUbaiGNbr8l1Dlreh2mbmNQaR3VFy9xyB+MW62vb
HOuRDNmVIceST9pfXv17V8lcqFhXmFYKDjz/xRHDBlKXVuIxir6mYGuknYmLEpy8dN9sYThuzOqI
1jyDLkWU+9sxqhKzbIY87qhP0CtGb6c8b8+ld7cKLzfLVZHah0xBKSi4RwcomB0Z/nZlTair0Y1I
vGMfg+ytxWJxZy9IMA2/mlj5I4wv0QqqFZK6nfug4wK28THNhiUuec3cTH3sTbNfolpxWMY+y+xy
gRGXOc0U99ciS86oDNzzyueiQ0ZoTC1OqiAtXtcL9nD+H5xoQejgxhervlPSSBMKIxEvENlfdh+r
jkQcUjLdEKS0H1p9kq03ota4UD0ApwfAVl5qk77SLMbju9QU8Fl1pQ5eHZ8YUFwT8+D9FfuDEoFu
kOjvbOdZ9pnmtftp2nlKPb4iPClKpVZMCTJsr2JGtuBTqqf+3Qu6VYv9ZT2l+xKSPxxY5q9F5z2D
406/xCbVw1N8AaIC5v3UQ6SAtus2XMpuzCuK+rV/glJdzLLvxBZ63f/JOzASRvVkNS6CbvLPx/5/
Hj6O8wKorfu8YX+wAAgZNFnSV3Uyl/a+KHk406uNPjG4a0rfy71NRIKYo8PyQ1kfmMxNLF+eaLU0
PO6cx3vvf7SM3PO2cQLL2Zxqqweb1voJX8vE4/gST5Js5nsRcIC1uqyISabJpXBQoeI4ThPC3RPC
ltvtBBmyX2B2Ksub4Lw4A47QGaNk1Vf7WlkXJC89FYwvnJFXBlCqq6R9PqUg6A8UkWS1vM03eKpW
q3A8hYx1dB1i1QUeG2jxTdUviMJK/4HRiJawxKGfOBDV/zcxkUvlm74YoVb+tOWPDC7qx5p4hj7J
2jSRU7Z7rmrgrGBYFel2Y6tsRe6C2P7md32QwO1j9z7Krl/XKjtPm/lEVSvAHZ55KEGAWAu0061I
iJgGvzunmPSVluy5cJTx4mWh44WzvesBCB3oDnc/OTDFxMqCPKYQLq9EjoxAtwlXcUpafjc60dSk
04jbM1RslMTk7ic2lBYm2dgKcgl3it3o7n28gphnV0E87qWrufctMrU4swB/mXN3VcZ2qOkBAc7y
PkbeqJxerlQkWcuVeZBh2sY1tLqInLoJX3gZYPPRKoNRl7jNJl2qlJrfdjH7IiR+WX7tcNP3QsDG
n1Id2btyYnHMCqncpnQoFISoald1r7AXGodWqgCdAqdZsDcoKbLGI8QHTenfdZ1Oa7uFA6L6SdCw
0nQ3E+2QImvwCFCBnD9xBw2QNQ+BL0zn0JylSjB6gnNzpzHFDzyvwl5odhFiarCHWioLFGUqRnnZ
6OFNzFIDgHtkp9iX3aIVwESfcdhnzkM4gEUcCJWyYaUV+DA3jkQdu3yYvksDXVOFhZisXfMkqbII
qpPhA+r+GkQCaKcEGNEdDhlNj+JIMUDWhfjT5h6b7TL9PcaqjsSAUmtewaT9iXxgitaUOfbO4yOl
vP+9+FyxZ4HByktqsNZyQA7uyRGn+aa+ZgeM3OMFGmLzV3Q6/9xi/kwNwxlGwSERqDaKBBONUGxH
lZ3a+unCkOC06qYmBxpURsn4qDHslvOitMWshXq5sEdBPq5A8Zn+6DFAlwA3P7bXjcO5xCYyNdLZ
3KYFDjror0oQdbfUnHe6/BBnG4wxoGrvR6xg1m5LCA/SqI9THQQhN8npMQ8ejZvPJgnrpCHYVWxG
husMT2N1vrRnJNsJ2PPAaFTZ3clT5Dknf1aYfVYz0lZ91DVf9b8p6iCksWd74qCU8+4H1aeL9o5j
2JQn4cv9xL2CC3KFDFPogzLfNMSod62otGPBFPHMZEH2aSfMAHrPa/eFQmQa9kF+YC3MFb4YrtfX
YA2U2tRPUz8D5zHkJUaQVIbvAqEZ+M7sZAe1VJoHokokeIIeQbS4E1u5F1otYDb806N5X9d+kuAk
+28XN7enugD41PmVWg9Nnps8imWjj46+0PSZJmZx6LWKkIubrvcwSzBRPyuX+1A/19eKWgHgEe6s
A0QCjy0icPa/Pl7FWrgr5SOvn6iE2wiK7c9jMqZSLpblLA74M1A9esILbehHe2LCLLHOkgnvW9wC
usy13GDu7k4AkeW17sKCmc7aqwudiJFf9ZBa0a9hHcJagiw9W55wxa+/kUv3o7NdQJXdqryxdtev
k0YeyFHPWpAA9QMd11NVWYTc3TJqYgqIftDj5VOjDYFITr/CLxm8E7stXe2M2130r1dF5HSFAkcX
bS1nL9cyu11QzSSBYgKV30cp8UnAoJad/mKxMe2q6HJtQ244uaKk6NDviwzc4iKAAhOMmXEaL7Yl
CkUK3rrBJ67zBPSRMyLAdHfx8uK1LmoZjpGsP0fnVwUsYw/3OpD1N/BJxTC94sOo7qYYtp7Vur5I
rc4dFHk8v/vtUVjHC2tzvGU3x9jevatWpMc2kuzthzeX2tsWcx4RpIfhNMwCHDnX+BwwrSty4HKF
HvOGcHXQ9HNnZcKNf/Mu2wlhUfS6IbMif2cIAXUNAY9wQ1wbiaC0maoMHkQap8ekqmefo7WTNinl
x6L5YdxZETRdKgU9FzyBIfR5dhhI3iOs99PeTyPZ7wRI9G5shmfimfPp2AWob1A1LPgfXDS516CP
EeDC7j/ZYNtpZzXpC533hW1mLXAKSGElFRh3uAv11DYzAPFdvSCR2KFCVMLMyhgKU816R0WUO+BR
vUGiDsijHvcgQiK9X/WeOEEQXl3XVS8a7ZVYMR0kELOnFycE7g2eIFahZ6U92uiZ9pmo+2//R2VY
BeuD3Iu75huaC1tVh4E5Vyh5yekc0LxIfhEo755RQC5pIrmrOcW4ITWITX4N1qU/m6hndgYMXfKT
7jGlv8+h0CCoVkI8pSM0LC5fQ3w/mUcd9KJIvKbUiP/V0MT4JN1DFNsUJJ6/9as9Yvs9U4nBHxyq
QV3P/pTDcAXefIkykB9NT32b0KiOASKZsnUeaK0cGiu7ulObbmtT3RyMwy0dXPbft1T5/Lkwjb1l
3EkQTUaBwGW+9vBMuOoDrz89FgsbsI4UyMo5/ODuFm/hmvBGzcdrE2vgQVINxS5gIvLNIOH1JAgV
Kgm7QwOX2i1M6pjNfT6XU/3wsAm3ILZ9APavQOcpKejtta0haveIZpArLOY+GuiYSACAR2FhLpk/
ANk430OgyoqBEpug13DUcQCXeLuBVZzMu4gNqJ85/3aBFnVkLazNKAOiNU5nFtye1yfwMilV23Dl
JAkifBkfxl23JnsNWEM0O8N8b9brejZTRbb85Mi9Zbdldi3TFMn1fS1uYNM12XrpbqMZ1NlHx6sF
G2+7+l+spOiHhetg1Ys+whxcbkdlWdwIzPTrMJeM0fxxYxNeDVButQENU8VEci8QwK21Rs/rgtYk
Ws2u8AGvGK+tRoiSrmHEU6RCuT+H+9cR09F4R1lNSpj83AiAvFcZNusehcGTG7FqqPZhMIWRnzZY
B3xULEs8Mgl5FAvj3MSX+HVdGYKt0bd+hltlex0qIfMVmjAZ5z1SveTT6Gt1rtCJQG7Vjp1bF89r
omenAcCcNBB1HwjDtUQb+bAmtLFAJ3MGX//AMnyHlvs7auMbHusNxNlAAIR79Zio5fwyQaW28GFV
ymEz3+PQLqjqsUhqW/A7QyN7gKcVOYZiYNyEjJgGLOtijyF70L4YEOaKm2vy46xMQ9LLnE0sqcII
dY8U6jutSiEQHafkJ1aso8wUSyklNUbPUR/YGmIU2xQfsNE11EXxpk53I0KW+gb6tCJjcodqNXSk
RUyHS2j0qDtEVrZlj0A2yez8rg3f6ALXaEhq6/KZN9xXkAPBm3m0WgmcUrm0SPjBYRoRRraGG6uo
+CnqDAUiE5Z0O31aokMl6fhlAmTwN4dpLf8r/K+a/BADZIaZJCgMIzau+A1Mj1hxRYKwDvHUbgqF
pE05FXdzY9qmVMgv3kP04281cSExuhvob1fx29d1/IE1Qlyp5NKe3+LKRwhidFaR8j4vUotfBg/j
UlMtUcEanwgXtpdqCnuDbDFR0HFKg+1QRXrQx+erwU9ns9+a24C4Z2MzEPJOGUC3vxD2mqegicVQ
aiDWhAzFTjhupsUMJlLjmPB9YS+r3Lg/0C9BXNKnOWyqnObJerPrWPRyQxgH31+FJUWzujfhn/j0
oZAvfp2AfevJu8gACTqPKConqH6XCt4PxGwqN4fhBaUkhVNRgXEvl4FCJCwmhbAjAdhhnjHqr78d
57M5iRGz0bt3PttbLkvfMHZU7Th/30I3/Zptvy4yf5+gHMGiE0jKH1aTBu7xeOiGxNp1yag2D3sd
GJ6scwrhi2hwqskkwQNnspLb1nUlgZh4FTrYgxXiTFc9YBSxEXqIYgdHAAPJ6x4SbFLI2eVyp60j
nlZhtLkkIbvEZNK5QqM8NGUDKxl9mYMb/Ze9VH5/1udPBOBowIRrClXVL4LfSFQz4AJib+t9FjqG
Ym+WnvR5a9vKW+IcP5gYEX/+zXHsPuRprQQB28asB0vQUsyspYBKIZ5clARELvzAUJT9WpPpGr2I
lILKHW24HUB0Imqv1ZieEGaA8TSKGn+Se39ocPn1vZW1cIt3BYDbMZKJMAh5sldqkhTEEKNE4TIs
TnetLefTnjbR6tbYI0ydo7pGOVkkac3YeNXsTJj7DSC+DSUg8mJS7iv4QiAKTCAKigduE9LtZtN0
VkzWJxYGeGW1xq2AKOnW9hCYb/SQ/GSWPhmbMF4CG5MOVZqJmQpyeBcNlhPKUT5ooveuOG7CLHJG
fGnVoVSiHehY5jpPtw+WyZM89ujp05bqwyokn0bzvmA/rNzbdkkeWJnmiMFKwXZlthIPVMRUup/C
bD5PZpupWn5IV0M+L2ITWDYZY/tyrtkjMLMQdQ3RckXvDk/0U4GKBFzdHahLy16qT1GbykQhS2kY
bvIfJM+YHb/O7Z1zdviCFBH0M2axA7MjLFBZ4KZ8ZLcc/Jr9+/yUlT9xTKNiLqfd93+mqjjinHvr
15hnyuWxbrcYrnRZXbxPzOB+aoxCwI9RD6qOmE7b2GuDGyFSv3J/IuzlA2nb7yjGO3YcDm8UT1Bn
ygEiRAPrQ8RMO74v3Y04ocuK0ULQcHbJrG50X4g0WJj42V3LoI6z96gYYpKh0EdrHKyb637zPsLG
ic0NGEspoT/WgGu0ojq/+w9HAUB4ZsS0ilZ9PVX83bFrWVggNOZ32gvXMtZ44CUfytYTzlTQyBHc
cgAdd+CqE4+nHFCmaD3H/nKNVqBTDghBqlVmF1PVm6lensB68U4k8/PLNRNMwdk1Oy0OLM+PF7kX
cOFsRn8B7cxoD3OhKSiOswfNLYlEtzGGeNsbUYTu/ZypCe7cw6foWCQpIvRn6oQA7sa8dNVm5U1Y
NWvKdCbWOmxkMwnDt+i+4Ii5C08yEaxc3wccp+xytSAH2o07iUowm9OwcbkzNq7mZ+Jydtqm828G
YsqrP/6KnFcOe6+hyfa9Xu+hexg9ysWAEVi0IZHODPmMiDgQlM7jeypAjYKL2D2kiljEKWF9yCLy
twRbYMY457Z/pog/oJJHjN/PkBqNcvLk5lpurNcgI73sv0d6eo5Vc7o9W153COPZt6DcTQ2bBb8z
jFdlIsqM8D7dkTzxCAbOeUsGQp7noX3YA2EMy3I6MIKT20XONRAeIIaOy9gBrX7ZcdREHFq8yGrB
lRoqGryw/oWI81+iO0hMbYIYQMyKAedyFk8tACz6wBKj2ktljpoqhIWzAhIr5pTmVTNPTT3AF69/
RsH63/JqgYU59Ln5kqy6vZN1TNCauuN0J8o6rfVRUwMqjtvEL2E4azthGFKb02vVKOzcDZhCTIuP
EcgUWCphWQorrrUH5WIaj8fBaBUlDUOSoHf6cbqBx4fvv5cW9unnjHCVYMwK7zVL28+j97Q1dMuG
TQ2/OXbKkBfuaRGB5znxAXJRn1ZNsMNDGiJIOmm08uMr/gPuf+kyZGlVOuppiZTSfgvsKr86UyzI
KXXM3uPoevML1buijeMfI6Gg8Ays/Pc0KqMnIC/l48G8fWNWm8CC27IhFBxLpcnc86WGrK8UqpCR
Vxu5LYSYrISbXDufsnoZ1C0VuE4escK9qBxr00tvilKUpWPXNyCUWNAthtG4wqydtJL8fh+YW5Bp
wHliZe0xjhf1LvdAYuSuD5BTLcEXiTvQHqxn9j2r0oFoHXoDC+59s5RN3cMFX/+aNN9QsiH3vNwC
+lSCRKdKROkKZWKBIJALC+KcMYsk98UMB/jZOblrh2FBK0z8IMOmVd+EI+o3lkKfvwUb+gnjVEzk
JGzHwqtmebBzIDth2pGM+Wp0hpCLx9TA7iIzo3FLWexp/rg2P0iUCQPUmg8fc2dIKV/VfvjLBNYK
UurSUM6TcWj9dA9P7FW5InGeMxhpJAJ0btJtNNYVT/239OuL350xPLMnB8HY+Z5xSa08tqOuOiny
F7WIj1tDvoLjI87D/8j0cQtYYoNAWpdnBkZJzNq2c5bEN+Ra22doyE8Xw/k1TH8qlkHk3MuC/R6q
SFCwoiQIhYafH98JKQ27ZGW5I/IFs1nmMeMRts9Lz4vwYdvYz+SwzmW2hCrLeHFZf8aass9Zm6Zj
JravXsYdRyNz25ZQ0d4QqGFTNj5ENL0lxVBuVCEsSPpmstzYlWDShiwKwaABwgxwUs7FTL3/cKU7
Tazl/v+viEqEVmMVbQ5ZPGcMNxMaeTcLYZ0jWKUk01OfPq3B/Afn1w+6bSOCPlo0UhckJJxV0fst
unnJpGDORGylqRr88Gr8v7hPwL4J91G885vnJz/Uze5y7XhlzZoYLZMpfSw64JjeCAr2L4STFpLV
0VLR2GZB9sct4SNmtB7JkRZJ3gFv9b8b6mZDd9RZe61kZSsWMKJs/b8XaM3JdI+QmdvKm0z5SSCn
jtcFLC/snavXhZHMFUQ2t3goMWC8pKGInQpGo/VfrlTWkiBeF8AHpszQbieLFh7CvY1NVEsh1H/A
zqD9Ou6SI6DsIVOTuYV5UZvhWDGLLJ+48RZEuDgSJsu1lKUu1Kx9FcFnBKzAY26YRfNE5pXZEk8p
zqCHcwg+2VZHYmOC4Twyd3+9l5244HJ08T7kvL9QwMO4j2cvZSLlRoFohOkoiZwcVZXdyrYE0/aa
9G3MP1lCAvrr13EQqSCFDpmX2VlZ1n44QpgfnC9x3VJ/yfSx16Z285cAhOCeurWzrWC+fjl0p9+w
dbDueMQ/jX+ChKuMWsvfLXrSHIv5n1e1WWfErBJqyh7Nt4a4L5XGc4ZXFE/53xWB3V7zLuBxqnYg
6pyfbZrsT1c63NLTZqOzpHxEP2fSM2G6paIIST2g1gIqwIJcqvfw/Wp/fHTxginNaMarsS0wlpzQ
qM0bU15EOxRhsP9LyeRFpEW2wXRhVwDcLQomoFLdSluNq3nYMBviEk3biVLMfCszrYpfgzhnXXq7
ca5jcInt2OugD2OOSjRUnK24EJhHtFCEKZxJ8o9LvEUQvzRV5TNRnBo3N+0uhmy0ruiqkqxvH0AK
XTCN4B+VVuvfeSNlEL+KqfSLSzixvBdWSHFZKX1DhL6T8qKVxVAICM+hyMYmN5kE4uX6XmuaUZ9c
9NBU46HY2srIMUa7ihFHayuvXBdgLteJr1Qe78jZ04qbSujEQhcwyNA/Z1bRoOvgDEYs+UDtAg/q
qBcVxurbwbovzv7vppq40aZSAkQDe+zKs4gvVdSa43sauTpGCmA7LWCBLoxI5/7pgwjfGNFN2Q9v
6N6bYFPtan4k2Kb171uIYu1Yp0LKSZq2FOUHliIS9ut/VmS0vwJcLgfDFj4/bbTPTivTeCOvCCtz
fvpXRqZ/Ss2tIQE34Hxqr71RVygma/Vvd092uAwTEMdoXfeSspfRp89bo8G7xnjdlxV3Gkmr/ks+
Ye9WL5yMZs1xf8pcTlLaFFh05z0oN7cxn6lo51KvdaJuJI2SoOhWE/a3DVVuIcQKOdT5aUdMt+oj
4QRKk2Ge1JsRlGG/dXs9DNw6VFti0Fn5MJRmQXrdKCR/DiNrkDrSzyobCyEiXmsFLUXYs3iiE8i4
zV4LQD/PVKRGxCne7Cu8Y0OHRCRIYRjhZ1NpasrIdtJW5O2YjgKq4BL45n/LI3kXLHvPxm5p3oV/
NplWD1IzpuXpkae+5enzJz7nOpuUxdVlKm3xhRDqv1IaHCnlY9sMe5mFjgj261HO+zQDWgydmfDL
UYejWFufnFQRLVDakKI4xIwolZYJJYhsEimwhS1G1aQPm6xkOAZot0Tb3ffpU9fsUAaHzK2SHR1j
RJP+AuQiWSVbtESPi0tmlqJJdeBdifSLedIVSlYZSspcU9i0HAMcCxeSiCsy+RirzP4LORiGxT2O
Mt2gTlCcsrtEafFEP6BzHzvu5R6Uf3U1VzSUYQAXD9za3H9V8DH8ht5dOXYMGbxQqhaJxbpY/wjZ
NRuzWxeTfANIjKpOEvcMgJqrBCvmJRQ1Gcqrp7ZX3s5IRYhfLN7AGjDFjnBrl+VTGftFaq+hBV8F
kFAUXDm1avyHHY0vf0emNouOgWsaNASH3hUk1tWvFuqoHqJbYip4mU9AaxsR68HFH0D22FllddBC
H12+/twr6NeWgX+WNwExb+gr1db1gNV6UFVDEOnf3Xs5YCnTWFGXFrR59ztebAEFidp0tGln10xa
Wy1tzJGxBMSuQu/qhwVywuqh4M71gRl0s79/mNPhCCQOjFd5bMSyAZ0rZ0aBE2MmlEo5YBoJwbDu
5uUbyzqBaqcbeG+CYlrvmPgCwdNSpsfTY8cDtqG1SUC0SQzm7kXF+9z3zSBDHVI3BkCRtMcS8aVT
9a7rZSf3KX2+gwuZj33j05Z9nzs/15/pnn6jA/hNQLxUtLKZfe9XMDlQ/xak0ERh5BKGdculIRYF
kCfdY+pCYwlUsCKkZ2S4gj/6SzRv5yIKdOx0nA4VzFy7deMkujCuN3JYh7SzRtlGVdR5/mrF8WE/
Uj9SVhupB9gsj2LPFOI71xHPylqiLt0hf95fqFy1oefBQfA3J7WFBgsC7DjQQZzlQFHzUTnxF7mt
E3uUVoK312qkYJ131mdvCzVxPXiuOUOEVc/BDWtsDjZFi39riAIkC1CJeXI9nXUaDwXj7rQWoMVn
Pf2dGOtGU0qYo3NvjBY5AuRSPL2p3kT4BwDmUzPP6s4YlDYMlnNVDbg/Dr2bfRYfFdJFFLqg3p/r
0XBTN+eC/cYxrXGCHVUbUGWxQWmWWCxYcPR/JD1z3EqSHRFpca/LjZEGGQmth8PvNz4tsuzBZ7BA
YdYjspfUQ1hHTFZ7aA0poWbI5aeKn7VfzZayf2876j8zoX/+NQzhmEyY+GzlWxvbelzQjKg+ypuC
sTh2YxK3yuAJf+7WfwF8Y800uC/WghdjrrFChDiizOLh8s4pwLJrCy1za3b4TttiYLRGvTxv9BqP
NvssDd82wt8ISmb2Ip4s38aaEIuBIYGSj9pSPDaF9mOmnJ9067o+mFP2PuGw2jetDM452fR7fA98
Lva0OqzqfbcTec9xUeWqwd0dGJRLaIGWi7/nj7XLjTuY4tDhW2Ln2X/9SLRBc1ZaBh0R+7Hiw4Oc
TIWj1slAUvIvziOsJVxs1OojNuj9KbrQ9rC0n/6C05nckFiykicqWDm1SFR7cRnB4krf2G8WuTgH
kGCVReEidicWHa/Dac8JHZInF3TYf8XURU6+s32SCslKVA4OtCJLoAGgtRYyf9ulfCk35nPxS3lf
IIs7dIPRQ5CeyxKVG5iyGT8+p33OiYbb/IX2pdNUin3gCSh4L9QWYiDHgvF57J5GALz3D6IJ+nC7
PBlg2jbdbajTx2LMEfy3RjEj+lD+PW5IcKrqUA0kxdE2qVSEAk/TFGdOqMlpzb0pV4JZIp7id09+
jnfKYz9zX36PqcXbjo3eG5LoEH/2+3cdd8V4tZ8/nkPNo5RbRk+GMDXPXZfbbjkuYkVe/cUKkAii
jO8QkONWPggbWU7ygkVkn1n04FTT70lhrNb4AhBgM+dcePrW2YOEduJRzf8w3A7POJkYFgwJDXbz
+ySvqSu0bkCPkxmEMoQz08rXdxFrDB4t9sn5uTA4BjTkInJAguTlBU3l5IhFwSvx3H/gkSCuPLlk
k0fJYeMNXBmFjFRDnJJxs/dTFfN3BRJj2QaPJ5PZVOxIJYc+b+ZgJ0jGZz2ENm3sGMLRNgACXXsh
7TjR4buDBgvmUIXLygbeRd8E7PmA2uvlbq+zBzExCj3oeTUUlyt4jjk0nU51vp30E1oQvOziOoYD
+OU52rBWHr/YRDJOVvwvoYnJzl/9flwamDAWQ9EXvEAMwp/0F1I9fzQyPKzXeScStI+P0uJ4ZRc5
ZFzf3ZYyy835nxOZae78ZtGS83CHzHABh5KSb8BZ5A2BiucluFaFRzjYJ1vmqZ0S9fmlAQrAwgBv
VeomhRcbGS5iuq/fNCaEf6y2gCfqmbWYlgtziazMXPZX02IbalVJ3emQerP1q3WlJI+WWTNqOAgR
HybmFLjjqv33kmjPTDaUSkxuD/FbdLkfV0kMRhC22xO9ISTSlMXY/2zg/UeJXvUDym8lk8g1rtHF
ezjX/c99BmnvcdmV5mbpFliLjSmkIkWm6JpUv+MZ3GtJ/SP8ITx5RWjneDMN+ot0U8yJoKYi8pBp
lojMaKhrpleOa8XO5AtpG7JpGPwOjPVnWT1Nca09L34He0fwPKESBoFUhXGHOvjkI4hkc7a30lZ+
/wLGYWiqMyb+SQGzcRZn5JOgKMa8P+o5F8dfSacQYPfzK7De/MwBzZsyl8eyq6bb2MOWtpEYYNGo
tSRpsIy6ZmvccCFbL37rV8NLDt8gWl8Q4aGuxPL5cihNh0YsFmOuUJ+OUmunlqqetZ3i2yiGWQd1
4P5PJHHj7FDRbBmGBFhkOxcKiKZgn0DemAsnKXs2QhPqpl0UiAajfgQQESWSfv6EzjUzS3FvXH0/
BsNgGQFUXWixdSUak37jK/Q/CUTVsMPHr8EaWnSoZtXdp3v16cIvs+LZTcx05o7CyA/9OTgbocT/
m7tcPxofKJ7Fi/ygJYI1bK/j//WvvDUqfvssIOhMNUVGLirMQdClLdbe4YsTvvUDLyfXowv4gO1p
DE6QxZGYnpX8tCiy/pcBtSyG7ShW1kHuUs7yJOmQiIVdB4DMYjC2FG2Qibegm0EzSnNBsW6k38su
V4kHDB6ohetB3lW3fSncPiyaDO7PEUjUvuRo9uMeCMkYo5SBtQ93b8vi7endM37f0z8r7WfD3wvS
sKsrs95d5pI6KpIFCvf0QWFagIjM1c4SMmIfWxnzLVubPgLpq7b+Mtf2dmSswSsHdoDIvvB4SnC1
XQJNIdhSMYyyIjiD07uULgfWRrIZp6rYfju0YX4sJOGkxza6vnBHiR1nuA2mcO710Jqq1iSxc3M8
hmBWqvp26PecMoAgWTBLNiq0gVmnjI4sPukJnuupqhCsajlYt4AKoaS2CXe85/sbfhFtu5DTiiCS
ne7KUAG5A41MP60iuLxvu2acyQTzw4awJpbLiwcjVgbITR6wZF6meYSG49GXvlJHleHQ0yDuUmFi
VG/83At531gKkbeQSIYzs5nkY8mbl90sfVZhstRK5bLdwcZp6gN20WUa7SdFg1vvvEPmT5cySiCS
N3RhkatIsoeiGcHm21Rh5FDAQ/gasB1Cx72aM3/Z9BUtBq4TgI53g6D5FcN/McaADs1+AnqQbhuZ
uwRxWhAknB0kg/KSiQMdNCt/F01vBMs5ohv4YvmYlDIeESizKpHmHz28oX6ceJc7Bfnmt/XxcYyj
iLWTV9KY+9q+GQBp+jORX9T4Kj4vbannqcM/9ob8vKvOzDCD6I4k3hgZEfVAUIEk3Wkz8McyLEfU
auolTN9zBOt6NHre051AklHBy8Zx53ungz5DbjCyNzhZvlV2q5jjxTUM4zQJe+GBUJJKjezbxGHK
oA+adXLi9Ua1aXFcCF4AEXSLHIRSyez/Voj6katH+5ME5kqMgtt8pkTWU1fKbcj4T2PD2MYGb2K/
k4ICksCebPcAuC5JYsqjqmIOwIXmd8vINDPy2LdwMeFKIKZegjPcYdegTUJwED9yp3jab/ivo3ie
nxUF47LVtXMIGjw0HreC4rNxZNagaCBbtp94L+N6naSV4nPDzXcz733s8oqQBjTOKiAZln0sG96j
87PzXzBCCEBizuZ8Qt31r2H+S3CZJSaGyAAOayL5mCTjw6/G0sponTw8WUKLBbDdoQSvkuEdhsLp
WPfEV92AGz1FWD1U5VfMF+aKBhhjzrF5+FCUz54OtTGB88mRrbfwyunr5cCJdRuYJdea8tqvfqCz
ffjn62ZwPWWRZXVhyxuSFZM5RiO5gILBCMkBx9gYmTtMyOeuamv53LbbEq43buPBUrQqDxwjALAi
7QFFgbpVROG7pcbBD29SXKdXpXntqMP3AoWaTCAb2pvjx+R21GjAwqwjwPkvejSxNhsv+/P00I8H
FhqtEYYt6VcKFUgH4/vXaCIgdsWYtZIo1VFKTlrkFXDwzEjXgh1BJTEsrJl4AmhV/h7ro0WOfADb
eEdiDQlFDp9TWxqz7bPptERf4nVjOy8PbciS7m/wFl+x/a0dexQqKRi7X8s7pHcbRaP7+BcOMWrJ
2HKKrqo489AzrAgkLvDgqAoE+lGvYzcrv9oKiKRneA7tCO6k4Q0FeHeNw+c2dUWG0AJjU5nGhQoQ
o0dZzO4Dy2vhwFnPrGvYbTUOSTCM7uFdGobxDj3aRiT5Lcocqbn7to4vshufeLOC86UkCOiod9XW
llkc1YryK1FyfnRi7u+x1luuOTWuefRimiVSkMnbOIGwvQDNhBBEvXY4LQZ0X6c5QLVcPg5a2Svz
jOxZ3njyQTKYJwpgIXPz6h+diB+41cjpO2wAhPfw8SfdomE5megpO0n3EpFwQL6tgEsPf15TTeo/
86Tj7kVzQcWLDBH8TFHiPlvcaX6ilx+FS/f7lhHHcln4GQBtorDmIEI69K2lmw0+ZBJOSpoFyIRi
pWRD8+OxIFj5T9h6Ftypp5F1JbrezVsSU1oSizfe1+GfOUygJKVc6ydS/Lph37FRtvB7+K2U2+0p
zmsVZe6Mjf4kRPX4M922mv+fCZWNhzHSYADpS1PPEVCjgyvoXmSx+eco855yicZd9u2jCTeZuR8+
+/h9rx0phb4t9GaGxskOOdoHjVRo9ufLCjbsw+U1lVsjjF45ISOD2jWaDtygRkRa3HwiUrMJ13AP
gUy8wvrh+GdGZuzL6y15o4TuN3ScbNPAGkJb2CYRifV7Ed1OWEgJN5msCQcIKK+4Mn6flykv0O6e
+XrvzMeAQdhIYQBGUqAtRqDKWCKdKv21sV7DN2/0VC2AtBXpRyS/GDkEIruk4+WNTr1fCRyRrp79
VlxgaJEr3qIbSPUx7q80+asq46NE7LWB0+r/oD2mH0yq1a2/TiHDQNX9hH3w78CKm1Zk6cn4xZCG
VOVxQoB8eJwD27FWPCLeGpYorHfuWNHbSbEwqP+U0zywE1t9i+yvvecuSmBvGNfpKMeHbvCpNyh6
rGFouhoeZdR73E/3PjHUHV8iuf3XaLT4CEgzzxbNgWY0DuQ8r3s+54N6B6MrxONvWxBKTzr1U0U2
cLrrhmpq8fYhvkSMHscUdq64wX40hbr8D5JnAEPZF0wyylJEaApg6Izu3pX+KhLH9miKqfYfcs7v
obF/nn/vBpLvISfxynD2PHY7LVzv9rpYUtSCMYek2+D8vjzQKMx9milSG+oN1QTp0qvG2+BHvYLn
qDUb7ilTxE499GOol2u1sTgHZjDPGK1KWKUwb4apV1jv8PDvtN7r+Ofs+QTAXhFOhAU27hWU5/ZY
czm32EWWhCukzRqZtBu5Q15CMU7xLd66rWEDrznWlH4ytwyQtjPOqlcyxRy3C2gZeLyYe1ISGC9R
AuHJoVniNCAq+8Jc/r/rX9VMjJ4mwUGSBURuqGXE1+fKHl6Mdrq6vGoGVcKY6OczNigiWNjbWVmW
fbVlFFna2/9qJ1Xw9c7tDOB5NypJq6W3JKn3OQdtVlwTYjUpPImDeyaRH8VoyZJmvx9Ws2Isy2q6
wH09NkGc3aV5QPT4SHhPC0XKRrf/30A2RQzK9Co0lJNXUx/1BAtBtmbqyrKPb1L5YBhgfAEVDULy
poGh8ObBX0u1cdlchtrtAEJhVf87luyKkwMRhX2105aNa6UvI9LPfBEGnFBThyhZ4idfK+i5f3Ka
sJpuUXu9hl8KW2bFDg4KggDu9cWDYtNRS0up7YUJTDXh0SC12aw49i8PYgZV489t9of3bSSMusMA
pI6OeWo7pf+tP4O9p3xarUNbBI0kDOCgwjUgea5TedgjeO6b7Ub8apk6uwU2I0YWUv8m4l4HKNX6
UbzAdOk9in41yM1hYmLZ7elu43CwxqNWTSiwelSerKKx+K1nBN7oNyEkp1Pm7Ms9XpLG41IlYiGR
Z+jN/vGERfKudSJsQydpR9Xf3S3DPUyzzKSrJpoDlpDBUeixhguDtQkadvxlUiTQHVJxa5TkRgFw
OXok81J2HS2rwdp/1kySNJxorhMgwXK101POhtMye7z6wyrg/doeqHfP36XhfSxYzhdM+7vEc0No
3eELXOuulmAcFUeCesiJu+N6Zmmbl0YZB9GWKz58x1HOHDejj3SX828ziN4s1OsojLAVhUQ8Msu6
113UgPq4xF8yUWMh0my4x/+AbdFAO3qY1bISfwh7Zxlc/uBVG57cj62B31J5NGQDov9gSYUxvN8u
hh9UsttPl8aGefyRgOrGyA480TxJ3/ZxRNayFHQUF0zP8sCKsG6+DKv8QKKnpbbMCdTnBmcce7Ec
W6OIiA2yS6uSjXA1J+OpXjdXz+eZRQ4LdGFdQfsRK0/HYj21rDIYqrBEdhCynZXtPAbUY89QOPLt
6/OJ0bEj0eaQdfdnpUMywj2npGfcjOxhION4ZpdmIzlhtrLUYtbgMUVhqLXyOhgH86RTyd4lEysl
YqHdQrnw7WAoPWzR67yGNHqNKHIuXbYMeT/rIaJ5mtHlyvEa8Ba1mIrJbmTBmMnxyQcoQDZu6Bwr
jwYfYwWR7woM0a53Da4yCGLfkn8/Dvli1TClEY00GyDarsp7dXmL5Gl0Q09fI9dD89OwjtDEaxZR
agwX0rUSim4lCzf9VBXJe41VhJaj1dx11CEeGKGz6V+ucuuNaKcxkO8HjAgrtYjuhsd4vjsWXSpV
rYA7SMeqloy+Qk3x0ViElMVoBZFQEp3AUmsN3NGCFCRwCZA046WKGU0uyzMWVoRXzOdVIbkd2Jft
l2/Ck4aCYTRXyCxqbbdUdPuYfkIUO7Z+nEDLKiCmw+E7uMfOoCdUpxBKbEim80aN+WsbxieF1hkE
78yOFzBTMwVC4Zl9U0ruWukJLw1jTYRuyEACaCPzfLHRMWYEyCV3CTc8P+W1H449sic6ZZbxr3Vb
616ytUmFPKW1WuL8x/1ZkOR/UpkrS1uOYm+79ea8Yr7KQ2W6p3XZlghXRsgtywMH577xkLxrhHcD
zxQ6ss8qrA+bFPR6Wz/y7F/5zkhijtBPl29VEkRIPm++UVb23vSop3v9sRjWdSVihqBRJZZ6j+Lg
EG4u3kexNJ8nCqus6XJxOSWZYBhCyVUiD0700nHrUkoVht/tcRkOYXkWiisNukubNiRuLAv2MDwC
VdsGEpoVgQtGBBlB0Uyg0jhe67zs/g2Z8VnMw1KvgidN7VlGGVm8Q4oziRfzoX3I/VAnF2rb8gm1
qsPV37ak1oEuuWJHk1kjgOxCWad7u75u2PsUnz5y75hDObjrbTZ2lyXwRWVJDR7+PYlCYGW2bBMr
tt/5Ird03au4bEeoYgcx8eA2miqt30Vt6/5lRotpgcBLOKEAWTza4ZFRFWM6z8sH6Qpnm8Lh0Xbx
GdGqP2T0JO1+/00lwhPg9PIQMif46AiMVdhGcJi8FdQm0KpMZcbTCFSxCsN1KITt+MOErVAExVHm
tc0NSdbiHrms0rLT4Y6aQsjWi5xaGqYJVpAFnmboSHST47ZxRoOpaht9WhE+3BqXAz7gr+RmfCp7
ChYTFfZUXgG+mqwaqeA7C1lF8YznYtuy4RHzCKpqNBY0saFrPdGbq/15c0xrBJ6CvaUADmxdebaX
CldoJPCAXDiNtbRFSqAMk9jja6JOTOfN9FLWESbE1Xd0FMGMCJwmvYmyK1DzcBefswYaFy+dwPmh
gJMbqP2/iRlBL0vbADOaKte5oyP7suWUvkmDzhtOp0P32HPoFi6r5it8tokT+W478eCQN+BHb8X+
ESK9dLm2Cgcxvlox2NZkoOY2RZPBKfXHwv5xH+FdPxyynyEau8frKoZpdrIh+EShNb7B95aZRZGM
UOpTUGHzUQ7Wetj0tgEC4TV2cWcBt7DXYb00i+lE9UtpILBARUTHCI2oTcShzqqMTNsfHbjlNs0A
remvO1Ot5eMxLS8vYroe5ETCRuIl7aG+wWo2bvINcUPUV0Ql2I5HEnXy/Gx+sZ0ZR/4AN0VPrTgp
1dfWnFyF9nlgZt70Wb4CyvLL0+HVGGvpBrn6bJADr1H8SUl9NBNKjpIWcFI/zeUPp7RSVuORGpPX
U9azyq6aTPYQXMV6DTvVYH+r/kXVJ8TeFHeODKDwlRRWfQ9IkcqaJ+Gti7IdIU5Yi4WdApv9QSHO
KqNUAc2wVopqz02MQm0+Cudud3jbHbHIczCKOalWy5ANEP5vGNbKZSNVF393/ScITeLSl2CLCtDR
gWIOHYCjC3HrHhcKP2JehpkycO6OiDG75/GQsJXEr49moRMqlgMQAGAlmWiBENL6XaxaBUaFZ0Gm
yqFP1mtuh0Rtx4/xCI85LTAz2V8jq8C9Da/SaCwZgma8J5FEygZj5YAaQHQMZuTglke2E8c9tBUm
vJEzpHZ/7lVLgakh8//9KLnRak8sAufIadQYqMYS4AzP0VmagHpJ2uTxEsN3a+Q1ChpfkR1E9S+g
LohlQocteWPOqvyneCujEI+BJDcTA7e+I39Kjgc8DobCUMG+CetsYxet3Q/G0QesgW+0oBxcAz7A
Z7/IGD0SR4xkPNDcIm0vbf7G0qNtB7IOu3ldWRYhFNZfpCKDP7rC+QmOyRrowWkXzgcw1HHJbxi+
TX7i08FLRROf2wh5p7KC/Q7CJNGasc2faRknEjJKyM4uffu/P4gYxQ17bRlyIO/a+XOMG+YbPp+b
KaGmvOLIZ9BSta+/KajmgsIcHn3riPxo37Ou4a/e848WYRN+lWKhQuM2xqdXfMrBUP+3P+ilvGcY
FcG7IiA+WyPsO7Q/dRWCcC4A1DS/aro51a5kB5vkXG9N86p5ue1nuGLaoB/Zsk7qZLy5SwUGgSmK
/a5ZloxaN6XawEEA4AR5Xdc+MEwpZx9kfBj6/KRuiKPkFUBY4rsfloH7oh0u6fQ8XTfb6gAWf+sT
AoxoWW1k4xI1lgkJJZ12B8Sf5OGc6DUT/FdXdyzvuO+aYqQ5fq74LRJkph/svhihvx9dCkyHPp89
YJ3JnbwFFDwp+jzKZfe7/1seCPAuBYtAirpDFdji/r7Y2y21KcTroZHUrIe10rwCKqaSx4mBJokr
+L3vUug6D2qcCwA3xWLj1EVp+H/GuoGM/SBVpBMwXrzH+DI/Qee2IJbshsFm9UFehP3eSceeuzMb
m+s+MtxSlDJZOngM2470UvnZ8pvGhWIya37GczZ4FtSOgbYL5aCz0xuNMOfCKi7U8r0Vbf0fRI/g
BnZ5txWhNOHB1H+vWs+Hf8WMaTKrCgPeFCpXutr9G1zcpwc9FNIjGVjKZ7EMUPofK1ke9jTNZ1va
Kak33XxfEMlcgwsf4IMvqHnAoQx1VOGc0jzFE1Nd4SL56t4rWdNMl0Jhe7NY2G5ZfCubJZ4MZpNf
BFt7TuoF/H7CsQMDrSjWyNZjxgcF/sl1RXbrrPD8108EDcqi6HC5jnYf8YVfmfGEnpXG40fGQi+7
XExemVITmkbiT1Hdkq4jVpST50bwn/2cgqIOfCMcGB//cfgd9JVGCG/iL3R+AIHegHoyEORlO2/S
zrP3fhMPjRUvosY5bbAnwMx6oOamU8aSD64URfPzZvS+ZSFPpBPibw/yw06h/U1G5nAW9WW+Gxxa
qkU8spVsqvWGVTiaVL1683/dl38CEo4Cxxml+GhMMtsKsXp+AnhSzjYiNjSzbP+kowPPzA1i0JZg
EFyrN7XPYwITjAyTthiITl7iWRiyJ5yjcJm+4NV2uGCuV7UMCrWRbm8dHYvaeE9UYFiHzykYzh5S
NhgLtCjrBt7fJL93hryQR7W2meC3U4FiwnVEQCyUuAjv76SxsKi4NgWOmRKO1YYa5GVhwxtJx2fs
KggYt6wLITVLhh7fAdXeWQ4JraJEjDQIcxrTiog/GIqvddbu+JHea1PsybEiDMAPdVuNpUmrdSfO
CSU+w8EdyC0YpUMD2CNq4F4Q604zrEVHwx+yjZnHA47ksNrSurxRnRxs2klSnpVjxrLNIt4JhyP3
21Z94JUlrIVK6yKMgvN9m32M7BmkmpuGfipbp12ReYDZWfG3ggPKluk3B28XyQZjbugJZeNFjQWi
ZoseshG2kX80f+TlSCHQD48NF8Anjwa4R+Wv5BN/Vg1x2jSTwO+7juch82FyWSY3CM62A4S+nr0B
6wu1FCJrWkKb6ZyQxFsM0robrv2k6xaMHjKlgjzjzMJDOi5NrMnkEcguPOXsqd0Wufcfp509hGK9
fBqeyg/kNPZsCXH8mW0NOgTV+Sgrubj8JD156y2bglTeguMkZiIPGwAjma8N4MuSQ2h8eOMGnbdb
yIuP/1nOWjM2s5/aRZXXz5vF5NHXHCGjEPBQ9K3jGqy0I7uqe2x6o9TURkBKZgduWs7EiQ2PHWpZ
uTp+YNGPBiEd4yyTKDlhGaS3y7KK0xpDuA0YcR9N+2Sw5+1rssfRB3meWXHI04EcPjMT+vZOAZtE
hSSnAX9cArC1D/1HNSvVvErFLxTaSCXIkpYdp3xY6hp0FYr5eLg0qleU2spTG71H4xBMzJH/fd8k
tTcFGvvod1hzUXXuYLg7EbzlD0BSWMezRypsvWNu/YxxBh/4woNTaDvFCezKL0Ft6Cqp3lwtmpI3
/YlIJxk5nfrB8FA+W/7QtSmomkUP9sFgSHRtwFEimvQzd3pmvjbRXNMjJMdES6hz3jyJHepMk+kS
JHWBqxyf1V8cuGFPqklnS6RvwNgo2F0BqDttuCOcdK5JQl4I1ARTYavr4g133PSq82ubAno2fbqq
RTi11+T3pypjxRIzAT+4FZ4cY7NT3ENKE6Qs6uF4csw8uFFHcqG2nOTp4fvGXmq0EnPFLc7BRiA3
Gtxcj7NOUA5F6Xx/96PWz3tJM6rnF3aDb0uVGkqfXiASrropbKk6USB3ObBPV25k7osK9fZKyYrn
Gc1X1MAQPlIGnP9hyfIW1dtetEAjm0uMoaPJ6bjJ1f9TmLEiv9mwnGYJu4VeUegBX51o2U0boiq9
GoKn1IhBA9vJ0zdiO92X7zlbn7vyBw2/OQ2mH0Uk0KzPNxCg8ojQ1C2ZH80ib6dJ9+WVWZntsE22
lnPJM1y0ykZm5ELd1S6VEDoPvciGuuTgSsEWNru5KpFNDkWt8Khe55GeL5wDN0MwLUpvd7y/CB2B
4JKGIr0sfddidz7+uu1bv2dqJIRxZtjUA+p5RoIoSq25Bys2ZWAkuPd+uvKRKPcjQZeGXy5sqRZX
x5945nEJRkhAbVFNrwYGmNhjNKvSvPWNFVj5tQEhNyPBOj2oT5qlqoldQM5YG89rrPdfdc03c4Nx
gCgP/gMn6joR7xZvxyqyLOwtehLcRPA1oxH6DkmzoPVmGK3OXsvHx5UXO+iNjmwpJTPPpAZT80Ec
GL5PebAR5udhKQXR9GTZDE6Lt5fd/WcbK3uk2emZAysuQXueoXhf3zZPGZ5IXrOGq6CPGhIcrMLa
HS7LXLxrBHKOZjyAcfGgYH4SL0oDEp5hS77IRCcHvfcQtog+N1nsDru0/EqT45fDXVUPWFCu0AZe
wS4X8MUSXeY3ZkdT01wfu8lTCO7NGdH6Qg1FeZdRZbFDqWvQIL2/aEvevmNFSqiock9Ps+ml+N7t
rH0JCqkqWC8lqvbE2yL2juHoKkxEDStWcThrJB0UEddAhfufKHHXf9gCVCn6Pnt2ZbWFmdnQLX/l
stC1LnKiYoaIuR1LJO5bUeA9bRVfim1BWMxaw+3zHdjPvi2iEqcaPNLc/Fquprg7XghivW+UNMfp
9H4MnMpwB1B/NDPX2FpbAbO3slydYBagXm+I4du9v4jatjuc/iB4ClOglLC0ilbR7xWjHUhUOU/V
93CbcSzqoKgLnu1ixUrsxPElOtjlj6URldLjw4gzCkJ6EIGsSdamd2wsVkLdlOzgB/zEVCf1YLbO
xQaNNl0VdsoGm8cnrJhHbA2C/sLa7JPKZxrO0YV/X+3G5vm/kSMoogSR1wjTNbXRnubSB2GZDZIB
8FI3m/LlXNuvorOx9PJ5roVszBlE23Ocg6qGjRzi0q4ua89IFBo6FuAeCT1AFdl8iF21k6FVpx6p
B0hb8LIzVC59awrxWML+pmhY64mXUbAIYQ6Ws33uFIxuBSnq23HJNWyRaphmdS6nr99FkDp6l1kV
ehXzvY9GzvowRBtgx5c+gB0zg01xTKJ4WRMNcdv5DyRDrWA9qvPwUzmvHcxfzK1J5XvL+8tqVHPn
qX05Dlkk45fuh55u3gmXjV47UxUKCn+vdP25Z2LMhUiawmer1xo2DpCIYzKhkuJNEY7xB27JBxRM
pyHG2xflcQUxIi706e4KQ+QqnlQ0BLRlmQPZknqu93ABT1dDzurQdBkyGE6lZhSk9v+inPS+JZER
3CN6aVlkJ+j7xKPFkL1zYG1PEgu9F/2cw3qC0ReifM+yltVt7WOguqMTGYcWUMMMmfcT3pi1d7QX
N3RrkIBcL9eeF3crJa25BonWrK3DClNWJhHGahbbZCeBkaQN/gUot/HSXsiBLOTr4KKpuBNPVvbf
7T0t3wtBA05vhmNZvz96OfjIGYQ2oDFrt56wY8MyBmemNAW9w9SnvGGF/H4Kj2PJpgXnIhgf+sfK
bMwNmS8fAvfX8JkG8arNM9lCXs9ya1OvCnD9H/gXSIl205INapdwb47thQTIihpvE7Bf8WM9dZ31
hvuakxsak+o9+S4naqTQ3bhBk9Ujpw/BdLUGOR/8YRV/DROBIh8f3YWx7zTHUXzbyYXPmjko8Khc
thw+CkyA1I1q4Zj/UzGeajCzdrcOS3KTwLvgf8m5Llj4pT2KenlwdIOdkRRH5l//KZJ0HrcnLGYg
ltCg7ZxkYyvTY4wnWaywwlZW6G0Uol446ZsU0I5pe5STH9Y4JAX8aNC2Cc22KhVWeoKVpvADe4JZ
9R82ewcX1xdR1hc0ncJPBvTiw6lShmI4dWU2pUR/Gu1NvSlUt/+oycEfUwGPSCUaAoM7LdfE+f4F
Qo91ZbSLFOdEBR4mQOp8O79Jj8Gn1AKt/wDNie/RB8b9GFKLmsu2j/U44Cwn+41t259qdCg2q28Y
a1f0dboHAjxAECXmc9h7UHDbGUMnxfM+KtWXh/pC28lfwlAkIfTTsq3NBe3PKSGSHGIb7W2WqOS7
Fj8i5DdL0Rw83UE2qSxjCpDRoCSqpBhKJewQIwe35Iz2ViS6aBERNGlyooSKScxb2uZRDNbZYIhn
zmuJvy1CXrg2hUTUJfpig2wk4lP5tm0HDzHA8xT32nvRjrc145yb85XvIZ25+roUG764NRAOiCtv
fFByfdj/xgzckE3dSUwfzHdpn+/vpGlZrGNPK4axvu2VP3vFZsW+TaB47bqG3x+TVy7aGYD1FbvS
qj5GfsI8f6UzCtTp3dvUgPgZDXcj9OTIlW9iA4f/NDtbVbGTw2dBwr6zuzkSqX/ShhwjMJ8HpZFR
OxIfIrI6W9eZX3yvMbmSfeiI7dto+po6SrltL43hmTq9yvriJARKHTGuZwzbbgyofSdXo/xTTWm3
jSQZb0lTS27avCX6D1CesUDJBHBpG/M22fjUEeO9TErcTa+rLjkWzACjIs/1IvHyl+mkCobgYGPZ
PwbgD3ZD1A9fk6UQCGKVZVg8eIPGYVCbZ1seniKfyONqCgyu0Q1HdsCY8pzciackO+tqvWwwbh2e
k/g+KGUmtYpLD+UIF46tG78kGv1rVQz1TJKG1KCt1r9Eob8zov75rWRaTHH6kaBzBcQmlse9HVWm
gqGUri0mMT5JfVjkSblzld5TPHXc+Tds5KJ3dpWmFRo/oa7YH9gzAybpAbb/oQ/7mHOBlWCoR7og
nTPm/DBKKSNMqtsoMFDTc4UZ/3lWx3k+/VDXlhA4iHwEdcrla91JFRet02CwZF6bZHiNmacW2NKZ
K3iffewZhBUoCJgLISqyN/yVoEeS8mvAzRFV9dshdL5nweIRsg/6f/NSX3uDVdJQT238u4GyAu86
x+aEmd3zB+EsXOF0DgM4fLXpGOq5ml122VLIxuT5q5OILcpMY4l4iMssa89IBQsPcjl5PCS9aURR
I62ftu0T5bb5lYjaBbWayGRS8ceFj4r3a6K4knu/LlHTrY/kprN0lkd6YLGBZYqPvJbQs3HMJNxg
HNQhnMd04+pA6bzPMr60YXGNLD63vUeG6dl1F/hDmR4z3R0LGAeYzwquCIlqXQ79qUuxGVESUp6R
r5vl617Sj7qPt+2cHTkvPHRmqQdfc6SoHxwrLyEEIBp87ClbO6i1VbFQrAmXUiyrPKBIsoSYlP3G
rxFjpyma779ymMuKO34CQ5qconSYPUMKn3SGes41sARiEvfIj/nMSb+mL81BvFFRzy+N0ifV4eXd
1nk6zswGnjjss788zxdIrYOSrxJLmjirG/Qv0d/DL4Z0F00mt/nsb/L/YrmQEzfho/VGsK+RaL+9
UE1X58ZNb9ZXjMVxOFGR9tTL/MtenAs2qYkFQ9o+O32ceWtVHZ+0AxqCK4j+wfLEj12Tl/+Iq7GO
VmvYqGqgVi78eytFsd0h5o8WTN7098PznZ5J/uK9fRlsz7KDJh6Ti1K+oKIo4QHxc3XTWwrcuJ4c
2FcCYFUkHvWUtwKp/eB1BmsE+Z+2TT05H4GKLDHnc46qoptbGEF1m33szZOpm8Dl0imIqWO2z8Y+
3cHyzhkB67DBwfKFuxTRHYtJpPp5IvK96E0txDnMq4PLSfoGs8bl1eKyJst5w3RN6huiadi7Od4L
+b9kRNGtTLzDq4nY5uvEqbNPUwk/2IlYy3EXJYlw50myDAszsVqDvQ3mY214EB6FD+b7ZmRGjtmQ
R78lezLmvFdhfgv1OhIiMooFdli2wqvRa2GBuOurXU3BinaKXPAVINMPgEv6D0Oirjvzrk87nSaD
OJPnjh1T7Ven79S5poCDiERHSEYkaMIuXlzqIsze7H81zun/zxy2Ku++Ou2DjOGiHn1pTrILUlbw
NA+/zqBiwza6NZYXx0gFDGhtg3lZ3byUgJ3oAcqJpd3YfqgAvGIZtkG+/IJ8gfGkq2lHJqZX6v8A
sWpR531MuR0WFMWo3VaGbDAdSs00mW9RNMMHppsCrzNx2jO/MHdM4jHuwWFBwXaDXlcl1naDy5d3
3C1kuQyU2Q4cBRO08l6n6RL/c6cyYaCctL/YyLGMndYS4GnSj8FTMt4jrhKrcRe4/mBwalZLLZFi
ATwscXFS/mnUYvA2leG6qawX3Aao9WdyBieEVusO1vAMR6NiQzOvy43yTIVocGZRSEqI0ew4rxEH
WfKc9nWx3BRBA1dZZKBipQ50K5o28efzOOFoHsokSAzNIKSNDTYl38KpYpfGXoH1H+DdFT46Oy79
ieay/0UwDrhlPl718Lkd+1X3n9eqFQIzkP2zu7Rjy5IiMvb6yogxHow9jsJjZ3tCXB9X2AC5T3w8
KIovEIieQ5Q79kPUnSxcKRYygflqcT/C4QloiY3H3FlABWzK+owpFQhISvjlTsNhksK1Db7hwknS
oW5/7HvMWIswhPXv9OqCy6Q03q4rGtXUZlLyYCo77fISzfcYkeDGB04sHN5K6bhW45m7Bs+BBxsq
Q50hi+DQ+FYfH/IRIcfe/cYVoNOxsNBNl61ZDMXGISCz5a3DBLDfjVnK5CmhzBJwCCFd0hgVVfAJ
UtXzt62CkH8PL4aAJhxU9zxJvdGh1jqKBYGcxHx2TlFvOLlgldhS2LZCXDrbJEMeNo4FKR14DF5D
64xGSr6XE9ZeUyCQchXy9bkb3YXWJfSNGW9yRWCo08xE/WgBEFYkDNMiSNEQKX2OiQHK0yWSKjE1
wfngYsmj6Y6WetbO8GRCba7de6rMU8i6/MwpIqn/Ne6Z8ZtIFoDu3I1Q6/zX3cKQnosPqsusnRsJ
V5iau5a00TT85+6K2sBViKbgMH3eNEgPmhVr07NjPMD1fMo8RYX9UFRVoGMJrSWoTWKk7B+wluEQ
hrg95CgEkXwqzpDJDoyY6YX2C/2NyjHuY/a/4ilZxpWcPtlHuzlFlwJHDNgiRrr1y4icdkACDfkc
6w7EiHu4kI1bqdP1GWrlS8H+TLcB1I6Ux41PY+D5L466qJmj9bs3Kc9nFLSi9A0LDAHrIyJd16en
tzKQa60zsik3IHKufkdb5cgU6hlXzc9cDKf5AjucewwrKmonKmK4VlQSpusQEwHSRvKa4zqbE4l5
wzQgN0/PrqTvqSSw6Obfqc70+m3YVUYVqLnhyDtXsYsr+Ljcc0DD3kq2vLwm3kz7av/3muUKwylK
hpe++H26Y659fCEioDjfZ5qh8JAUUui2TLrwvjg4FoXjFSe7FVXjUrHiOiOqcj2LrXyv0vv2ycbE
qlNsYCjLEOx+Ec9dqalYxycdTScdbZXCmbQledGCnd66jObBc8euI3YfvqlprKzcHgqqxNTMiQFw
eL7MUPRvNAulkXyrcnyMfy7VucaCJS70jEzdZ7fOEucWA8vrp1AE6kEygPUnXesL9Wr3KXKc0SyW
mTqejE0J8oJKKyhhk6gjcdXJHUGEhFTPNw7XYu6AWarqSW8RErw17LwVzgsbQUccZuXXXduIapNu
oNIAFRyRiBEXyHsjifcHVM564WqeQxVe1EDr0bfHCHObaYWn0ruuSr7XL9x7Icq4wbpx/7zuCOfE
Mva8jzBYpVL0CbvmCwon9KQ6ojqNAa6JiQnTSwgyRfHC56hvY8cH9hGIs6s68HLVJDH/VtO/HuCQ
ie79Yrf1oWQGolVihboQ9VqbKcbKyWrQaDExVgEp7I/VPpf5PgfsGzrLnIH2aVIaxASP2WslSDqq
+C3wXZrXTbEwvgOz3ckeb0x3h4B0OkvQzVJAQlNBtoE718X8VnrDBk2x8zqKPiPu1CR78hM+8BoF
VO1feL5w0hhzpBCAri1f99qSgMHrbyOHG4gdv42ivoZXdiqa4yR+/vM2wggVrNYk6CnRklQFD1lx
W2361IEz/Eif1RSqrtolBRVpLUaCkqt98nP08XDWILGfZPtBLL3xl0rIwMGAn2aNab8APGlrY9An
f3l6p2B9gj/sOUAKYrEmiDEQJ7XQJ4SFVgeTI7vh6MbizHT6qMn+e+DQXxK6bgvMoe/CWAPRBsn0
v+5b99Fyqlkd3y2QwcIO/EosWZXcrmz30ivzmfH+QAHg314Ontyo2FptZL8474boBERanK8h5wuk
4/MQ3kh3wabZOYWVkpEeNOPoDXqoz4VRTB72xhOPf3G7ax9S/+W5fn5e5p/TI2wJeaY0f9UwjbHv
whoCWcNEVqEfMTbF9mCQyBSrgiyVz92IF3hvrc2/wauBUFCnLcAeZwDXow/dmcX1BI/BjnSZkls9
Kmia1dXGQXjZH1rJx+6sQal9Yd0n5mHxW9BmC08IPP2000o7k/R/j1sDcU6yODJWsdDthNh16+ql
nMiTIL/bk1BN+ALghKFDu4o8Pie3s98QOga/oIclx3c8uCfxXsub6sQoLPaGhjDcf8Cm6RfkawEw
Rw12XY/MOJxd2rC8vdkYVDwU98ukT28D3hIA/FkyPYVBPuR6sudU5MLJYbdNADdntf1JQkMgalB8
Dak50yQ1Wk/ByiYZfjVDlQCOGG3RPnIv8cZLCWoxK5+6fR+w8D8xPlIthFVdB93y9eVcrvr11cvz
k/f6S0a/wfIXG4QjmkSQGuNRoFst/uf49/2j8aQq/NHtduCGjLERNOD0DYj+v5zH/ebt8afxrWq+
93N9xLX2x1Lj3K76EMne0ozoSagzuaCkuTn3R3go37F7Q2b3VTe9IS4b8ImPCiX/BL3vGUh0ezsg
uW81wTDhJ1Tu4nbBRKxyBCZdSM3PcXqgIwux2i2Eti3UrjIUhZpz0mZts9Dww7T04gikEcWV024L
kDNTtdlXwfvU1qADX85j1kapJZ8pUTGoOVkutpsqyyaNZzNQe+aQCsfqikuGXdnUFxm+wHnthZCm
QPdHBpt1+fJuev6HXSF4xf2PXs9pNfZ5UuIXCjsZnmbZ/VYWM+a24W9xcJj696lUQh8lunFMSpFL
4kXajJsxCXcpI6iAV2j5bmU21E2JLcyexkevCg6IRUfPPpXSt4OPtiW1rEEUC/Kr5KuebpSQKEpn
J7nZxTwVoIHD9AWerFH9/qEqpehmaVF3zBNsI4R1LBgcV8c6AZRjxdSmWQpcw68aXCKAyGrBqRM6
rwjWyZZtPl1dopZEU7ai0jvq67hdxnpB5cjUrDRAE9kjFJl8O2j4jM/CnxOf1MnAmiORiNMv+sJM
tvXI3aT3kG5WMcdegKscXVZE+n9JM1YhdswfUBpWPrPclK48qGk9Y91T/abn/CG6HnYnRtDkXPmo
8x8p0zlScQPRy4dLsHqIn7qOfiS7096pwBLDSM9B+ckieF5K1Jui/uJvn3h6K6uqtVyA+b7cxrcq
HgEFk8FrbuA59zl+enQ/u7EmwzJ3Nwn3iJt8uR+RFYwkF1CaQiG9dLYtWCIdAMECRBvemSGLvlOO
ISm2hdY1VlkmLOhHU9Pmncpc7HzW5+y5IIPkCi4ccStFgs3sbKhTYexSbM9lYGo5HmSTwb/5m6Rr
+ibwkkLPFb+hWj9u05pKkvvyynizLuMVb45629WxuSAQF9OYes0blHvOzkz6Di5Gz3kn48REEIEo
oPPemRRqA8U2flx6B4D3P4XHWTvCKyTeJ6bVOnTbSTSgvKq7tDbzmnHVNwCbLhabo8WS6zjPrBSJ
hLad4c+DjBcqtxJsBTAAXRSXvuc7qLhwIrdxemvLR8ml6/aosBt7C9u+PpH44V18LsqiP/O3Ckw6
3nt/4f2SJHE5MQRERWFbY1ypcPDCkEbO7jdtVbAK1W+LYhTrtnhbd4lv0M8PNvTNMcvAv+QFjmYI
cFie/cqsd2jtqS//uSKWV+vLbSqPlrRNgN7JG0F7y7DQQOkb/7pAW24bJ3XzWGnAPftIKUfzXduJ
iqKPzqfCheSWSiMmxgtxXjjfluzVd3SB25GmqbKIShgeog2bPNUVJaQ4gpf/etcvGiN7RNlO1OuP
QblV//XoHhtJrmdvktyhDbjNryqnWg0Xatw9DrGJPwEu9TXxRTjQbR4CwmuS+FcJWtQaaxJ2qm3T
lZXG9tdUEnzth087G2zIShscQu+ejORv+oQQVxkjBqgzT7EgiIYj3V4DJ1PYIH2Tehrq+EsGZUxb
cAmVYDX3FWUwpNaM8gK2Pgp2GgN6/65LxH3M4BbuckIBYdcRHpMLrdwvuuAjd7uNsuqHN+axl1Ux
n6wPYNxqEKA1K6OYNZDsrBjYUQ3Gfd2/t13eYrIHGawGUCvOP3pz6CpwhtJl+1esXCLrUBLqjOLN
HYPbp1kSR9IpsW5fXS4XyLXyrARRKFd+hVVCaA1YyoccJ/6fkPWME+XQuXKB5H4x3cA22+rrce/+
h2p4GiJfGemKEaO+FqjJs60nrejj5XDOHZP2el8pUSdWNCeDHK+MNsZ0A5a6gA/TE1wF4hCLluOG
AsEqIRc/Iu22BlupMHu947aQmQTpTaMJE3Kqb5ejV/+Glc4m+jcxOAsAiBbuGtDYeDEVg1lpxDSp
usDuV6j7jFHiFKjrwh5e0r3g67oRul11cZ73EcISmlGT38OODjAUBDXE1UHGgHKjTwGJzabrW+j/
LXn7AJgkGK4/JC7Z6sPABPUm9UcJSMKUOCH2MMoDdM419TYCCydpS757M5GyTp2Uk0hU6H/WHkFN
I64VIzMcWh41dmLX6qVoKBk+dk/w4r/+jmZ2hjI93+jVk4is618KPHc2uuZT4ChiP+pkO9P1wGsM
ABLXUwfHk5fFKUdv7AJB0suH9qEEt0jMYWJkTWwmF36OYl8LENAVjDlK3bedGGhMUumwH3PmtN/3
nvOEGR/SEH/NnHmjIS6KuGNC19EI4UYfdIgZrCLjMECR7QrjirJN6wJ0ozkB7jNv36Sm0EEAB2u3
jKPsjl8zB7OOaNPofOXGj32ghm8YzsV/FkjvEK4Nrfn59lDBeT2ZyLK0qDDlkioWer7oHBNY1iLj
0F/ZacEGcEwgohirzkbIrix8817YhVgJPAvtTpu1cg9xQLQ/4gvGzP1Pekiy8MfsJUqTNyWFeC7L
t0B/8TALephP9SaP9GdjfC3udGh9ALhGQW3VjxWm9Y1sYWaqGT06cfTTh6+E7rOd8ElBPNuJqMvF
xWepdX7LUzh0in1ndP+Hk2K6GhgCAVhGF12UO6UDOfxR4gMX2ls8/UsSr0NRCglXWhZPnQ9+645k
fUisxzs5+CXDfUuMRIHKPtE3/8fmeTMEwaBLiDfGHGyXjDk+WCfOXevvB2LrE2pflH1DIzZ0Bm7D
c2rTs2rAJYz2QQttrvxfYewd2RHTQc3NpcTU/BqGzwsg8cJevakaZ3vKSQhwn38DsDwNo5F65LPc
sXJzX7LUpcNp9+tc7QyQR7FmQglU5kEF+cLTJnvd4ra5pGRzqUq1f+RbdhWi1sIqPpx0IcF1yfEf
uRwLSlErjlce+9RiPtq1HB1XsvdL3maBsPd5/el6h/z7JwA+iaBBgBoerZDQC4iNFy1FdWdQZJhW
ElRmiM8dBV80fOpkP0QfVVCRHzVyR5MIsFzKTkePwQphczaCioEpdAiphDJ1qGdJ0TkyZ503XOXE
fS8iLZCsiFcuSQmO3dcaDoA0nsIrC0vpBh1hlY9hqj76cI08ufU7eqYUi9TqBfxVN0QvhtoecJos
6OUxmt2am6aHoN2AoiadCYScpKOUpsZfUT0TePJatZ5MEr7urcVEEp+ZGBb6BUo7LeF7+DH//awK
jRweaErIIsopzC7vLDm0ZPQ48QgDDaD+FDyV9k45R7VRoB7c30eqcB+BnN+gwIWfdFwqXoYLyrB5
gIy6ydTeOUeDkUbZz3v7L3yzEEcKu8PIXCJ1fN6svNTfU6B7q+KH73gIsJ6/Qwl+8S7AhRW+FNMQ
BtoVPIb4UDppxVdFOLGcpYv3Icfz8Cg6dTjjPTvr1NSGij0wDAALIN821BAtzo7OSo05yGGVD1GP
a/VLSdmMEDqSk3ZGVwmTfzaZhxPOB+/1HuR8f4be1LklbiQAQiV2t2KzxJ1v0F3uDO6Iho8pYewE
X/LdnJl1epCpAskXNtqLDc91cUyRTeTR6HS+WbWvh+9f7cIQhGdGJTM/N7WpgHAzjYb8TVraIR1v
wFhHfTuLkw1KNfjksynSbDSpE34f2a0J6aE9E0Ji6mipeo3eN4U0ufL4HkcXEI8eXShR4f4lOMpE
p6mYLp3n2n7bN31xuELkJGJAawDR8yYEM/qBw9XniyDBtl/ZqgXxXgdewMmyIfuCU5Z0X+SJegO3
WSJ1hebTJjjgusoM/Ma7eXNygGOlM48/ANfG3xnMput4EpzXFEZflLVHRl6yzGRAe+Qu/boz3jp1
n48qKpooGBszTewNQGAgCcjqm3PQklk3ZPIRj3EfPf9heq03zTz//1jBS+oaTtrNvYJPrBostJBR
qTamp7Y2Uo3iclCSRw5C0p3arhTEzDoxsXUR+eU5du7rDDXL+FaqnqvpistnQswv6WRlCJaimZ9T
bMvcjHZ21B9x7+8wKAdtAxlWZ4IoQHsGzlj45/tp66VbwgP7WkjGLVtdf+Vmhr9BnO6acquuSkWH
FaSKg+JIn0P2z4Fin2rR8W6vqSGHipLmX7/pBixDkIs8NBofx2j0UuaZun2GQieb2hH2KjUEiJGN
grkZncuL7gJLEgkaU+LK9bh59JskI0LNrlFlQ0O6gtBw+IFo2lkCRtyr4r+/Tiki4eJYwtEe08Id
jaT/X4AK1zCXL2eXBp0siUl9Kt9bcW1TyGgzZctGi7onW3vWNqpGoGnvQnZ9HbGkFiwukYvnpP3g
aB7a1liM4tUc7qgno+aahDqXxq+YWxaCjXlKrcWGJS7D59Om2CXWNKesxoRmqajeY89T3e7wovqP
LB5rqg1HgCW1SZF7/P+Nvq3GJIbKTnW/XHNJZaPlkRvcqOUQ8fOCTA7WNCIEybh5VcjFsFBLUZrn
vvMx6FhbsFHW2givtZM5bvc8gMHwu9AKtRuEsr1WYKAr6bxSUIK/f7r8keDqfVoeKNbjU9x51VTw
VUp61Hrs7Uqw1tYkpTLumtLtzn157QXErvsHVMknwvTcfsxBTJTH+N0O2ifOdnd04KdZRJTwEocU
kbXOVlgkHpllm4G8IOsyjm2ZGpGiwJGAVJOKLul4AasGY71DvjBq8ia1HWB3hpiY5cMWvG9Cy04u
DmBdsM349RwkCp/PtV4WIkL3ZvBvqSueMihTFrb+GpKqCXyOrmBtQMEX/lOT6yct6HvCzZqq5MZV
BXadZtTIoKogEguSy20oTlE+rL9ESsmiYHQ3OzTp2KkqK36+uweoHSI1H9SrA+aHCBiOHxHo3MIW
qGmnIbGTHmQ3WEInZuEj1qOpZ5urb4s0xyeOaZcTQFQkWqVx17cQ9ECsivTzpXFVNjsUeE1EcLKX
9w8hLM7QU1ED8D7BuMZyBbDd2xc51XNqNdZkVrAV3Yw0fgslkmWEeXxqhsCHh++CEfbuqQa2HaOC
PIAa8FotSnCvcb6/scntp5evtwbrgWn7TXr9sXAEC9dfvo05B7PyXSGaHL/JcJAcKNGQlWzYOS4T
1F4oggKBOiy2S2C3Cfh/i+u0yNmH6vNK+d5q/FcygpKt52o5vqv0JGKtRcrkl67oajdgpc0EpGH4
UXkE2/wEd9aTIsXEyheH+GDTgGLxImaLUZe4RoL7vpNlP5TZuayuKOum3uSA1IexIES/W/Rt9hTs
+msaOM/C9S0u+fztXcHdL8gHyDHsZzx/kEyV/O5xJN+18tbQsczqXtJHvY4VIxrmCXfX8gkwkyx7
+YSMY1ppnq0CzLPYPBWYH/XkHnGuyHUS9i/eJpgZJ6TGYDiPlU4xI4XOZsdc6DgtZ0UDbio8pqK/
g1sbkg2yoJv48Nb8LTpHkfA32QDN4TQQCahDAroEHH7CH2lDySoRWME8WQ9cY9jPVb+VbeS45AGq
DgOqC/Zd6fbOrh74ywujHtEZeC9WRGPgDfMwmbze7fca8cGHxCvrTUikzCFmt3YGoeTmMlq8R3Dy
ytH24DSjHQrN9NoIXNr8Y8GmgOPp5QbIQWPlqcqV46kg1ppOEmgPlnW4R2/TMCmRWKmCNTfy+o3l
EC9HkrHcMtVI5sW+lzYaNZtbfatK4xiBwEG/5j9z5mEDZltU7f19h04cqj4dpSIcV/HuPvLEhdnV
Oin8hoNGjhlhUHLfcjGTy12tQF8elasn6xAMtdlyi5J6yW2Boqt3jjDNF6Hie/U3dvjRuf3N+ebz
DQyVzhGfjfXKELb6jJ7vhGwR3XMcQfkp1iBgtZNdsJPIMzteX8RwYKzhe9gVC3ifFXRGY2tPJVYB
Q1aNxcky4niA7yzDgdFgOhCRcj9F5p69mVW5PQJEnfzGDr23zYppakujpPMJqytmMv+1EBXW3isq
3CaZchtXdDys/JxzvcfVrX0IqsQa659vYbuw1ooY8+ROpK98VkIJ0Itbw9ZHzhVxxNRLqDRJthDQ
LlpoVwVXGpZlw/ZStbsNjTy7hocqVBYc+yDoT6uS4bQ0IP7NtHNjDJ7WBJPXUdp106hg8iDZLF0h
AvCAhzPvwwi2vIQm5D+D9Db6yv0UoTQV0x+78CR1E57swa2MxZkagDE+OvEPVU+pFxYzR3Ygrb9w
87RBtVKQduqf4OC4SBTniS4Hu+ocKtuWMxwK0oyPHnLaPnQSPMBAbLg+7NimSPyaqPeBky00/G19
ssSCJsshCKMS6KfCfSILKXk+hWVXvz4XJMlz0Bsm4fM1ztzPgCz2SIFFsbYAQR2MXZ8TBhRGAPDx
+GxrzTcvPxgLBD0gC+p3rpmdWxvDux+cV1clQPdt+wBpJoUHjGBi/mbQau2kled2GZD8uy21IRhY
+S/WAWojQVDxwjZAoKzq+IKO6Lmhm437+ZruZCJVbVmSGpEz7d2Inc/ZaSBwXW50mi6b0hub5WZA
Mf8b1NNtYoVm+P3U4BVZ8gw1a0KzcDOaOQwcz8Nlll38kCt6+KroLSsVA05oZKgkUaiKjTl87I8h
yzT+hC3X3Qvn9s52MlNJ3GWecGK8XOZRrbYtjSZGVsu0Vc0o6VNf77U4BSqLm7wTrjkcPXSKntls
c9gGeLAy4tOVwMMPldNN+Bl/X94IamXaDuS+JUFCK180hoGwH1AuhHL4RPz0I93yBw5qCxDxvZij
EahzJNh7p1DZ5SJuUQdu1QEQM6CJfVxL5Lkzn0UILdGZHHImhwxSsRo1LN7n0CGAzQo0okKoSOMZ
BAc5/oQyUALlOYKPxUhnex9ytnyykKhLdx8CH1OiKvAClZsda4cUmiHGaaUnPhHRUHN5cryb+COx
bD37gnNj6+k7il6ui/0nngKY4AveE065TGbnfnNQJRnq73qRFDe7wl04JE7734ONim06TNAHwVFD
nUH0izILcJjjGFnojKvmSGpSGIGLUJ3vdxkx0LK3KMa18+QQ97BFvaGdEOJ8W7a1Vsn5mFOQutHI
6QrYpDruYFu6jRwTltRAtgrcbFY9K6w+kRlg0M8U64OskB6Bcdp81AYJ2rcBVo3XMT1xxEgvhCRN
cz4CIoJv8S7NyzFWYN2otmRHWoJxYfUi9gguXpRVlOb3tmCBVPNWvTnExnkZerPx1RWeK3t0bOW9
p+LSkDAPpWwVM+QVJ+PepCHuSWHleTaXcvsOAn7v4/B/z2Pp0VjaobTh5F2XCJS7bS/zAXdtJ55Z
XVwZpsoMGPJ4UAuuRhPIcpgbv0xcMTUdFxXn6pmpfdGGKKRyvyLfjVZ9jWcYR8y1DVChJ1HajCCy
gOMsH9SKXk0RYd05KRmUKCqB2xaajsAH6wohvotgK8puEh1aw7j9fTn+EA9YvtlacYo5Y+6yqlfJ
SGLq0nhIjDZ6pEledz7X1SLV9FlhdAPYjcrJsJKaTmk4wlmporVa8wQa2sZYeZszG1nlYVmtFpsz
vuRRIPdtKNfsrWB8Owse/0F+I8CM8lTYjxRy69d6f9q/V5eSHCzBnBtF9EYDpwY/1UgOFyBa5OEm
W2lXpJygomPud/fLHoS3kl5ulgecUD5ay2s23hSgSf+GwRNeIVvfcRAKrcxZaxd6+iHihAIL5Hje
Ziag/IDHQhiJTCudufgajdv1devoYg6RwFgKFjT6T9xCkqo1etlErjy/YfwFslvfx3N7qzW3qsWM
f5WEeE/jHSiZDXPLBvukHJtC0GukQp3aAEHJTqJBLrknCZul9CG+C444Fn0qBBUPt67l8eZE00R8
HxNrD/zmV6/cFgM8mVDs5AmyWvC66AQymfhhjgGmM3oWyEDiZDNMzTP38fACS3uPAkU9aH0vsigJ
83dSxJjM3h5WkZvYZs3S5mWrD90EdDRxrzuzpYXk+br7G5q95gKYkGxLbDWNerQL6I+97pyv52vu
2twnyuDs5nvmW+PclBje5NHcBl2DY4ec5FiNXGXc2p7KpDmMQv9QpMkcK+wBpvcYHpkfIJX9Wwrr
4AwSOGcnJnNQtOxMOQx4tLZ58KMRc/KRVwocq7xiIgqCXMYiHcLACHMgzJ/fsIi0vvQ+ciRp8jZl
0CeNGv0iwZWf2VVVLyieA9KKCbTFjAkLFUnMO694+I/q2x9XOkyC0teDr6K6cbpxmawncoY3XAzY
OjsW3RQ1jfmDit1Zb2F4ZHexxTg+Y4tF30S7iq3fvNLmnFcAaY/t7BP2sFDwPmJ+rOECdrdYnLxv
tFMhZViZM4bYhVBc+unIrHtoU1BzxfarRfsdgxD/NfM1qpPGsfZIGeYDlRp4/Fa2YhTM7ki9A8rb
WGp1HUWFk5Vb0Ywa4bMqglf5m1E3ZduFeKrW9fNEspi+ZmIJm05T2HVaut6JBlQYYUoaYoNCiPlY
1kCm86nfY5m/NvYDOHl7cfXGsGhRhsRH7ffHxQzhWnCNGwtDuv/JVkI/KsVYBNbq27FMhUNDvGgs
+lzXSz/w+JiSjWSYVjqd7xR8DKvri1iCjTaK+Idj6hGX0jHETpnEpvQj7DctVy96N9kqmcXe1PHP
TjHs87rYnmcv+VhTcqZmi/5dUFkMxbAs4L3WCmHM4pajJpgTgoLb2oocZmMEU4Jr8OFWei6y5/kg
q1IVPa2VM5Qum++ANQf9xoyV38qjoy5otrhIk4hwZmHH3L9glLDSFoHiyOyYhm5kUxR06z5rvmmZ
tTW7wg9Xr4LI0sdkxiefNEfbC7bERGKKOSs02OiokRK98xIBhzZvTv/0MYSypgCEjGtfWj1Jejfi
PRf+13qk6XoZZSx63xRPenmhpNI4J18BsWosDINY38Nh6RPPQiKHpnlLAJN7lUg+/fpWbxVudikR
35d9sI2d1bJ6qB8RrNqIejNjNaiAklqXLLrWhUMHRoTa/crd0d3UZdBdryKksEbkCzOTfahtXQKE
uXzVO1D9Z9vaabmtYui2BhO252bYpcmHFiH1gDgEnE7JKM3nZb3DcnubWwvu9BlYchNfcoO77Psm
LQdzqR0f3ctrNnUqzqHgTRJQNhhgFTq/Z9Z5FiKzsnz9KibMl5FICH8uSrSxbIJFrJU/bgZxl6TT
8h05DFtu39/LhiGVbuhB1uecaAbddsAbgXJvVZd1DqziHs6fdD5pyxsOgf++U2ePvPQ3fjUoySTc
cT6Yg8gjdOezLiMSHyAijZCQ5mKcEFI7t8VgAMyAlNblHtW066uR9XQ2m9w+lg2uuWyI5VFkR/Vt
grBi0Wgm8Qt+khgsXHLlwDBVS2nhIbXUGOTlxVtwH81GJWJwxLGjbDr4fPH4VOp7fPeGQqVOTjZp
344LGNGCY0X8gIQZzRWwUhRiNW68UAYqhlGM3/I1toKT82oOTLe7Q/sO5zKVk1k9Fej+kzllfo8m
5G2LY2sGXNL0/h90f/WrjqU674ZCQdEdheuYftPMfnMAsIcjt93/YLZbBsYvs3HDBjg/rYGZ+kvj
DV2PAk/OkYAYmp6f0OuilQ7MvoP38zUilXW/8M9m0wbN68qwpSgPGYjVe7o6Gft5IeprL/27VlKH
zVUEy24VACeJMgocrA49wU2YhwnSkw3Ch5atH1DeP4M1QD6dltewJSz0+px3L5nrzjs9XJ/cbwes
gj+bFftnmyKm6OrAbxx8D5tkEg9VxnOeVDiZ4bxIde/zbG7A+xMT5w7ThdQDU7Unya0DMHdLiHH8
ps0rZLF+1gBiLd6EfJDeSl23BLwgRJ/JC954Ov+jgkDLTiYYvMreaMNhkwpudclYzpT1ZUc4BD7J
RCFvtL/QhoYwxe1WOVTOSiPkq3bvQsNxuHDHRcSqbU2GCZbZ8DM+m1GauTUOm1/oT84VmxCOJfd7
N1L7LYa3IZ7ePiF+Bi0J4dHdOh0lfxLfqC85+XfKNErvxsj4e00F+fNUkDUQ3st8pwobRMD7M+Ba
aGDtvjlmCNMycxMbKF+I2c06tg0OAF9M+nnmHR5SwxkYj5+GOcA+GOptW9EQn6Iz7C7ZmJ/BdQvj
sg8gh9nisKvU2XGI9jc05WaTDiEkVtt2HFfQhXGPU1Q/LPQNA0q0p8j9+dfym0eUcrSwZdqVNuLm
u08JN+jGqLpkvZm8TZ+wJQJydGZuGUkObxc6wIKl3o1cl75Iq2GPwTYpfo+xXDlRyyStuY2IG7EF
fBkYV0Pfu6VF4s+hsq5PnA0LeCpWNEBjDljZGPftjeVFRnYrBW+ljp1WpkEDLOm+lBZpRwVUwTFm
gOnCbszSzc0gmM9a5bEMvJzXhjpPyxp/OUQZaPXKKgf7pFVeXDhIpMdzQth61VwJADI9NJPzyJaF
uV78RMyr2aP9i0KS/rbigW49wTGe1evDJNz8u8dEyL8BX0i5r11zSnRuUJ3r5kSObT45+tlrakOt
JJUYyVqg9GC0IkunmbTDjv4gi/HAi8EzjRJoNYE055b6KezpHrdAyT1atVO29kV57jilO2cpzBij
rQnYBl4nx8eCxxvWtDEjm21gA8DaIMQ3l0wPtByqTFA1R7fb3XHmX+a4EMXeWu3CeHkoGJpMsP/B
kmOUvo0207c3FaojQM0UWy+9JmVseRCrM3JwNwoaZ2UgXNFvSvnR2Uc2W/kT6uha6vhUtvoANxO/
iGqdeMqh2trXvyWbOq+vsOQ26ivtCiaGfS/FSs573jOoj/a/0hCwXqcOqWK2XJHKmKDrLdjIPWAh
nZlL/isGaqUJlzcTAifFnmtvo8KjeWx9Zxl5lkQ4itrOzQtFFv6OypNvRyiJEnDAvW8hUHUuNKmL
PH3VSfhJkPcPWaJFB/ql/zo09qr7w0N0YMqToivFZz/lsGyYomeiShSLlN9dT3OR+p2FI7WqoG43
ByZXzRTwNWf0k/V32T+rOEt67Pnz21gOR41D0Iwv7qW47GKQ1MOf4MoqxbjKGfBirWNQwgL9lsns
m4DO8y3bJWXWadRfViN5myo4MDBz4uwURaUWQAe4sQIKeJZZeqOoSnPSKg9PULgASpilRFJpThiP
ZGAtjPHs3f6ZRBVJ22xrqUUVF9JO+Opiw75qYixvH8ZFQL6Dvqq3eIh+YNzQR1FoHm1UFXPFGWGJ
e7ZspQhV8f2NY3LjAoO0nO9HsnQOFlDJXSpnUmrxa4yMHkSz9AmATFQyYAWLwUnrKsNUT0lCCLPu
m9h1Ku8YeT38xNyBGEYA0f2h+EozU8QVCvU1v2O4nXzDngwvDbUgKKK/emCz/cYWFTIBc/PD2OyZ
e6SEejB9p80vPYBCeeszBbRWnUm9FEHc0d+xS8RmlBIzbg630UWWkHwDVB/h48KWhjm5dTREtIih
gnYPyI0xu145attDP5/sUrQiSGfU/NBGNQuotlJ98VID8LE0rnPxYNCPKQLJCVHJyBm5cURKGZ4T
Y9aNLy64Aw6si3Gs66H5NaX8TGr3WbRkfY/RVz1UOtjfuHle3sT4ebnUrGERG6TOllVDhTfUWx9A
GHOhod2Bz0BICEvrDAs5A119XZ+jV43ymx2N6E3h3iOX6Kzx+3KBSVPXWxLUpLdvEVhUcukkxfbK
KkVv3vUcykTZ97SV4A/MIHbhovYC1XvLZfz5nQzeH7crb5mfyaytrolbSKXJrFBcMLZ7+mMmTnid
+N9Z/czwHPSoDXZDmCOmd6YKlyuiXgeFpweNgg8DC3kMqOIKF1DFmJUlGnuPsUxsuWFTWCUAmC0S
WZawkloU5Zz/pAyzP0yJPNpd580wEDl/95nbUgTGdMLaGUyIH57g9g3N19oaIgVRYUG1HR0kdz0l
0+PL3c3sGV8J2zrHUAsgdntxLDPCOglXDXDQE3O12gfisftdRUyQEVhAA/QDLX68CpreU+vtoral
I/bDAGU8ufyOOLc8Evitu7RUE1g8nmOVfK3541bsMtzTIGGqQGR3GVnPdw5m++PoruWkqz5k9b10
ZJY4YGw5NtGb2eFCm52U/VGVvRJLC5WJ478a6bbH5lstVQbCwFcMNetZanWZH/tibViX36fLFnRt
d6MiVD+GnVuX5T6wo2zMoQEGYTSE6RRd0IgS+AFWk9fy4BvKhW00O8kgOO//OmqD150SUiGMU5dr
aOj3/LAXFJLA24cfWnC2c9dOANQM6JfxXzFpeZXDR19MPjYlyi3jLx0CCI3aiAGjthRkqMJ90W9n
/2PPwXwTt0tgaESK7h77L/GjQX3QMSmUFD0QpBmT/sXKc6T2RzlTpfCaGilc1vY3ZPnyQSxChNYy
NxFvbZdmWdbs5FKUgrDRkkGEGRB0OPkg4nUzUMZ7cK8dFM81TfoY0GtGwXIreOaik3LvqFaZ9jn6
aJUJ+Z1+3V8vqW2ZFuFk9QNJp6RecUxqHpxTQKPn8CyUytiwNs+0AwLACIKRjlpgHsD5TOsKJhLm
m30yqhBlTz+go4z6v57PgrRlRE6tm/64cKlWaZP/pSa4Z98qf+kOZQGgOkgsOTMrkuquDMYYtb7I
M/F9Gvy8gd2XHf+oit4GfKr98PJj2iUv9uP9JmSb3BsZnVsPHKyhqSV8Qyl9Dc/KtBjSp32O5D8m
L0qiOdlZuD9S7e0cMLBRXqwgQm48GM8+gVwao0E9JA43LVp8OHThG1t2ozZa8RD/mdDlVv4YbiqE
WBpNPYyAiOa6ABzEo/kiKaciY7LJ5izLy29pBW5SdSXkBLckHkLZDUS4pHh6B/iYLZeVqbF0Llo2
yfiMwBRMq9VwfgdKk88QcwsEFIKHNSTDoEOyQjrWQIsgk7h7wfJ78l8sRgmh1t2ELxHCYqcajWDJ
ge9yj9s+RMXEQdDiE8WzzSMnlywW2YG6MQfwjMnHuS09MnTUUqZPTmIFMq2ElfKmSClQfyE1z2dx
ptRMfxMIzQC4nH8YgQT0VOD8Vtd3fHfeBy2AGn6p6v+URsD1xSWFj7ITsMIWnWVJy+VXsY96Bfy9
hnWYsPHc+/vcs0ytM9sJ915oNBywAndQLpOX/yMu89FCDElNe9dC2KPvJYabXTNE9U4Xj3sTf3kr
+vYoDymkRx6tP9uLYzP7NfwSiHIiYEgclmUQMlwE3mPbsSah2vvDMhY2tPpvLKi/XoC4qsjXUl4n
2vSNjBrJ2fUrwGCQo0a6jPDGUXom5DnqPaH6IK/6N7X5Wnalw53pJjsyeSjWPHkJze+zMvJ6YbW3
7bIiM6hKe78xWqehu/vpMUJjC1tepa3K2FjSpwz3y5X3pzVu+I1nIBI/e9dJuqO6F2t9csnSJQmJ
9zbA8knUEcjzuRPO0hDxbFx8r+0OgoKTewR25KWPYW1qgEabH8PQFJTC0Vm9RsxKEvjRZ0T5TWnm
+Cs+H2FycqWBmCAED119KGfCtL2u8VV4Y2Qnbmmm30oAbKcvmbk0dMR3+5gthhqhKi9jpxC82pOx
USR4Vx7ThN7U3KVc5i68BR/wicQ0ZKWAPTIjtddC5ltggn/AR7tzyeuVukDIOraLE2322pc22PdU
CZknwLq3Tjc9aL/MnvncBfyDPNuPrkfgvyfjFu96sfih0cf7S5mY856h9X0YlkI/ATtp2pFrSwxn
XlCVb/VxCt9UKTbVZ7CyuCLtEi7+F9oasErN06HMvRFDdw2AptcPgkls2mJXb4aIfNwDkPP6YxBY
uDIOiOVQzZT13cUhWkJIvS2ypZ+NEl1t97vrJEmMu7cIVfuKASyccHXwHpXsFN2KpOU0ZdQbUSQE
Lp2G5K3rCk9tY6vvH7RAZPCHwJdJp/IcZyYAJT/edDLUTTkWkNgeemxVOD0KnKyAoaiIB2IeL8Jt
ztixRNnecpM1CN/HZeQAtaYJchKFuxVwWLN+CkpuJRDGgLaHyuVxaQIYLkTp+vFU48sjLtS4pL6N
MqjDOEHJcNez7+pJZsVOOrNvH3qOr06WMsMOH82Q8AnFXf0XFCRC1NLPq38RcPqsoN6j7bHu6+Hx
8UvoRP0Xw0AOD9WtkQoPjB7Ij81JkPJVNlodpG0kmmwx1gx575C+XdVToBHGkOGCPuh2A0FleaNj
9vzpfK0zuwfpZlSpUrUPzSQg9E9Lxx1d6IEARSDEa5oI5j+scjaLH7hpz4SQww+Z7ygr3Wp1/bjT
QwSvV008rPX3IVcP9odyAIhz0SXXN55Dpg7kaZh1PT+r129zZtUI+P+V7QoKl0haFj40JlStS5zM
52Oj5iriX5c1anM3+9h1mtecF3yanQXWGhi9GnnaQszqc1viJFPwpFvgTA/8pSAC9t6BulJTnrqq
vd/b/A9Isqkz1VApTYoxrIBMqTOd8ND1VO4PWiZG70GiuSpVJv033b9ryCav0X3cT5Hua4AVoP7m
RJAnIe5wf48OsIA/3Hjtljn2FZkJEG4F83EegIw5D7euMkHeVOgUkcWXyXWxSPb8xWo6823HtZGo
yKjuGE3az0ixaCVKR/aGzip1fdoh2WfqvsgmFK/P/wrJrF45LDMITYSGWSumi0wUWg5u0OYhIJQ+
uYafCQmvW0mNQA4oNuw8EdnQQK2Gv0Ut6o5SrNsnPtMI+bHrEx948oEBxgt5BgRXKJOQoCzAKZya
RhevUwK17ESRk/c22+ybxp95LgPcgSyaT88SXk7908MJm6EmquvmxWUIyerTfaP9c2OxacugP8n6
d7bP4KmfYoScmbkotsvm+MfTceu/65Jx8TLgHPP/RR+BbSDHsBuwo8O+gxZhM+SAssjmQ5QcLwvx
28bi/alk+guO7LpL2Vkj/le5tvE1bwtcCK5TmDL9ONGVxL8QJjhYJUsE7waioYrirMSbClARVfx1
NKvbII67mgaOiza1KJ14z7GM4FaGQJl41nRO/sFj5SLubgOlC/9g+H4qZvlwc8rxgqPjmDLtzGfP
pFUtRPIbubwlx/9rh9PvKfTU55WnwlxOfVJ9rTh3c4qBegXw7Kcvy5E303YDKXYv04LC9+WRnXF2
0+E6u4WCawW4RMnz8PwDpHh3uwE3c3wTaCSFGW0kzZdGWfu8bPktJyhjNgHu/cD7GVINvXy6iDUr
anR7MRMFUcJqoAbGLnl37n2LD6DtEc1FBx/vrWQmguH/kixkNRXKQ8nysnL8ONq59BA7K0QcS0VY
BM4MKBV4OZGn6sxz9VSAUGH/J3l+7sF7zGK+XAo/cc/0U59B/pfxV7N1hKXAlIhBAgJWH08COLsr
xmpYSn5iflC6g/rzpP57sRXiV6hW7PeCMG+ofBWkEmxEgzYdbYyzJSj43E7UJiTp+jWUy7IROYSg
aKt+VQKU/V8RpCxqcfXT97cdNHr5gf5BArlhGKxfkF+PBk0EE352BtK/SD7huvxK9NLiYi5yR30P
hPOHc3kUBqRWrBkt2lKtMNYmhKOm1MuS8qUG9ohWVmB33tWr43CKIgJXeCfYAmtYnRppD+53eC6i
DMvM+bUep8OgRmdZ9GNIV/n4gLwgLVA2DMGp2Oo/zvr2sJuPpR5iNhd56cZDR2kDfA+e+XUuajKT
iBBpHy3TX7Zzr+kZ1+je/Rp2zxDAy2dEVNl3+S3nVwidUJRfdM9zrQWvi++KWQpSVE0D0dO5a9/A
8qrAEsxMFeSLEL2R/QzUWZFlDfuVqyDqVgFS9ZwI3SjCfQBUHwVbpJnEcejctoE1jKZ+x5bKxEjJ
SGHya2L06MUrBebofFwB8fgRhP1aEAoIDZOIxTXzNMi+bUE0BlxQvg0VnI9BJ6OixhGxxBRsJDUQ
1ly00d4e3R1EiB2urHx+1B6b6uPuRL+aOQiJjGGHBni6rMOroK5W5EyElqA4C69kTMN4iwySoIW0
qNuLY+rQZFdeEq0mFijMY0d8gJawoK7/Ert/XrR1TduoGi6la8DJMVmh/f6BU8Crkrmt0Y0/ksBC
8Y7i6CsQdJDn1B1sycUqnyqJoQl0gzYqWdCwhPXwsdaX1KFXd40aczhBe1XC4YtIEIfNUHzCNxbT
+00HeUpvyWSTWvXpqtbxa0P7BetBOsgQ/yqFBm4jGGjes0l+WAgCu8gwjoZo3M/NCAbX9uPqFkeC
Teobl2tTf+WHGHKS9bCf62iGoxH3TtZix72z0XfPTD895TaWnSpUBDLgl4dnuhZ/Df73nGi2jvFB
tVl4TRIbEOFZ7A7xWWlh2LcRJoXPE6FYgjcnaHGG5Hk8p2U6x5ujcQACktnJpznm5fWCsBs2Egab
1oR3HGdvbFn3ijg9TnqcrfqKT8lMFf8Z1sbW1FWcqC8zWA8VQbzypLctvuScXl1MAQdLufvkjabv
YHfi+bCAo01+SG7BmVE5V2f49gUod38Ll1NGP+g/SbDloadDY0KtxGpfMrAnpq+Lq01DyXbWtQE8
H2aas0jmSDZKoIDtY0b1V5zIY3j9cwI9rpT6AG4W2jyx/odq8ZB/npthPMlqS64vkiIffQF+DCCl
Jyeo/ot9LhtrkBqKJCouK3AyURYkkzmITuRBZ5mG5wpu1uAouK32a13w8wF+2VhyEDoKZ29T4OB+
/81i2w3Ajju6PUKiVjiuzEoDBRNdRaBXJKrpZXB3/HEGnSdb3GRrONJFWISFo/2C3chDyAp1QxV2
qPVPAl0dXwL049n98o+RxdKT0mwFglBJtF3Io3EjbqLAqfxwgiy0mxRYEkbLlAHSzIW0mW6YpIbZ
XSa63s2KBYTLNoiYWKKRNGs1d2zvevfeO6o1/2/p3FfYV8SN94l/zFdHifBbXOD0iYhpBisu2t39
QrKta3W1rNjootYN7IgalHcP2OrVanGJFUVUNGNUSi1fI3NGdYzstZLsrKUayv+MAQTnjuHIY1kh
m5IP4CXSjSYGlgRnyWSW2oCUXZG7y8qOsLt8SjK4LU3hrpoPsmM43dHHY2j4egDjMUXJ5klqf1dS
elqlJ4ldMY0nCmqWif7QXFd13Miwh7FvLTW1JM6L1pBQ+7wpBgCL5JWgdkPidTe7yB2Px3RraOSL
+sOmfdK60MJMCtyw/FUpi9pfu8kDUnVChh/81fRv7E5FGo20bVm9OqLOl0qJO6+J6UBwcIUJs0dU
3sFQNJ7dg4xFnWQdPVKIcd/XEystnDrpEbQz0BU3pzL4xy0/BHnULyMZrXRMfoIxJdiYD7QXkBEN
Zj3LRPjBvBTeBSYOTs0IlMpfpHdoY/DRtgBV+QUKsoILvujUEZicgn1xURy/sLZX7ajCdM+M2ykt
+rvlFJEq3BMWX19/4yFeQejSVXzBi1Q0Ah65phCFWQEJ3i3HQfi3iv/xQSHhK1rBDUvYof9tBJYT
sSLoWR/I7PWhMDJeiCMe5EeKzZvD+owO6avGT+wP78LKlxyrpmrPx3G1Nd5RxYw69FdXnDcw3TFd
cOyMZrfHX7Tugd3t2bWYer7UfFP4IKWDLFgfHjhg8qrzwRa05gPL/kVr9Hee/MkQkGq4U8p+0c9n
GXziP+pmHzZWGCWHJHaoylK6vIFRejcv1t88IhcEe5N/P7U9GrSMKOkK+mxnqMA5FECnJUMCHR/M
MozJ81OJraCJnmbphdi6kUEvLdASk1iGbkpNsv0XmduZdsgVXoNG5O2qHSlH6z5BPIi9/PcApyLu
HAkQY8FuD/WdOy+z43rUveVbM8WMf4MbxDo3rshw8//Je2jFqfbmb8FbfejxkPBSIvI3aiLxPn/6
Z75rkoTv9AgK/bY5xlSS/phBoBaJQyIb7Re95ouWu1gYqkO+Wsn5qq+GICtS1YF9brKvWY9hg7+V
zOnLern/ueAkPLFSWXPYUc0nSqzIQB8XxnImVUqQts9Jd+9wZnLWpVab1rM2rqiSSubfGsqsxz+h
A4bTZSmdeTJ4IE9jinpbBSkzRpF/gZml38YCZA+LKL3GwqidLAGyZ+ijVcUceOxc7Ocmsu88CpRw
hv9cwddpwZLuod1hQhgExpypC73btItMpNOcwoP8LBfo7yXSmLw6B5rD999ZrRy+0dy13BKJ82Y/
Kh2vKV9K+VuIgP7IoRBu7a9czKO9R+0qbGFmPsyOFIcEuK57r5/X8JHqnDNREWDcZ2DFdWa6QyiS
MUa7JcBlSGLSvVor8oOjvzZq9G0Lqt6HwxrOCdibYPmksIuwK6GI3RZo9Yrwdn+GW+MPqke6n4xN
uxNxseojlShdAbXu63gbDZdkoRAHoaWm9M521iTk2B7IU3+Yxo4/TguP9EbhvQtGdC3naUYlkIHC
FsCrZw27ykC5VTLiYBkJefZy24KAkVAcvuZbxgBqojekOiVMywK0k2eqXjfoN6AEju1AOPLTqF5b
wzz90/4V9mKtFBeWLn2b+Y46FkyoZzHHgHCfaY1sTMGvJD7EAK/S/+iwpv9yoEJ45DecVrKu2PCn
8LVmOvWGsIosttDOjODHhxKWxWBYiPjhvbYNWFQa23VHCRGHcJYrfQxJ+I8r0lw3r3yMAvwOREXt
jtWPSFO4i22glXK+3FEciDh/lnN12GTBIWSR8c6e0tJOuBnlSRSsNm0stwfCuYdbS64SSUMjW8T6
QBQAd7JINzQIHWmDfFMaDytqIooWO58OvquxwpC5j6b4f6g/0uJZ5ps5QbqNnGE5fB06d+aaspbR
TCvqaKMVvJ4sEiDQ0tf8BZsfnCvHvAMmhbfW6sDhM6bKosPEcQHMMxyTULvcTxEdMt+tCsCnDMH4
KXvx9gGZeATLjW6faq8625yZd/XyO37BIQnh9ejVrEUNXgwnxe1yR+NxA2laAeZH1elY9s0FMGui
FdO9Bz4bBr0O2DiGRqKaCnOmD2ytL/AHLuHaaptwBfCOr65rTwaynRszvkdIw4REt/Ehr0m/5r0X
uMdeeNO1qNNswq2Hg0MIUNeCmYlq2duTcLwk7c0B7jsMeLvnsgAu+Xcbb3EnVgscpg+KiDULF2nJ
8DvJyQXRApiOxXVAWe3umebodtbI45gpUKzm6gcXzY4GpNTEs+xJAzCfH8a9FOXU8OEwUxaiNBy4
E/upmQNrJ09CL0NbQPMkI5KMkQc6S4PTPUIoJRTxJU99NhZBiZNSvqFviclMG4MP4d28+6Rqer/c
TauRt8xJ4K7JhQ1e37OUU2ktmJbYNP3P6/RCy6JDbNmg34YMMUfFOLhg1A66MJeJzJ7iBaoqlI8p
Y0uVHskCvpQM83z0qWQgr2Siy+ZPgwwyOvLOOKEKFwuXpOFnr6deEINjPUnvghJ0xB4OLpquiIN3
39g0DMoB+DMV+8+Y35zyz7wRO3sIlve+s8U6DcrtdSKsSIOYdcBRMg445+3IJ2BwoMpdBCtDpt31
PDxSCpKB9yBChPob/E/EiD28vvvpp3MGz9YcQvu+aIQQOg63AHp4IN2ORVSkgDoQcpdI1J7LnDC5
0pRolwoqWfvRhaQehZuLnvl5fBfhoeImEVe6wu6TNGKdoN5KpinpAgiIrj2ESa7jdG2/CjkYGRzi
LT1+1k5j6yyLCMDo0YGkRoJ83UkjA1EkufQASlp9QeIX6PNAZoWxy2mVDVvACzfvLFHjO6KIPbY6
y7iug1pbQpopb+R9KZWf6ZnCT0YeTEEztqt1WLDtqyiDiDA0po++GEDGcobVaWekmbAvYCzheng3
QYPU+/7VESQEGgaA9WSIUxBvGdSWAkId4haFy9/USkEXUbS5LzzwCkC2jFC3P42YU+hZVpmZ2dey
ZUHUyPhwQuSlbIxAXNrrkRGcqM0hbJyRu5ASWX5OPGB2huXMaz7HM/a0ey5VHDieMMS6v2WM8Fgc
SxUSPgA8v7CawmfQURJlPtU/LZRoyRsAXdBiXM62PvPKI4rYMpxot2iWmfyqlYi7rIuZzqrz02mI
ChqoHg8TLzgmfsNht7HuDv+zgmHoi6awS/oHWDTlXTeAGlpw2+JbIK9j8ZsxQR8inAYOze2qQl8F
P44Gfk/uA7wVFU53oi/hPKEGKp/xuQ/j0WmA2PZmdV2t0YdIyz9qzf2bVeKJhjlhKyi1+0JMUOpp
P7cpbroum4dvIqmmG3dB50jon7ywN2eGN44aayORTiieQTdJ+u/DF76irig82wgMuV5/I5Xrht+2
8p/FwSgL2m3znb7qNZoJ5CqL7GAZ5EFjjso4MkOKL5Sz5yAeXzU61RpcrsgguWMS0JvsCkZyPa/O
R8y+4NOEayoTFcEX2dG3k7xAgWZmfZUxR+5pQVRd6mqZO7tSVR8botT6n1DBqM8IVRUNSvcggr/1
kMmzICTewfmV8uOlty0pAvtvY/mmHfIAQmPqZ6kMqLmmHqcseeCg7hcBwx9L+Nr9bIb67jSXFosw
0P7EsOZQuSgI9a+QxxJv392UHktBeTXsgBD4eVVz2tH0gui3bOxi/+Kv/+p262GuaFR0X8g6SBHX
vR+XxFPr9JSMgvJ+VVO9gmrmvgtKT+agXth3EnHTWxeuvU2dGorjTrQ6Me9qjazqDlhcYZiK+2ms
gGwEV78A9WO6tfulhs5V43MGyAuZ7uHznMxchQ8ykHdkP9DTzIiCII1NbqbpGC5MySdDvlzxOy5+
Q4CDBaAq1EnpHdQWUcAqVBffk4g1VD5KB2IR1kRBG3q5BipEVAr4M6jjtPL9ZtSPp12utRiTL11u
1ZxHMmnVW7L9AR3o59uSewXxnTN6hrsxKE1PImcnCgAu5RwZYxnr7NqWjx5NEoWE69lZXxafF+bd
/xMtGLDOcUPQHkDx+FhH1C+m3sYKmjKE0ArdS9DRGxdBmDgg3qUHN+LbC14aEvFLr1YIA+b8GJtk
2ppbmlyYHBDd7xauY4FsCs/0Rgyl1090TDtibP2nVH19nCX2d17qz3UAlBUpt+DiGAm3/3WIwD5r
mBYc4UkHjNPk79GwIkKygIme54DqTo3hlxL/iPnGF+91N1ogLNZ+5ARTt6xiIil9l4TwLDPyPdgG
eQ1xofBNNSEeYuVXCDLaTonXXMAVdZ3FN1SEoDgtF2imFN+ZzpmwYsuVWWd9Elx0kdFWyQXk0/Q+
E+6Mn4eZogPM0l4YXTSeEg9r4e/n9hE693yciWVHHME0HUp5ZzXmMikTtldXLjfkcCgnIf+NGTLW
xV3Ip7/DdzE/juAxIzdGVUF52RUH4DBY8bHBbpymokcf6inY5Yog9OadkJ5EZzysqDx4YYnR09lX
b6+LEWNbWr5qx7y4xiJIdULPv3q+lTt6+jXvoV28yIW9L6W035ons1OYOyR3BlQBbiH538zAhA/X
bE+q4fjZq5lGJ/5SHLsC5/a+RQNRIBmZRf9IJ7FQWTK8VBa9hxiMC72zP3/HOM9bMPf7665aUqA7
QGfpGYT3wpNOgrjl9PQXW7jz3P20zZffPZRg7qpAZivSrg90z+SwCLZkmS+eOiRelIHdVu1bv1ev
o9uO8rbJHypT8pXogLFW8YZrqvkH6ke8+fMEfaMaJztRR7Y9JViRWuNlPRpkzBpVyPc80cNz4+8U
0aa94tjWm82xDnXt18hZ6IEe6cgNIi6ys8PpNa/lvb2+Do5YsY+2b9VRopVJuq6MQNCWgqJdU8F/
FGueca1rsxstbD6PahEHNDY66kTcu6+8uAe4s6bO3Uo6uWx5NOw98NcC0Q046K4bJUFMakLZYuy8
lryFZYbAz60glv2uxy9tcrwbTLgpptQF6ExEOPsNhK2AL/5PceJgkMHOpC+11+WBEHEq0AOAIC8T
Wo7OWGopTzj/A8PlYljg1nXKzdL3/CWfpfBnP8xz3hexpoQTd+DXfWB+QZ0JflWkCyhHDWsJ3o9y
cd5Gwrm7tVTTxgD5NMU5ww4peLtjzPDXJ3vigSmvbxwHqjOaM2xEAVAukduBu8uYS2Eyidird8w7
c+lUM7I3j8d2DswYbY94yf2krIyEw5X/zFBwrsDbRp7BansaJLeZanKfS8lUZaEaPMmQKN3JrJS2
w21SFvEok9A+TCwpUP4zVO8dI71RoLXejo5pJ8gPg7sNTt63Mjlg/jA9zVUITv8C4i5ssbQ3ufdY
0hWmRw423JbmS158k+HhqmY4zngNDGme11PSAcPDmXPkksiULgOYTNSnINF1G3lPzR+kWzRTlL5Q
5g+WkhR9GbgsZXLzYPVMx9rLzfASgJpBliRvcMxkma6ET+LazGUDheFholYLkwyVtUeBgXAV3xYs
xB3htYCU2deilBFzkyS1sdGEc5ciCdhcHa+j2WkOAc+PfN6Xd0z3lvTy+Fnjpeq/eibIBBADnHpX
0Bo3ADzvJC7nYgWvXBcvZdYaLzIuQeMmWg4fSEmsvCLtJFXaUe5Ha4KJfVhn1RWJIBxnvMmytSdr
/ZWjoEtjRwC+Li3kHuMrjIdjHCi9xx+S7syHk/0z0ZK+TIEMDSJyN7Xmza+wMQaYOwGjp0LS6DtN
Jf7W2DIklNA9Xv3zC5ATQ2CMroD/dOlz0K3RJaIRL5FcXEStcuHu41s0WvgQ02b8xYaUU/JAVKNA
IRMF3ZreRLyrrTx4NmEp6VS1XPklJi8//GUaBX8WymgdtX6j3Pp/V0szBUiti2stsAJQY1KESmcQ
/zx+H5rsRMUfJrIScmy6l+r5qmfZ/UykG5h5EiSIe0H5JDGQMpz26bykKrmhWBfhs9ZpW2YMcDQN
U9K0oZlDSusOyUbBrPoqAnJvcifKRQr6vKz/9GTXudWSMkirGJl3XwkvEnM6mghMWv6Tf3WtzkS2
GQk9QDi+Lm+FcYn5ttO1n1g9pXqnZGrHlhOso7iZPzPQ/VbDfTBSfkEY4BtNWBCdRVTkzgbkkjHV
r5rza+XqENSwawT/6s/w66+rDvevTIsyfd6POMHYxS7UBcwoplkoLUxJxHjJM4gnOgPUczzxX2Ie
ELPwNNy8QcOMjFsRkeuQQVeUsU1+YM1ZZqd94hqMyIcH5NqvMTTumCnCDTrRHNISPsk5cXegJL5k
6LWyZ5r3sk7z9tAUvfG/FHicpC4zpWJ2I2KblCQ2uQVVx1bVNkhFUkEggmypBrrXBcOskhyIpliF
wgzM2GpTbQ/yVEPN6BxosabTCuYLiYE5hrimExMa2GCSTSqknxti49pFqJllqHBm0AHqrtMn0vr7
YCeHlDTVgnBuUVl8+vMXU+cjA+zVc3sBHU/HX8amYuV6Dz34quHFIOnyPzvUZqqoweAufyH4zZNP
aKlSa/3A6PJt+NKvrbhp+lmYCLhg+Vr4LhjS56wQhaxWEZrtr9Yg0b8a1kZQPeXnptkccq0QwAj8
KZRJcvfIPnAa8z9my7sxnDXJQwQyvEeblNUj8gmVfJiZtG0MCrLcDvZqgejcAFD78pQ8JjTk3WF6
3aroamgQrINgg4JJmeHQBN9zmPgtKeYj5N9fxaP/IA2hpPr7eSyQ04Gsck37YJZn553P9JP55XuN
RMVxSgcyhbflFD04ttHziLdkG5v7zqrlz6iW3Fq3SI5p/J8yOGkUdQU0VKekk0Xxqcp72wLw5n1l
Mb34k6u9Ff6v0Lg+iBMGIuTy2JmMCmughpyIy3Fx1frMbwcEQksxU3scSfPcT65dLZpajBwSPIRu
5L2Sn69Gs4ANjNTFSfHFmiVPQF6mNRXSjSGtgisIiSv1cyn0iyrQWJADp49vUC2I4OqkcdVb/uJx
Qz/C5TDxm1jfMmOu3zRD5PCdCku9clladLVxtqsRMeP96IeKwfvqDzPOix3iHONyPtZWGdTRNDGq
Qb2WF2nzew0nFryGiwMzgUVIGrS3D3Uv01OecGfRq+KhRBub2VKFEiA1Wqds6puNFZjue5JwyUci
HOf+Z8SFKG+/8/pRdYaV+895s498Nr3hH+DWUAyCfGaF73gLnQyWI6ES+mD8EkV9g+U224S3eNsj
ObNb/49emU4Tcu1xUjzKnpxxIvarHtMkX0mJ0UBoD7aEDg8hJ9J7INGv+DoKYNwMmQvYhnVQCIRA
K5dVOYX884YkdvkIAe5c/jvlkbbsLc3sqoppZJKQkC1Bx09FlgHs6mZM2u8B4ARRAnBTGvDR6eEq
oiyfdYqS6nipdX/1kAAXz64/EZ8mmiUxY8DrLZc1KHQIFtdQL3z/BV6PVUVxHjZ6JBbFAoCYlFAJ
eQfqT2gND2HTxD2C1hzA+roTlF5Ys9+E83J45V1gOsdMS62TZhWKuTuBQP8ajhgVh5ArpDrDkL/9
ca/Ef+TtdK5Tg6OTetms0EnEy1UqqpDUfC5lIA9uNGGbcshxLfMfC/UcTIc5uPwWpJmBjTk9F+1B
V7DfYrKxlTyuSWMvU2hGXySm6xHAKN2ZLZClKkuZfHkFqxRxnQX347t5gKAOJNzKmBxpcyzxZX5r
xqzfyxpkmGwoEb6vZTap//0X2hecRLqvjmWjKqnD2AcZxGdynjG87WIzmME5Z1Fz7t6UNbXmg6Xj
j5r8HlSvObKOO+camUVdjZRt/EeEQqG7JEMtHxPG9iBjdcj93uLBLEulZzdFel02tH7doTMACbSZ
30cqMHbZeuNDMZjwFkEyAhDqyhMeJn//FJRWnplieMx0QEvSgIXV3USKFWqQj+xeCmX5gGL4eltZ
yByQuFfR020gXdOQTDRvcvFK7rC9goay7VU0UaqnMMVodambKzIlSDPRz/XsYpssA0Dai++lt9/R
BIgEwWbpwujqKEebWcNEnDvrYl8LJ4gR7EboJCYqRMI+gxSh0wPYOo7C/WNsm4kbyp7T3Ck9OlxB
JIgvcRfQn3DWtGRoBVRL3T2zwg9N5UnjAdP3AXCj9KzbsbIidjwovez7xS4iCW4BtxaH+/oYA+fr
hRs+PUTqEV0ecSGv48afJOFQKfOZ9rpgeY08lKBHK7lEO+e7gqdD0NaZyJ/4tMhAFf89My83zFNx
+8IT6z/wmKBtPCtwORFCaKm7KgO3Oc9RxWnuFVS5BylvpUUh4pE3Nf3yz1ehxqKJ682LY+wVFKjm
7iFxNgw4CI5gwtu1mJx1OxvX+1ubfMlE+Zg1qnFy900lCrl2NolMz6btZQ4rITKy3vKKU4HmiJGi
dtIPKWF7/D5ARGijHmr8W+xvKxH8d/CC1RlTVpdXofm44RKiYs6qV72lSzQhrBa0rD/QUddkNhCq
RCrdR9gugIHSZLgfFHTrn8v5Z5dDNnvYsCBe9+9jl1L2p5FRY8zOArTNsqNOFpQcphnraJ4rvPo5
OKirLl777TbHASHrD+dnSswILlUHb45+hjfdPSR9ymdsrlUhKMvrbmC2wJ4CjXjTNivJDUAyubm9
YxTe9kQbWXLRYG909LuVvvX7LyLmkC58KIfSEWuBcKVbiJKRH4Mp8FdnB4UzBL5Sq0IOUsSuuYxS
XMR3sz//hd/Rj7UiotfugNxJfx0K/aHUv7u2hckEiRG4j6W93Ks0Do4Px5pBsE5RwlEyDJcDd/IZ
7QlCKckifVRR+oeRl1ReRPp3dfXz9TwrDMDVLd4QQSksdqmLgXm5dfJHVLP/OmAZae2ceMuvVEOS
kYRHOz6U0o+jLrK6aQV+fYCtypJEJYH9ZYLoo3ylJWmggz4IjfG9xVGM+gOJ0SfXpBcWzsj1+qXM
DQL7xswnmFOWfPkX5llBWWU922AoStcIs7UmbXkHhyQrYZ6KW5LFZQop+PgChP3PIF+oFZmjYYLp
8JFnQekFRjT9ikaCXxmr30svrNA4+ErzmYtBncVkNXTqoTD8fhAJqaGk+j0Xqgyg4lYQQJ+6XidO
/frCgRRjbr7JT8tKRiiI3UNwh3mWG5sydJ18j4MdhNsKKqsCoWu6ElCqAXHJSdgn2eLuQy08oXgq
hszexZ3tHd3rk/loWZ0+DYRqxsVbN7Ws89cJBadbVxmn84J+gnqbxy3wbCUV4rqQyFHPbz6nOcF+
QsjDXqPD7Pl4/HAn4Mbm6QzVRXOxjKGC5USHvxKwzRQDUOSRVw6qK5pb906biYwnb0JCV2xpFHos
XpcEnrCUMyzXnT9/dqiKRaMd/gaE8ZIgBeSPcuqcOPhE63vKS0DVqPVjjD9ShInfl0KyatUw0K5v
sRdscu3z0OThuWnK522y/Mm+/C89SN1P1EnDGq8dVK7eUciOfO88LjmXg+knBYDDomh9tTKpLxBX
P3l1Mr89P1vfz6dB220mHr5OgRzur/4z39oMTWgx+JO9Nsk9mL0TEWy/550YvIX8XhB5+9r1w5Ld
Z6eDIP3FUkDuczXmU2VUj2UDDLlpzBVKZbn16YpRI0ZolJecWG9mM7NOXs5zxNBMyMMGFsVkvjdK
H3Teaq7BYvkVOczMlL7PmQCuDkGvpys7GYaaC8vvd4XVs8Aq8LTS6uexZP7bbHsODStKHH6Q4WEI
m0ZOZvMl7QYg9s+ZcFrwjK4kisMByuilRO4mIlAlaqj+CwBaLua7iaaGIuQPH0jZNNPvInYnS6dC
3W3KVEWOu9tZHrMwAzj2DDbTj620bZBcbEFM40jUGczjxLPn68nqmIBWMqhMK08I6XfZzQDVAD6H
92Kut8Zae6hfY1bQpFC5gb7fKd5ePAL8durEMHO5G6Kwll98m+32F87L1M6ooVS2wRb+uzsuxWgY
xDkQ1RaILc1YCJWNEgLiC1Qr9EE7exg/uQE+beFzirpb+NumtlapM2WE0j1/Uk8KBXx7ozFvHIvS
9BM/6jBShCucXoLyKPoPr9xI04TRho/89q9MVKQe7pe5pRV5DqVdnQLXCPMwjEX+9/NkTDzKmuJf
ac6lv9KR4zbsEYkiqv99ynwvdOTZp5DNbajBYl85vpcWUcc3pyJr8j2sSZwcxT3ZBNmFG27NINzp
/VW33AsMH0VvXfuxMtn4Kz1m0yfN8h1rQrMNkCdVPwRkU5sfPgoXL2Gq4wSHOAw3GKN/R18himpp
l6jL14VOpk8/jA/QsFd/fabS3GheWqBqAi77RCK8djpuy3GqiEr6A48aDVJbq4Buu7DECvL8nAVW
1/i/ABfeDlr99nXYmhTCq0iHGZxZT+iXEkgJYVlswLX6fhTg8Gie/Wu48g+n9exUmQIj5MpsbFxC
zOoHckb9Wk1qVjpLr4/HW2IMGVTmA3Mv66jwp567oyc0KQmEMr62ttjTC4PYlo9ZoQRlq319XD0G
dHtBsyxO1bvjAYeUvE04fjeght8S97Ku+MWDYTPQy2duCOhus3XvtRwFy9BMdvfyMsHt7HhSbw5+
Plv1psJu1E6aArafyehuhQ2FSRK6HWeDtosEBE+PZHnRI+KErAkNIR9htY+n/NZngUMmAaA5sRlR
kHVgzLTmSR8twQNrAbfm3R8CKjBfnEZQsxhklJVMR7BQ86KeV2DG0ulTdmH8QqLNHwLQDnZv0or8
NBnOeDhIlXHlSxgsR5NkSziXTvMnwwR6zz2pqWCBXsqDfllUwVPhyGzKJUzo0rvI9Ojn37SNTkRQ
u3dyy7OmaFLHiC2XtcLHeTI6SkLZKNctzVIh5J7eVczPhSTZd/ReOJyqHzv3O9ILbuc7I+rtXd2G
AFn2REIf/UGuH/XUXZxWQlNv7km//L2Mnt5xyrr6kBNNncO2vR6uECKQS5QIiDY80LFPSHUaEo9k
qLI4qTLJVCGK/36Dl5C/bXf2KQcvxUx563G73vEl5nSoAiSRm61oL6imErRdvFKy1h5r1IIh7QYI
5dTOZppZcw1L/5cMhHnV1PNWG9h+zsrIZdKQNY5EGudRUGLiQVTJxaeny/KwwwD+hEmYVIP8EcPN
lvUFODsOh9ohHgQpx5UAGqsJt7qFmCDUtUSoD3NYm5N6bpKXFsLRWFFQxtELk3hGFcO9EQjz/JS2
gizqZXzpPokr7Ni1IvtF0pF6BmyzD/Fn2V+c8IfFgdhQsGSlSbN5mMR7b8t83WI+qX/UVwPNGU9f
JMUOWVNNenaEEXS2YH9E0DLPoyznXALd6Zvu3NFjpFkCN7hSrBRRt/19xc41BP1VK51KJmI2JOQl
lg6tPuzYOGHbiAJu0paBJvd/aW7+Vn0GmXDJNG6HsSJ52b3G4nd7Ibn0dIN8/VYQ9tkZfg6N7ZM0
fLrjt+0bPkWNvjz9zST6bpGlxnxjnbyPKqSnOgimLccQ2iwK/wfKpi7HfeQUL5/JyUhCmBXrK+x9
p4ZqqzenMFhZMfW3IZLZdjdJE9Xn4E7vIXSnWfUskWU766nl3q4DeQFesb4E6lhXrbNvLc4jscRc
bHHXWGv/tcADFSoy0R26G3Bgjxa6dVKujArW1CpVsjf+78B5GPlosDPAVPHGw4vFDQ0wIQH1sadi
bwyo0oIyMx1IidlZJTIritrfLviQFUFS/hfCxc125qBM13hBYFSRw9wfafbAOTF9hhQ0xDVHp2Qv
UGgomMigIIOUTZk3sLf8Mj2Nh1MwLyfIRUBPdeRYf5m/wy8mugca4dp5+5f6KBXmjw+CdwcW6jA6
DfpI3QsZnuN9b5i8NMXTmoLVlWdyV3Vs1BQ4NTgWkWizFde4LJxHQNgQ3D94NKDNwz2Uh1r5h1Td
stId8IK0QPAkn/LST11XKUA5zrqDQodYgaVu9LtT+HCJNx7eclFlfO5ayNh4vZUa1gSo+evMwWCJ
2xUMyB2i0LsfFLPjUo/ZnpSdd8N/JWyoRiNolqaoKY1PV6MPZ9JD/D9CElr1UCNeaG6VVEIgthaN
rXfu3VNcPuxRXtc1IOC+6KOPkJzTq32RjflPRbJOsWuEivqcQZGKMZJYQg2RPqpGNvGAYU/EyO7j
8wi5Za/yaEdCjGgdnSapLV/Hid98LaSdeBjufLAX14AQ6wXRxvF+uZN3MktxM0kPDmSKEekRhNgm
BqcR7vLMC1oXV6sMsQ4pEgNqaWKjYZ6LmWgINairo/FhYVnjpFAe2ekcf2eycJ+lXwIU2itg1aDJ
eqrLYqajGmK/KF7WCprqB+0XwVQvfCp95l/b1v+FaFnw/ppV8ZRSxy/ab3bXENidFmGBO+TihLvH
qp5tuAJn8pRN29MXW47o5ptuPcIYdxYdOiY2exKLmktBzPbaCXRebAV6YGdnJJDoWxD7ReunDDwA
my9uUBKQNyKwYOE1LH00ygp6nfgy5KEUGN47BH+TejfqzthCuIW8V8Ozy1WqdQlB1hqk5nhPpwEK
/b9shmWQx/3uN3PBz/dGRHXNNEXQInnFmiJFbsQv1B02AoMAMM75W6mxk40gFYUct3aDWE4wifoA
uRG3+mPuq00xC6SvOsNB3FZHyCI04AQd0YNTgg3pJEALjcTTFUCEtXxisKax3uixPw6ES4VrpYcs
Uo8KuuYldfTz3ldT4+l4mkEFrHdXUDgiacn4PpOu8BEW9GnTjpY52qPSbshAsJX6k0HjQwvJxqk8
WmQ8EkPDGS9Ms5kMiMvaJA1vu/DZdDEaKnNLbGYyAEjhzvFJ9bv+8fGu4XkGa4DdhVi2gFI5ukJ1
xUE5MLPFdu1YddRJpo3wDAPeQHGNLxjEz8Tp+QdPgxSapR3KmA+kAAEN5/ZQfvlxvng3EHEcTrR+
2Ymiva4NnpdHD0pHpLKEIW/6TkSUITqsOgtpdab3FyLz2W/F+tQM7Em28ffHnTV2rbKIktXugMMw
zswq/LlqwxeoECEyykz8byvMzHksn12ug9RryZjniyHYUZZwolz6zvPIup8SXWBRTYkEt71Jkxyq
1t5g/1v7mNRTSJ6P22eLzM411X8U/SDDYtPc8ISPww878LMmslrQkqdKyggUX9Fr09YSPVWQ0nD2
bRQFe533IhZSZsNE0bbkh6lDBzGtEWYyCiYAxSXaqg/L+NnqwAyYTWyo53fhLYc9TXY3Tv083xPo
LdHSvAKjfIQYZBAHGFir0z7c0XAujVR4NEXlYr2NlrvkLEQ5hLcdHBiuRZ0XxvSsFx0soD+0m8H/
s/MkKLZE5DY0DW4bXA9y/yqjG2iBnTIhSKu6+/U4PWA+vaYDrTqKvbruadV/XnMKu/o7VsznCGcM
360xovwmm7IU2uk1j0/Ub+Rv3c0sH+UkgoObm+32SClAhQfuYRzU+xsFhXdyAFywpQiK6+wUvom9
t70d0t+SZI2nzmNegWXl6s8FUXWjYyjb0UQhs+fmC7a7OY03bdJJyr4BDTXJv3iNJpKEk9vqVww4
q8y41sHc/926iwM4hN0PlFdy1Ck06X+OWYr9hvw5V0yZPiLmRyg8iKWClOuhSvwLeKvMOqxdqo46
9Zn3i4/e1ZhGx3jkLaegxKUfKOjFgzS6KPRN4ASc3DCC5qYkxaK5LumcDVIoCiVyYbC0bACxVfoS
kYmDwKSucf/qiLTwSTEAHriuwa44/98Ks4C49X2cu9qFXroBTJtgSBZlaRxV90cePlM6CO8QeQo2
kfuoecm4QG2flF8cZU7H2/zS6nmLG+OJWrj3E/Y3kCGuhFKUg4WDJp7FXbqQWZS4GeWzcZ8YW8TF
DLoSirVpmVwcSnYFbZRVBYBx7h/ArajhluWVxo/aITGpT3h2bTKG68W2u4j6uo0ZfYceZaoBiLwN
7LHZU/lnXv5GPz1eInbkmiJbEm0Idns5yXKLl1D1p10TdYx2ev6xP1zMUETTLr8sA+kvtVUJ3i+4
yGTTsKWimFRW/AhsdhPaGWywqgxG4cBceZPN4/AwTLtYpcjzYyYCVl8jGI2ZJcJPM7J7GS/SKr7m
7jDQGorvVZb3Yw0tvUeDqthGnhgsl+Co3WIu2Y60ukt0epa8bJ4Iu7eMUnu1sfR6sAzw45tKOFBQ
UDzLI2KLjz4d38GDriewRuQ/JmmvHlu2MPc4zvsf1Gvx8lw0aT0dxdmDaSQTn8yjKys6iT+F/oHT
5rEGMF16SNYdqUJL4hS5SaMxjPoKw7i0vlP7TvQCsA6UdzL9iAba6L50b9/B8hO+zQhjvK9m2uB3
Srx5B3BuCdRsKxMSRUB3UmJESmyZxGcQ3Q69k3VpCS33v7IouF1jmySJZBTTx4aeLjM2bSGGxOsS
VWMrjFJAFwvWH4lQxh5/mf7NxUBCFA4LCP1Cy3QJt5YeXhhU4hl4f7Ipkw7gro+7mS+oL/1n1MUE
fnDQiCPt6bL6hZwX0FDhdBft0nhwBZXMNq0GBca423PvhL0NeboHhsKrLOCaaZnYyXAIHdDK+Dga
KK80Lxak/yfOUByYkomeBMT1W0pP1z5U9LiFvFhUm+cyBJO5LKIIIgBps1vRES4kDNNX3LmtDK+s
4mmTD4A01C8Hi6EJNYkjFFKtmfdjTo7If9Jg562YhvVGpy5dtjwnSm53YgrJGDiBeXxSyL3VbZA1
eXIvfkIC9OuC3uZJfNK2e7P6RqGWY79UTZJ/gvoYXxDxlJlsMUYg//IIEunrtbjiWfcaJ1/VuRog
uVq83uWyM/+OczVMSlq7g2CoawBsiBXB6DnNsrbiipaUyIaSEvcwxUVG4dtkexsr6q2sYLHEbTHP
l9vF5DimvkD8AzIHAYsxsPooqTMcEMLA4WhcWAPmHvbXrSRfbf3RFOXvjGXJKNqriIXhCNaHaYFP
zUbNMR6aOnmVJA6u8CcvZYukWtD3pabCg0HHy8azI4D7Q/uqW8u5/ALg0i5wvaaoM2K6LOqKD8yh
U+eRoCJR+cZ1812Wa8dc/sH+9aq3xwOb25LX4fYfQO1Xr/UcHSvg0LbVs5MmXob2bN3thEYL3oYA
p41sviSrK9X5or/vIfn92IDH71ZO+L1Xrx2dUOXXHUmLPdIcmzIMhkr38zzGb5lM5T2YhAquzYcd
Py81DFbpIl1inNApcnxxuNSEUhUNFYL1vMNMFDHkdvkcLoEIu+ObpkOZEvvrdcR1MifvjZ/1g+ar
850BT6lbQjuKbFhz+2Z22tGK0s4lvuP3m07saqFky/uR0uM1t8F0jwsakeQ7iLfqqYyTRiDcYLZw
8u7EffHuHMXkyY46+v9GnZLrV/Od3J77fSLxG+BFEhvD5IBwztdQvs9Ehle+c642km6xZYh8xdfr
+UykWeLD5KfcRJTuT+XfywLlHb99cU34se0HSDDq60fJJzKIVmiPN3/k07KObZE2E9Hov9iZaDNt
BGWCK23f6Mu8k8vPOfomBSSyTVIVDv6ARHeuAqOyevmySVXx4EgNbtkSzUatYu67b5bGSQEREn5y
3ePclx2ozNEbTsVO38i9Ss95D/5SAYKoFQRIWXPhajX8k1AlVFkDHWbNGkA3td0SL33EEwCBtkk5
rHo+iyyEvqsig3mkUCSJA+bBThOJRarVgVcP+HbzKwb5Bopmeir0P/QLl0AUHrAramA8tucyq+Um
/M8VfwNPl2J/vPCUfZHMsQmPtOm6Iu1atRBpth++NYl2XWNpn6+URp6R2myQ1+a2dMeoXUBth1kB
5JBWUjyzqRe/wFpKLb62UzaDSuLmOOkTyEsd+vM3TKcqbFF36/mRkjiZJGDSLf2IoVtEstXtl4kr
A2EHPHLOOxzUC9CpZ3A6QuLVgFsnA3gnYXlXA4WgAVhishHLpWHpM/MtJ11h/fRsbjB1ALP0WB09
5NltUlxDFAahkR6K9QL8S6/hes724f9rsY3C9JyF5oBfCFLjdR9MdvX0hol/M785aR4RuDJHoXZx
9LicSkOGtdS/z9Dk6KQXIvLwuGQ0i4ohjVzbU5AUKFQllrY3batzFevBpFp8eR5VWRA1LsIdAG94
n+SX0drLd7f6vuYzidiy6XwqQyDgrS7WlNkFY0NlG2pKO+Dhdp1adTQKX9MOOgT1MaPDdvzqWc4p
E9a1Eh2WeTqus7I72GAIuNFjRRZaoNoi0M+hcMOqmUZZIOB8I9huYByd2j04BOTXrwAkO9UJQzsm
d/pEm8mu6QXc3M67CpDXlQEQndUEpCE8rvUGW4LtA27ExxZFI8KTgI2jlfWjFkdlo72Z0wMpGCpC
8gl69tzYknuhu8PnAD4xrjhAZo8iMwCaU8PXyrYFiqN68qrZRdbLFAQD8IodO4fZTElI7G2DglTt
vx5N5WZn0Am1BvG+bhjOxVDpq5k2uAiOjQGRHmA02grNW54xR3th/VJQ0d/Zz0FcnZHJVBwgtriI
SjyPbBfu0d6JrhruriQpCM6n1SZUqjy+xLOpPQaYv2+lCt62XW4+4c5zsWFJRK6O2B21UxWdvIuf
zlLh5V4DNa0jLl2DNxs3GS6MFN2gW5MUsSk1jhBWYtJgadeYzDF/2ZiTlJa6IpytNJxCwoLH1EQd
bMbd5RLSYgKgnS/hqECP8u0uQSxkwqiEWzowU6pTofKnrEysSscoDikw+pR0rRNCGmJPtTh76CEu
MaOvhk0rYjRZViljl50VaTnulydQdgHCoE0QwoWyKK3aQFW55nVT2N3zCIvLYuhXbu9/O0GxB/+X
lK/J9lq89uhfQjVzX3mN/sixbssdGw7lPV7jySF2hg+3PbldnDee6Px5bvQsHqeVqkyKK7tZ+UL4
gDmHW6Wi00W84MNgsGJJSisDEObb4AS1idZgQluU5xN+8pqFYLg977sIunF1decFFz04FxhXLS5v
rGfeD4kZsWNvHq4znyk6T6PV6Wn+Q8yFzTpuc0NkWndbMrqpK1dQ5qKfHhCpSRGI7yp1R5jGPVQl
eQZUldOU7u6EHqChN0SiQ5BWkASeP5gT1CHEphSe4MQc6y8bH3J7vD+BASIRz8cmNI3zm1m8ABHQ
i4xwZb5B1f51bvdoavfZyXFHRbCOFAQzZVSzjXQ4GVnt+RfnE8bH5PgIVEO3ffvCDY6CNypzYlW1
qKmmN5BhoAMCeaZmZo+PifmXzLcNjzAkTRcQiK/CQxsZVfPcjcXOw8p8lDeu7ohiPCxOPX6t6kov
8+si+exj5KxOaPRZQuIpZhHRZrfYichwr1IMHsmmhmnZ03YmBZfm/eJpDuMZVOGClygTcUJuRJsd
m6YiuBkxOi0lo0O4xiHTJ8CEVZyrnhda67aPX1VR0zzDCf+CLWeeqzCfcNNfDY3xNsm8+3rc8REf
PHTcJoyK8m0WSyWD9r+7Z5EQMTiZOcG8KzxL7q8UHYR8H7pFZGWYUQ1acsLT8zSAL0qWQBxHopSZ
tHT1djW6fiGTbZf/WvSE4OmUiH7v7qx6qxpZAMcVRoMUL7N5LohVNJfb1B64OxQinkGGZ+GJdG+v
kcIJ1sa1A77zZILzcBZGAi3S78Ur/W8Szc+JFQ5lu3WVgnkUBMvWTnoythn4/MXqR6id1dSlixjz
6lsCKRvDVWx8PRfbXr8nNDwi8EMO5zYeN8tFKPHvgHM2XYVLRpsAwHjxkIQrkklIxRL1Vl6M5WDs
MVr/mTBDhCFBB0leR8WAIc65alp2//ZgewyS2zQv6h9YGowYJq5olxm2Sok2Y7N/DCC8JUIC/t5u
VFTuabbL2aiQqM2rtkLYUXoWx833kEAW2QbDaXS5SvIy38fJiSr4/KlylznE2+AiQ9IuNEXzCVK/
3noV6RCGzvdhFtkTOqWy32vUQR3RBhKyUDs1nNxRAbd6QjBELuEuLjjXsqdgt9YGc76Oe5vSIG2+
FQfAh4TNLxXlLO0PfkN4OToeZMe9eFCkyQ6ccOPte41wD+TTQbuvrVpQ6cqIGpmpdhtdujbtt9Er
pZUIlPhJX6h4ectOSSL7vNg/CQ9JcJUh6LPwzlOpOsYL0+cZ+lh5b1x/1r5ky/hPsNpPzNGlo3zI
M6SWUEncAe6SzRYvkEWVAr+meWG3lGxv55yy7ptlVk1i7Dq2gnhw+rTRWMeQJWRVmgudszTp0fRY
ZVaBSSawqdRR3VRv7mb0DxMQDcyh7f6sJ0Gex7Q3VsMFAJ1EchSCFA5raOqenk9lpUHSdTgE5EFP
Rcu7HpWXBQgI/5wRkDUKCz37rxaIf8Gc471bvjXE4joiKBLU2q2Lc1ADqCsmJUaUeGvJz2NWvcOK
uqAmT3rekbW9XLS5K8+2Qksvi79OkhPkigAkJz1Eb34mUlDBG1+l5kq+9Ujl7U64MOGcG50JW5wF
NWybqp5QD17Fra/fxbpoQ2ZK8YQDkWAYuJYrQC/s0GaL9KoI3XtgFy4HBad7ltfYVmBg8Yza7GeU
G1wnX4MKWPPTQJE1TvKTYuSpce5nbpgRKiTKtU7zoMqX8BtgnMRnGYEzlsx8arhG6uXW781+99n0
DJWyXrdFMXA84cdvlM++3eKvYUvsC49RzjwdWVfo7SOQ8p4jMq/zDiFdwdaKL7eD8sA9jZOUjW5O
3J22cekP8xFzpdyi6TV2PNKVwCqqdNZ4hnb7ZKoLmDb7agSOaGeGTJmp0xkxjyyGmaeb3RaYkNPf
NGk7L+C6w1sDKjYSHACDvoxRgwELfvpRnZEh0YQlIYg+rYL5wOrFucrkLQw5rpJSf2giMNvo42bz
ySCzBuAOAp6IuJfUTXNkpHbaUX32rBjJXAvnFjpeRvOAj0Xey2vbcosu+ygzll+S6dhVPz1IM4HF
g24USSGg28Dv2d674iMU8mG1NMtDbJ0C/n1VolmucAZ6mBhE/d/Dm8M77t+9ZBx48hdyCJI5d91I
G3uLDxmxzp3YSncdlokYE5iObtBqPGyRhyEA5u4Jxi2/slIaAkIUgENIJF1v3xeS6ewuVP131YxL
rh+N9jqlF9IcI+XCRA8gEwl6ou4Cim3gxQqrOCICtGm0mSFRUzDd5YWJb1wpiTwFxQV1xN9SEOAT
0VUsf3JxQAO6edJk+3ktvdWyPQ15ppuIYFo2mvnFo74/c8JJlue8upeieDhSz8br07gQSKJETFh8
/dpfYAb+zRxp8RQXM+Xu0lfUOSAvJ2Ml/Q7JqbmTOROSY6fMiqIpjVKv26cdmih0gaOncrhJB7ei
tmRfjInkbs0owWiIeF/QvDJXzRJCYC3xKm425Hca0Csv+s8d5A2uRPOvYGJFNPMa4bLZiaELfpRq
dsgWeWwo67k94uShxtlLc/u15a6Ajqo5P+yqLX40miJR1KImvsAsKnrqvsR1xOxDG0xXgLVfdl/e
rdVeT6PvJLAHYFaCDqC2qeKUCpOmG+svQ8/Pld6J9wSQVy+A25xUMsWKhdRq1+pEmwifReKfb/1n
FHq1WPCV0ZVVFLA4pc30TlAfzkYJ8Et4bYnkNAb7kefsgXh/ArF2a7FIZJL0F+c0MBBxh/Y5QaZF
TZRhLXSnrE0Ld6YYIfWUB11CCiW8rBu5oMUwd0rAZ+sl2LGypilA9ImCCZa/H+JghaSIB7jLEnCf
H0veHmBcr2UdMdUGiin3XxND1lu9NepvghDAL3Qq9HRWBlDVVYNuUCqJe7o5/htYgwyEco7G6+ut
dVSKNwp5NdlviiKKXFvkGFIV2gKCJkEP4K+6aBgBVPF8dTlWk4D9Sx32Rw8FL8VBZb7OSCQWlD4B
OTndqbkVbap149kGBob133qVf3JaNj28kJpjAWPeSO9mzWyxaqkyN/AT87DcfKfUM6LxQj5Zd5pb
qIlwH8pKlFd4EknQxUyrullWVy0az/DnaVD9GXVLJrk1t6gpL7xwB069tAjogzTNLqaNfP9cIoBk
VoAWcYkOTudWSDwVVRnkNG9zsN3TrRYwhukoodbxd89Ou73kJOBFiMpFOvArdylgrGYGnnuLhm29
c7e3daAlraXSD8ErLE6AhAvkLusqt5A7bq8c+5GYOjlYhB/SQcHKAM+X0c8yES6umGTS0Ik1l7Nh
mo4Kt9XmqWhBmwVxk6EtZyy3PBGLAhM1p/Sy4dUumea6oIfanrKT8+RvJiMtaHpXRUEHy+83R3na
TpbQqJfMoFbNIuhFtq2trUkAH3rja3cR6Pi1pb+9USL+B5J82kNfe5KemzmdvqqEjAlhMhbf2N4B
QSE0hU7yHRYCKIo16L4DrrFlykBCqMRuiFSXLg/oHZq/rpM5ZSgeAoA9k9hQ88uvRGvPeg0Fo+Ai
MxqO5zovGvaYYE/BIp7Ur6cmIbfMoUzQVafcBkEaMtCrjF8OOdXgbg+fPrxHHUKM6fZmgi4OWbye
Ax0Lp0dulNMnF5RnqNUPy0w7dm7lCaBwaZe7b6szdTu9AU1aMwMQa8/sSjdf1IWS4orz7i62pIeR
CaO+r0cTNQOyl+unUu2YYKYk9JrGIjOgxe1SnjCOh+ubRJIhAxRG0MJ3bmgYyUqgB2R7Pxv/jgoI
UUgP/K/RzKIycNChuT2/Dn6hUFYq6NX48xIsXjc8DaTENkI9RqNOq6LpBm/SGswP1l7NoEOcZFsi
qzJAQy4Li9KBCcHfhTd/GEwsdhAN7sdWf0llNpWXM0yHcrNJs0Dyeh++M0Z/6/z1oEZXtPbsRhw0
ZmSIQOVB8wShmgeb5Q/MkQxRZwunKNn9PFeoBKKjHW9p6OsrejScEiZ9yUzUzdD0YLOEAMUx5wRp
pGYWnRlvmuQc2R3EXQCYjWtzs7wQ/qu+/FnNtkVn6pAGeuWOZWSeqTgMaYTgQpOUuILdKjQ9QHO8
uxsFqT6w13zl92QuDbr1SfCIhR9g+smnH3spQXynE1KZ38tFyYtWi4fj1lp65D7aaFJj77Rb9sGi
HU7Zl7pn4RIx64OCXtjACFCSUADCBdiVAf/E15Vp5pybYnDRbhUnHHMPAECm+oZRgKAilMOCOCzs
7ySQLEmaFP0wDaLse2kkOX3T+tQBmJ0oJeNoQCgXovxKWkAzefObMgufkUIJS+pPXQgdlRDHe0t/
6yHgZUh5X3rZK1FQU4kxNWFrlP7ZYGRTv9V6fOm9uUFIZvh1nYAF1M/DAtHeqn4MCamFAA+GsWUz
kBEPAihZt029oo5t4+qbQsRlCNqoMV9xNOx81LFaljsygEotc2++UVRaD0FwDdeobHqKRv0e9ghA
vie5So7MVNgoou+Pd8JeVfzqJix+SxgE4mEcpSUCCor56yDHif1HwWIxV6Pfb86/xU3R44VZVZGC
j4L8P8tnx5HIpcpH7nfoJ6lMWjH15sNLKISVMkFoDqfARak/Mx5eWnvogxm8f9Hz0BzLahMCQYk5
YkVwUif24rIvinm5to945EgbrVcHL8eM0N3WfZMQhYuX9nr6pCh/EzaXZPXiU3w07uD33zP4Ogj6
n/0QVV4qvN47hGcxdKqLvv5m5sPjsx2dJzva7sMHIEGty9uHLUBt0z4XWXb2QONsYaTQCuPieT6K
aydL1BGe/0YZFPEklUJjFjrBSQsmeMXrG7jjA5xcFihpVkww3shAV8mLNBirY/iLipzWTVU5Ch08
AzHhKVJJ2AAWilIBxxR6KI9Tw55bPCZ0rl/l8/SRTAOr/dRbpJ52mdKgchUAjvxcRcEu9z7rvP3W
Q9AFUd0Chuh1O86mvZgUmrYeN+sIavsaq5Rq/y++ZWKMFNYgZYPfuyfJZYXN59R+cArfa+5dHv8R
euzQTKrxsordmcIMF7IoEfsAyiZB2q4BBvpuIBo5eabR093zBsy4BpuFOMxUc7Fzz5UcJOijItbi
PDtrGBu/44NYrkAIzgvQGEFkaC7VpIjiUbegsd/Yh2fMCOr4LO9629RSKLETDQqWT87CcO5QtVKE
rJ9FsPUnlHtYh/3tRbfSWVlfoCEzMbIz2hmvNIzgnqI9ClU9usuhFDd9/H1B1aFCwI+R/8MYtU0z
fTsEgimTdk0xEtCpVIyQVxxKGylXESRgg4TETbZwqa3FAJ5zA3tMBHWjU+/T50ejT1X3lq+bazmW
QH6PZt6wpSSOFkvtVSWjlk4go/Kj7pSK7GOt5MvnEDofQklCMrG45HIDnB8fzqWff1Zq6wpXd8ov
T/Jd8z3Qe/nY64NrquugQ1cIN+g/wLIfOSYrMOc00bFnapAxNPceYmHeTKRWJ3qH29R/Jdhx0YJF
+ichVcMb3Tbx+VGqM4pMDC2iRTrHjlRL5vndW56X7WLmC1YxQ/dpRNrVIyh6/+St1fMJ4fC0eQ9s
vTjZzGpl34drQXdJrxfHYk/VtVE+lUHP+wqOW4ATw2I1cHYjRRkY2TowW3Zu6R+DDcWS0gw2lQ0f
4iPPUVQ7hnWgGK1Z0tQXetOly4kOWame/y7UZOwVjwLYOrRriYZaJGDyGswWJbGXBm6XliDaFlnL
QgdxSiQmTtkWzPHjXE2cTWbn9yNzmAvJOgvQzg2g9uvPVUFs37M+mdu9jcg3+px+QDlh61m0ZSsX
IlVlKIfWhB+dMUAYi4FVXqM77PstJFggKApS4d30aNEpB+kDL2YVBNjUdiWEOaxEV9Apa1Skdxbn
kteEZtTqdfRbeuJRJ7lS5stNMPeFLiag9TzVqFoOSus/c7SNhE8U5G3BqXcPPOzPLGZRSFVxdPaE
oB2dvpB+JYX2kurlr3iSoqY53DJKDDk7vEtqcXMbSgyAXbw06aqZjAYfkefZiLMiH1oOmyVaCLNx
5U/nelMBnyFB4zx7/51wzGMnrnRtvGW7YyqyylpgoZu7GHhnV76ocIoiRVcGlTVw30WosTe9sdGR
JLmlRWfLwwhBgpppyDxnf2ykl54zd518LlTYfxuegI1qIhTfs6FL9tiYdlxbcYvm7cILqc75/gXL
lNlRS/SZsVcrJFLSp4sk/vQ7/iCxG8gGPHx9HBor8ogM7W2E2AccwNHweNbplLtdiPq8E5JVBpYq
U02OjY0K9NwNi+FK3OWuYeV2VeWSxYpyW9SHHrNSNMRs0TPXZdX5/cH/YBJHLV3M/iTuMFRskV/e
Dp/lqAVj3Y4JXdQrkEIlmj581FUENMD3MlPNiMXemU+L3OdUraiOSa30GMz4FaCTC3mFobfAY7gd
Szk2xAggv0K3anCKbPsM+dHpQd048GW3PVB3aoTah2FyDeDA2Mp8hgW5ZcNRwNzVo1608u7VmdOD
uKsT1UUWBlsu8v97a1q7I6z/PcxZ0u8UeQePJEYkxVaMy18tp/3j+zfrkq3B/xJatepBcLoHWKfQ
LVaX//rkQn3EEK3bOXGq0Z93c92KvjkED33mkPvUsWefgFUda3D224fuQ9QRB9yxt6kZ29vcJmm+
CSHybMic+4yzkyjiTCgAL1Nbdwmron1xh7vh8Qixm7iVKoxQC8y6L2mZyEpP4aNX+m1/nIal7lwV
Ge3sOhB+POv3IAwzgnIp41zpCOQyO79Elc7pSBV/UFw7lj69lU0jJwJ0WI7gwOAi14EJFk6o46Mr
03V4We5X44JUGKszIrjZsMInGGf5sCAHXYpP73SAovhm2+/BTKwX7Xe+Wyxiq2oYH6y7sQiX5zcQ
eHBJIH+HV3e/p6w305G9EH2zcZJhaXjaIg6EfKMnTp71tcCXImmy6S8+CYYwgQa2LKrESidttZIF
6bqE3k037m9CNuCBuxBRi0W+pkPO8d82sAeLclc5HECwbykR2Whfx1qayQZF71a7e95EHHEh+l4q
w78ZfDUAXONWDotjEi1/HUNDzxwb7r0XI2r+YKgINSlSobl+ETMt/jdMheDJhnEoL4o8KSh3iwD/
EperN7lpTWZAC+U5cVDb56puAftUo+OcF1pymGfTMW7iGY0M8EYZ8MGqkN11GG8AahIJ722mCuZt
G/o+/9aNA3SByrsiW3K+sJIC/xg+M5lV6sl8RoahTtPwIu0PEW6QvTCsZBavJH3y06YHYumtHjLf
PKeS3ykakC4gdF/e4owp6Avsr1nQyFXCNEEehBDaZ2HkBJ7qBuBcxhgv1gO+GJCqYet2o5RAmLdS
BEZGRskW022PKejJr48fesaRSi3F2c1o4DTjlpBSj9YBrJtRmwCYPVTSnTAmJFgPSRkaH692v/p7
tu/+9wUTguOUoUh4uPXuPY5gI8pV/DCoiY+9A0/FYafCh1s0lk8mSP2oZ0cdsb+MPn91ckMQTvgw
Z7LtKVW0LUjkqcZiToJZc2H0KmcN6m0Kw0heCPgdumqzIxLoSygWjDTuds7y+3C2J+cfeXfn+RaV
HGw715goEbU9mHkXI+qHiYCKzLQDU6T+os5JNGYSjb+jvIymJb7MeOxfERejtVKTZJ+MCTr1yW/c
BPyemlwl1udUOLFQ0XExqXIaiU5ZM/J2ng+WJ+U8r88hOlx1MIP351Lm7oSHeRCh4jPKvhPcPu50
HdIjNl0DVL36vgKGyjb0nF7dvL5Y4dKgsBahlxM6NGy5gCu6uuY+8VfWUj8DgC6K8+vrXtLFAVIi
Dut0RnfuSpLIBbMo2AoF2OCRdCo61RK0Cbe/7c13H61x+6+RoY5jUKe1qffmx0b1Gc4kCqtrgRRR
Q64dnL1rgtKlg5UyUO0qADYNc3lApI+QLlOxm4LygoR52kLFyRxw9/VtSs201B98PDdA6e/zln4S
m5DRjHjPJ0JJTASqUOLlW4Y4pbcPoWymISmmm+Ca4+vV8ld9PI8RS454Gat/cqkPDx9HOz5s+EYB
EtwZbtqdEJwZfuB3I36egN+PZeUUo2Z+FfXv9MK/rPYyN9OSgpQovUoqxA557Xuedvk/BneD3Okd
3xR5oCghVaAouYseP7TktfjDU6H6MwRaGfoXh0/RH7E+nViglADp5Slb7Xq9As2Lhh4GxHZuEVpC
TzzUeLjGiqIvhO9/zzA47GtzgkccyTO4ULXa5L0xtuhvBD6n/z3a+K+1+F3fGgXuOyhw3Lbb36dY
FMCm37c7o1rJs5vePBDmX4VVScfwMcXAlTtcJySsOfOQyLPKBmUBOQiHjP4NaC5cmtgWiE4Tz++2
vEO5MsMV8lQ+zKNMMDTpqsyXtAmhPEz919WDAHzFTN0wJFb97ZXT5Sbcf1TTF2USbMHDIUksAABz
bcxH41I42r3QniOMa6HiKIxDSc2Rpu4m/sJfi9srYp8foXVnoh81EGSUrdCKjI8M6ezVNlMkztJ/
BMxkANXYajhJPPeWjuot+KV+A1qw0yUw0rWEJ8/ewNWW3p3at35lwUmJP2W6h5erk1BX73DjJdH8
i1Ej9uzJWSyQsGH1MYJj3gWhUV/n/zQtfipmT7qVw2d5c4RghnfjDuDS/GY5ZFotZbzi9FThMUBm
hHRneMxsEac7fFkVquW2rWO9Yd5MzmfMPuj++Ep6fIDx8RbNgpg19kCLxkYd+XfafsO8HyEJSE8G
eeLuJxAHC/fxvg7u7i6DXLHI5D1wm6IrN6YJQXqv27GQgidHOmRuXk5IpKoJsX793FBjiMmpxyvg
LfhMzcJ2jothDp70MhA1v/rpz6IeSaQGZG3x8ySnUDvsrlIycfLZRSEQJyOWRAI43ySOrh6YazEo
kX/Qicf6XDQbGiZ8vWbESdVfkILSjUFeg9FYZK7q7BRwSyIC0t6JY1SUZvA/LsNjOqRpE0UPLor4
M9Gn5dkDK4TXrk+Ncaet/ALPPinY5ZRDh+QL1kWlC/Z7hfjnxiqdVecBfZRhGiCQesY8BmEifDpa
HqBe6uqMHQxBPrSHDs7QRCN/gBwNDS22DrJZIA2RA6jJqgOmGEDY1hikNJcGnDUx0YCga6nu+3Aq
oXuB4L5SaCfnro/JZXGfWfWhf4/UJelloED+uKSa9lgTp/Oa1yVjS0ExSqjtFZpFqn9gpWcxmqrK
JFQbXltaunUsZbXnzXyAo30dQPsF2VWt+k1Qn32cy1E9zyvz4saNaSUbgNXCdGIBFgd9zFPlWZNd
BpXkafPp/oeNLUSuhtQr1RbxnyGkT6utYDvSna3RrF+N4TXJc9M5B4WTZDtNRIXeLiLa92UujgJk
pn7S5iFcIh6LP68nkc3f3M3CrVFRv+w6eZE3Lxi8S9cKb+8ViQTh9IHqYJh0Sj+kqjStKl4urjBv
R4VXQ4He4EWzY+aPrHvMAzAZkWWriVKrC32RVqAfOi9wzrPFzhhpoFKWEfF3AG5xC/5hEuNyo0eq
XI+wQBcRpCWgkjlkH9Am8ic//fRUW3oRbfrSwz8emtrrShaFQljskMdYpRSF7mEsoAJ6ba5JWdkp
v7qtHB8HiRfZ0LAh627UtVBHRctFaqTyRrO49fJM4Afs42maOdLILpegIEOhKPeLQy3s4umW1ozz
/E9u7EqyZw/3ylULDz1Vu6rTQZuANUQfx2o8XdlGWj221SdPgslJKTF7FikbgHRER0hzI3c/a+fy
4AvQyTxEKLx+atC6ysCyJcKG04M9eheXJ1N7noKWBwIc8dOjnTOnLzhbbd2yIJqXfSp83HVrEA5H
yPcgO47DrXHRta9k9rCHcFJeftq52c9L5nReb+YWkdakkNZ8NN+QWjg+zMka6j4IoiNY4eUw9pGO
XfxJGrFIpoVpec3finakN/dMGEB9v8F5aOBh6NhZehIk5edx3RsCdMEx6Au4FIifdiqD8+ySVzDA
ghh4w1QGCbtemdUJpl7OTH2rNxh/WgaRmL2XRqA2upvdj9ptFYjgMFlIMOSsSXDi7FKCSU0e3ckW
Dd/OGMp5CIlQraCYKaNCaAtl2HFh7d+lBsN0IVfGrdFsM6pqsjmMCCwzkEbMEy5ntR39EyRPa6ID
3Bo6+qmFvK7jEPznKKGc1ERsSx/6hb4Ehwq2QjkIPhemm/WI7bF6laoMyeZJcYQdvLRF21FExM/D
cwf3K76MncSnrh2VssxOri96VeebhqQsIDaFvCjYbuDTi5oPcdnoSOBCN3RatUn81pTHqhG9bta/
KPn5DmiR3lTZ/QIjDo7l2w60hdhBMrprEfhnZaYRfTnIwsy8uHdGMGkAQZ948mDHffSKLSskrW7I
k336+Gkyeu4jQfPoyOqKZ7y6bTUzQXOvp20gIrsTqYxhjYZ740hIInbxiZD07WRjxXVLNRx/Bcqg
TzNKcXdYAKv67QrTAMAAVQJxl6I3wftArkZmlZwGygYJKJPZPhU9aEFaCt0rrOcJxdRj3FTgwiOJ
rKwNUDNlaWN13PtETpeCHhB4+/swfurST+6Lk9iE8NjD3wF3gt+YNCn3DDtzYqtOOC961zpd32av
b33sCGePSJJQzEuqAFt9oKu5pNNwJrWK3p3ZgXY2mSSVFfYCr0j3GX4KsG5e0LBMK9CM4/ULgN2S
Tiu697XtHaXg8rWyzmIzm/UyEgEIHlLaGI8y1OdBOuDCqWhAg7GZfbBgmnAObuSz7HMAdDbQsrG0
QXYjG15RDXODHgIehIWrn3UAElnlt0SAGi2feE9vPCPg2jWjomPpw8lKdbTgOfFKWgCP0OhMZXxq
DjQqttau6JEXT/XcCbN/CDTR7Dl6924Fp8RUgcVZZaNykAVYqnF8Fx8bjO1ph1d2TXcpwDD4mLTm
H0sj2hy6fbafgnyJyxuHsOI/8D/zytk0kpZh8n5qhHCP3HfQJhFqVfu21varOqFdAn+6+DLiUPDm
R+2K+VHzkDPmGV/mE+LGk0REyrrY178yxQJyKkEB2d8LzRT8UC2UFz+OLD2FriH3aysBpOyF7glg
xVa4tY2c5mHgCQARVJOSrwd2DeLYg/BsX4pkfwRIeZpF22JtO3CvXH+qO7JaP4yfdsftwEfcOxUh
+pR4dxNLtzt1lXxS+fQZkq2yzfU2Bks6YMWMeRRnool4WC+pLDgW5I60RzD717H4o5DAXfu+nlGU
0Gp3rnQ/pcabQPXTY2lbwkPpk3Fba47gaUbNj7bfVENHUAqX1RgSsAFh10UHRSx1oHTPrc7j4uwt
oCdYnu4C4+Kz+BLJr0IFSOexnMyPrOBcON5YpRxraK5R1xh5vxJ+zOX60KR6wqkXMpxUKZpnqlg4
8kzrKyKSo91FoWD9hhNv7c8wwcw1yM1Li1pyA4tfSnyKazoR+S76RwOWgHMmMFG/Wta7eHQpq9vJ
1yf+wfpDlZqEkY5fbzCRFVAvRr3K6Ch4UXc9iMlWtvEaG8406/B+mc10nkTDU6ATJch02ZYX8hD4
g4qJ7CjgGp5o+bQMWpNQ5yP/EfMGE4J4nSA0ckrCOKCtJ5vGp/cDetz/MKlszfUWdn1xauhfA/rF
W96Zc6rPoh8qYkS5sSdZIqJqxRpnPDxfdvQ5yY4SQ40cCZ03PFDtBlvKmcOtqaWVmGh3krbtV4gW
H+JxmdYGKpjyuk/0aairzEDVra8b0formxEpsfc+Ovu4m6aVKaA1Np0o7tMoQbwn76WN4NVL+FYX
QTHWnNbeP28+WPWS5cDi2N+2L+VG14POkdfDhZ9Y+7kIbaFet0PDyJu4ar4yt60mwg9oUVeFcvb9
hpMwpVEqTlehZBwaNvKuu7jtq/jgXq5WDTXgdweQL+33IuSJGeRODmqN7/vSgxnvq2QUZJ7cW5DR
RGlrOGjf0Z8OnkXe7xSs6GpPc7XGMNHwC81JNh/WJe8Bo7zvvQdTxjFq+pFp1+8oly8chyxvjRHI
U8w6X+n1xS9KPraADzK66GhRFvGyRcSEvEC1Y5rlCA1CESx7XZ2zZTPR1Zfv9aBoxy+2Pf/PglCq
uxgkI2FsubojuPJFTngfIC0wQ+anzBxpQpkw8jmVTkoO7sS6c35awxc30zY+3h0+OcikRoSgeO5E
neoayACsmqF+VUduwNZ/IXfyr/8vUG8ux99sRX3H2+LA0rVuNFWT1ZRsW8k+zAE1Oc0ZNCSXqBWn
yVjdEDyqJTLbsaw8ERqYMMXCWJgPVM9a1MDox/uwqZc1ocjnqR75ghgseeKGX1xkX/7qAqFd+NL+
W1Q0wWnK/DhWo07iRQbTdj15SCXoPjNDMOxwnpk3V5krEh0aKLrx9ll2ON9Atfl01XP+iQ9b1UYJ
ZcY7HiiD5lzsAgjdKAjjkposUjhZ7u/vkDYitLIeCaIzxuzFnLSOXZlu5EH4KUa975pOiAK/Srvh
FL2+X0rQCKMyOJFedu9n2QLFXUymuKp5huyKoClBRMiKuLzDiBy8lDqLVK42GP9gOsBqfqG1XCC4
CaZQhq1boNcWY3GuotMA+EsUasRvcwsP8sjuLxdI8vn0noDnPwLeqcdDOODaC/nT7CVg0flFpWrn
qipCROlEE1nrz9bq/XDA6OfK1z3I2MA6VggdktFeGFwb0tbYZ1mW+la1WGMZIug/6YvPdWKtmf0j
DfzSfnujCbwC3nhDlVslOr323/qTSzVVuKjLEh56cOUjNUSWr6SVwAUk85A+Mm/rxl5Gf9mYiR0j
5E/JhG3fb5nO8mIJkEqJ/pnWMjN7ULCHQa24W+QMZPXrwajZ9MaCmQOZlDJc/Pkush5MBejvngL3
cmWeoOwR9O74fsUB1kYMh9sirqGlFqjhLgwvmewFVTnKQSEAcb/MSvJwGiGMMhMqXu/j2omf+Biv
BE8bxjH973K+8uGM8yO7Ir/rCDp2s5mqs/v0SW1GeapgFSqkqnky0DgVVKWXkTtpYuq+GNT8s0XJ
oeqPSNRmzp1Op+VTtrxSVcF69O3Yq8wcpfqYW2EIn/59eJUPHEEQFRvnB655bhRLBGuutfkgogC6
ikNF4Z1K1wym8FiNI1a4USzAa0PuAyTFWzngi8XnkU9D+1Kg+7+R0biGDYrovu0hQj9F/PN+IWni
rglR2DNnMKP9PtHj5SmmZsHpjwLF9jOXaCVyIKNRsXgmf/GdYyX2Vc+lIiffAKDZUblAtnCeoqSO
f+WIMzr3+4TIwE76BKbkZCJ8Iggp7x/VEseHQx+NKONgiq+K5qcKP6/mnhrik2su38IfEmkduUqg
0MgUuLwSgNnf0/WiTgrnhloQiU5l9JL04Uvl5F7Ltm0mBjwTo3DSXJ/uBkNajfVu+o5ErO25sBS2
Lnw5fREKnTMY/GqJHQnf0K9yHPBVjguwoErryrcYg2RzgogVBlms/SZijUWet7YItzbL5TjaiJ4+
EiCgloOXQFWw6Bs4jGNUuwOiBEVTufXzq/P18EU0wsbrh08dnoBdpoObpH0hO3TANZJr+f5NEshC
kst//R7rek9nSF8SMrIYmCyl0uXKyNYOazopdzr0aoa3SlkHLNhfeJn0AxiBgmogRhzQSvvhdSoO
U3qvRV5Zclm4H0O6lo3L8g5KQ2LDExHMOLS8XF08tdwNLokX9T2EA1SZ2xcWb87+eb/o1IFjgMR6
XiLFO8ljKWQtOiyiTD7kjc/oFjX7KWo9qzzHDSgecLuGfhkU43eyeck3JraUvPJiD+YpkoxgJPrU
DuXMwCV41a/cYp8IpADrgdgNtZfEcZpqrdGCEKKst3+jzYW5B6amPKxxV0kHIl6V/uB8+MoHkWvt
gZ4kpXmuX5XM8NXzbTE+0Y/qEhjVfjfw8alOtun9aVMw4h6OmSvvq1RPGiG9XXB13jHI+UaUcj2n
ooyWPdkZIhUrCL/jsxZsmtgE1pyMTPxgg1rlsTIgk/Bktef/feL57v0k7tMz0FCvbuUo4WzZE/7n
hPHCn3gbM+VqblSrRdtM9Y8xfxN/dzHV21aQIAAN5v06SEtTw5yEbk0w491tkVnhydxi+J6mLrQH
GYmZOTSI8wIGbw2dIAe5KKeKW/mjgD56zh7pbtk70Tei21yMhZ9SxCGKROEm+vjR9aFxfS0qFrcU
kno4192xeXRQ0XwJIzIteNQmxGtdJ1B9rxuyNtLLnnd2lVBOCZJUR+Zji6DpQtxpSw+KswbR568g
WCiB01A5geFoOnpmsVxxLLl9ZmXZQ2Sz5kTjFQV3He+l8G42dHseOC+mEoZdYBurWs6bNErtOACr
BDgYG/QoMZIS6WZ6gkit+oZfOw1lLiom/FEKygAWopuz89aG6PCgNajjv5Oi5r6AKwvjxmc6M809
z7gTuLu70SCMfK20/9C3bldEQ9/dcN3MI54EtpQIoQrHGgzTP3l2ANZUg1jM1p/c5hvkrnwC6ABc
lu77/2m/C9YdHmKnoBinvQLhJzFRiVWCsvpKI0hZWHkw34XBV/SgWxCw7G1odtvTzCgB4be3rCGw
T0hZDwGEVsBINknEnzzHkRYwcTWB7fkEz3JaTzuxxxqykct07qPfa+EHcjnocglLU4UeYzCfq+ux
izUDqXYtOyw1vsYTq49jAbaz/KiTseKGuPIoT866spv2qQZRBpTQ7Efl3+/Lg/kny1/PU+x651Qm
K+3mo3s1pKEwcyfwd9GTZfD80yx2+1VuS18Wt7lFEl1dEhBDfQhnc5sqQFIiE6xsrvImh6Mallna
m8Ay+Gp7A5+6h2r8z4jPuwGlIpRSDbuWBvA9netRtYzGdR58la1MIk9IGkIpzuXc8/xu+Cqy3MYp
4z+0jzUwk3YK4qAmO5OonGlNXzxLsHFSU9HOrr3KFvQpJBegxXD+Ifck1RzAL0cWDzwTSHuKTcuL
fBjX3iIs7Y1zsP+xBLqMgKB07a+iBKKNw0iG1HtlIVA1ksP12FuFd6uoJgfYxXjUKVC388x8iFcs
sV8pz8RJO37QVU00W2wQEdrA2jzdWy/0CbS9txiRTtDiauX0BkegR5O1unWOGlOlMZ/QKlAi7tz1
IlIdFPvGCQAsQgC/k0WPIcyN4o2Y4ds/PpDIu+ogCJxeALqAtKDWGbCSBZcYIwwV1BTLJ2CIln7W
NhlTEgKpGpwzWsH7c+qCcVNrCmf1L/rKU7F+2T6D0U2O9EsRv9oEq6Lmvy2rgiCE013R40X1oGTG
oRgV7Ov96aNM1rhT6/AarDAzKpaHGzvzycbTNC1X2ikZ4uNWEyac3xwGHwD//MgK1s+6ZHn1sOIj
LSd/kMSBWhKBThkPTfCdj7jUcjWbs70J5FE1JwicYblKPWrHPy+IELQHptvBjaI8IOT+rgoieqmN
1lBeRxQdh1zr1h/qbi7RD0/AcyBLXk/cqS/04HYdWwq5x+5LMIvVhcpM/1ruAJy/AxbXab0x1Bp2
Tbp83ABsExCBjvhLpfdG+H6m/tfS9Q+lefO/Cg5bYj0L9UWDq3qM8kWLJ0k0gKHeFik7QadKwf+h
+H/rmF+QDG+LR4uwxSj6Bj+roiJnU9dTcXiWxvcjNFLnwRr/k17BG3Lb9I/QIU5RkYgCQXcQZIXj
EJim//yckP3xeIUz+s9bqeF4yZp9eeW7xTc+u/dmgyv3F20iYaZYnXKiEwCDVtFL7uj2btn1aANA
UTwTPBArg6V8aoF0wGPyKTdJpcpJqOtjbPOLRBTk9ZK/YtmKppoogOTMLPPQMqS7rj5KhHrzElGX
uD9jSMHueJOVUrVlZsRqPxN5Xg1o+1OAvM4CLAPkqpnQEKk8vDECsnlOE9McQm/ZG/oE8Ih2u9vl
Qm6mTT4t5Mk+ImBwm5dmZjDWWnAQHAGOc0lwG6dCqITSKzOKNxm6na6ajjuvLdVwCTn2URBSBLp/
b2NZfnXeKWYP0GvtXq4wuH2Z6RO3Ik0irDzz1s1NwKYJTLRT6b/gHpqXLS3YwMxO1uaFamyEXZEC
XZHIJlq//lZeGmLotcFfvt1geJEcWPoiwOjPadeJ5AbWRpfljDgaJvOsCQ2jcpOZ8f+YLY6REcYb
5++0kQDV/F6IiSOS0y8Z1KjXC4bxndvAXkT8TH4RADa5UaLMo40gn9MBwJBt/hA/bYo+Z+TaaSWj
y0P9Mdqamgqb+Sl9VY2QeSnGmG3EYSbWAh+OgEIiSsnMoYPYGpPzR5nnhex734k0o1pbIJNRaCn1
dp4aBNhQOv6GVw2WmszwIxvWVRemSMnzdjrLe7MoCK9EqrZGsY7/NTzuClC2s1frQ3z+3JHxH5Zt
MXlqV2I8Oewd157XQnhNDPal9Cboy5n12vFujc+Hod8czdelNmp+VeELayUI7wwfc1UJJQ2AYwft
+Z7RAiBz7f1UyPUNPCpckS8BNPoHFHpuGtjLc8z8tN5pXZBlCgDLTwtKEEwOCUo/nMQbN4cV4uzx
IodaRFa01/R4yon44wLoXQbG5SD3O3RNYuvHfddWD9cwRiOecy4C4frIntiL3G72pD3nMUfHrnw9
1Fo7vsVVkxofgn3B2DdJQ1KJfMTDKDQ62kuk4Asw84ZqbhcRUE21+VDlimCgreL4WAxbVfU/70fK
g9XGUXjvZeDSkQJwCiETvN8lXiCohLa+lfpUdNg7x3dPYSr3rpcA2OIzyzQBKgoGJASShVi/zToz
eEgBQWykczw7UMGs+Dctnr6m+Mua79ilvLo0QPPLWcB1UbTp+XGHJDsV/2Djr0U+m2eL4wh9yAxr
Et5ELtaH48t6rM8m64Qku1t1eDBcXibUxE2c/6cdp0RcqEGAZ+761/8WT9EaL88VEenmU4w3rYMB
2jwGQIsfhDFeoWYYTvXufQVbH/J++P5IUALZTB9f1xM2Bqsk4bLizbK+VUNZWoRUxizHoHWshCph
3p0wQKWCfHeiLgJam6NqGxnjAigycnLBbi8X6UrNDqkg/umuV4SQNzdweYdwCckDnocbj5C1Es3C
oiWOqTEXJhzRcS7yYQRsOBgi/D/MzhRGbayDu343zkl/iP+yH+2T4topBxFkH5Vtzxm8Ds1x7Wkc
0T55KLo+bGTFRNWbA7OgXZ1IKe28fTEt1+3bl48YNFpnW0yXaEIDAEhEalzFusbN3U7auX0Mc5PD
FoVz8sUWaCGyT9VtAhcutLDMyBtnmR4taJ70j3ufXs3ev7CyAjDA8x1r16uU6cXkQ/2hCHkrpteB
+jJg96lLg3kU1H6QvXnWvZHLrNJStoo/HQ8F8AnuqRkacFkJLZR+4/L5OnbYKAMFqZowLr6k/Flb
5Iyr+d5Iw12ohcharz9M7ChnOw+LHf7Ef90C7mNw0qp6ndeaTrY9M7TY0Dvwel+ovG2GwLDajjLq
7G+xr29UJCKbt7xFvXCe4YKiU0SPw84fDjMMkumXWwnGz2461PPfS3YtKA945scgL6OSoofiOoAo
bDoGkDX9wkjd0H/I8IiIXrvUe9tGdFUMS6yoxxUnwHaenU1uOzrmD6JDd9eT4bl3XSCR+CrCc189
uzbanQ2itHWdp2Z+IvX7Jppps5LbP37vcFCo1xWN9BuMWJaqwlEmg4d3vTl/K4/yZB23rb14GKvj
bNldbyYNcfgsqDA0TYuGmfp3Dt13hwsGPJaHNzYwOqqa2CE05kG5k1Kn4F6mZD7IKM8oydaeG6hL
bfTk1epLfsB0/yFjMKAkakpBi5DOMaEqitIxwefn4AS/1VlhQh2aby98ypKT9aFxLh7X51X/XmJ0
ImdggL1th+x/wE3IfK203QJLgzwWRZi+AQGOlDt4dQWWVf+6dsEnvAlpss/xWIDoHodUXGOXkmJQ
5ZKlQNgtEuJSGzj7z4TLB8/+NgS4RU49BKh5by9RSaMHxKcsJS1eGNACJA+NA7a59nHvZthFnusz
P6rUpQW55Vu9TtGgX/mM3Bx17lk5VSROoCVwt5qTCTjHS+DRFx2LIJzqcReB4SBIYIC2utD2Rg9K
REhzRfQHT9H1lNuVMIEw60CR2lI7HVsK9B71831Wr4+UYiLHeBYE5YF9v14Vq1lcyDeKySztlsEa
MHLP4UuDlTQ+eRXbU1DMFBfj8qhcXYZXsfJvgbtQuFBFm6DTLYIJsizPgjE/xXfvNzyetsquQ5Mr
dSH7LZQiXuOACzqT3QYWLcQhtX73aTIva8P/GZj73W5MaURsM5z9QtEWFRpyoNCuGOUMAOt0lEzi
BXYddHxfZvhhzkkTMn9NoQseweDxzfctylJJRw3L2l2USy8akGOqbVuwbeXsZbCXAPEOWZmxygms
09alLf9Ziupo6lOiONrvkY0QSRdK0MKmF5+K9DnuyZn1PBchQzthd2DTjt6dXC4oeavvsj1AO/4h
/CumAWLK+g3UwEy5etY4tLMzZoD4eEXDzXumsIROVL9sLM34vRChxi18opZged0EVwVMzZyf8t+s
X4SY9zytXbzpc/4Xg+1AK3WZsG6OkqS6/1WjADjndev/LDRSlfjsxzjQSrIaHCxFcD7Sg1ThtSr6
vcz5eb6+Ue0D6iP/tv9H2Hrv4BNoZZ7OI6yuB1SUwTHEBInGVYfOSX341x+0RkTOPW3IdonBfOqD
x3OlLIGSbaX2M+PiqGi4kLb/6uK0ajI+xrw+kTJSfiyM6/5UpE1+dIA1VJpFoXnRYDmcizQAeKfk
aSzr/BcdZGZLYzlJ6CFbGlU4CWsVeY6B4n3gm4HFZoGSvP23Wv2w3TTjRhLNUl5vZYOrwti7SaWS
J1ynain5bHZ3aFYVoOynfbv0JzbCRPAod2tOPRw0AHO7WKbVrixpwRg464+LrnbAzEId5kIodIQ6
bJeNHpoVKHJTnUz2rX7BvZRwcawZNPIwQ8yc6+gU16ede4iQmTsaOTATqYaZXTyxZKgIPtsvbHeI
SQROzFVNZE7vieFlbQ3+zT2aicLgLOn1QETyfmPUriEJJERovLzd8zCEp0FZhWl3u7Yi41UikMI6
mwF5Nk77J2ihvRwF6YWKuHpSpZnz2K3LR0C8+GYODPZ9vwGtU/tXN80FyaR0h42kuHpZw1AK/Exy
LQ2E0wwWAtN0+31+wxVuBeCGaORK5JfgAF+W26jIJ4Gy3KgvPInCCgNvr7zVJexxN4uIes+eP/2F
cLriCfLOihFXQP1pFixrxdsfY/BBWCFu5vnqv8NWxvaV54Ff6tgDOQvypK+TPQFcpe34UKp/z8xB
tfUhhLUHOIdEAerN4rVDEmIjqqGd+LVcTFVZiH4ag9zju9+KFGPqwpmzHEKefAO10f2gQ2LboHOH
a9015oNgdXfPLfY2inCaF3TK6MKBlRqINzZi/ZNgg4bQDHGePbw7rbMXztZqUtjsixQnyXUuPTDc
dKGRElpWvfPuKgZOej8F/qK/OJPR42P5Q1ZhiccpztGHH9WtQi8YRwN6biNzgwqroB63VCCgFCGR
RTqVvury/oK6bq4Z5Ie+XFGl4Ss9zlZwpuOmF2tyQPJFxW1nGua6gzOBy+CC1t8t9iOIpX8DBwKr
RjaMI6URHrahmF2YwKF+DeWHcDMphzmPhWXrQgkFDQKkqpRp0R+mk+e0DHwWjwl5CBoYrIc4FnK4
KVPWisPuNXOxHIbW5hRQJCtMh3Zk2v4MVEhOjE6ALwiGtdMtlJ+4O6LASKprxfsEKkoAyuorG8Re
VhZIyHW49RKsfD/kpt7ExXpkwACgUuRDj9n4MxyIILh9cfSBX9MIWn1XKOLX90NPy/HYdmoUD+N8
p06eTJOs8P+y5aVg9q0kVQgRati4ZRPKb+gSeO4Sqcj7DyvLDkxFyZq9ZzaOdbNDzpyVUBaA6mvE
JniCxm2AaJUIDn46ONEgTnfw7QSt3ukMPOKZ3YIH7ICSvscZ90zq8X5Hf5POcY+/NNSt6i2Ms47n
utW3vKFbUhBh2mqlXTpO1I1352Xl2Z9T1u/D5sZKcvEqaDyDwYlerqAJ+0jpOs8i6H1zLW4LlGgk
wikU1D3fZfKJGjoqc5UYeh2opWisKqxmaHgSkOmCz4Ins7b7DnQ8/ydUmG3k/vHfR9aP2OmoO35P
f+JYJuYmLw3KLYjAvQXkfiHUBtoYo552xNcDszoxm/OwDB/p1KuF7e0x88tL/w3n+Hd/+lJh779v
whCi6tGMe7JIeGSFag5fq40jXIXYhgEo6BdfgrplS55zBVwW7UMC5MkP4sWEzNWLoP0z20canwSj
eeEsuStL85cQt2lqeb2Y8FoyUTF1uaIKblOhEyPJ0jX54021PfoDaLWnUW9POeEHdTKTD83Vb4lB
Cb6eB9s9gcBrchoZ7S2DfM3SG57xsXGhvSZ7gPmPlVptxUnOpbJlzaY/FWhikV6fMkCsiPXEhe9z
PaS8Cjo4cRf+9Mg9Sl3Svp19rCKsIw3VwiU6tQNG1WWAKXwsqb+G0qhUnrfYvA/wLPx9xnDQI74B
tz8nNI0rLCwRQ2u+YS4MwamXAc0i6K9mYdxQBWvoeLquLypIjHKNTMk1nnEZibR9IfsMJXAQA/Rw
0UHfPamC/uT2oqDln3IwL16p85Rgxqkh/DFt6G7ygasnTkeQ3nx1VKGeWIi88GVz7P0wGX7boe78
wcG0zbcODPc6c8ak8rZBbGouiD9VjUHZLSpH7k7IBf1MTHVSgWo2q/9SW3qCGjoA55WBe9UYK2+N
dV6Yv5zB5PDyUNVYs8m/sC5AdW73Ycki00a0m5Eu3f+dSY8CALpeVxV57RgwZ5RKlcFOybUJWMqd
x4lb4IZtn1iU0My0+nD4WDHqegsd/JVW7UNiAII1MWAGIyTQeDddImK0dlFgmTYDmbkBIGpNdVfM
2O9IpDSuztC6yutDpYijcYWhKQSvzhwp151Wzi7Apz3bMWTD7O7KRgjYXPLNi2JIqVRdMuHwmnEB
yqnfnRnqMBOPQrOFEQq78voLQx4b/4olGhhKJHyNC2k8dVbUkQ9MQZAjjhpYZfVmtKmh/lbyXLGU
F3M99MJzztFZXJksaoCxX5UDRwVdWcEDfJwbY31lrJi5YH3htoo5V+CO/G8neavoXX+ZYruNQ3VD
ArmLb2xuBwWAFPEc6V2rCXcsWSeWfZXAa9Z4oF6OdJjAlLyM4JxjEDJjDEEUjw79yhi+WkilPiwV
kXA6JPgkhalGqcM37GnWGgppH4y8IjQuK6yLxqgMbjyM3F/oLLm5JHq/sPd6dfJcWqZ31/7PpIgf
gnE2IWXs+yTCkXQvsScMAGxr6I3G+pKZVK6JwjhCk/wq1u2S2ECYZZ8EaY2eULbvweFTI8lsqOp8
Wsck/ywII9Cibpe4Nh174cJwGZBTA4hcC9XZIFxE6ijAyPJBTgr3Uo3VhjVJwWAn8zLfMKC/VQ1b
MWFI1hYHr4cKDxf3uu+jhHHZqf53ccI+sQ3mB4bKnr7PQo04jOJEQRvXzpBtDlkw0EkOFDXjXcvU
5OASsOOnKJWUI458z72b4fMriRnP2tuy6LL+KyN1ifzUG67OVQxcGjIKjDLV/TCr4VzcbTGjIgqu
W/mIxb9ZyMieofwbBHqZA8SeBPDVtKKVepKKwqdmtIJORTNPEOJwy3tlzbiycNSIooAjVimkVr10
/s0EpLYUWSh4HKogUTh1nZdm0qHDZFD5G33He2nKRf8LUSVsFqd9NbYA7dwWiBgSe7ZuJQXoepyk
DNa+oqzOVgdlsAEIoOzoGHdehAF+oRn+esU8sUVYLEAOP8/diSCPhxLkqaPjU2DILxXgfR7CnzOm
ebM9j6rNb5/5fKXLY1sDxKsV5dyUGXO0Sw3cNWnghll2o6vJJ5KLhALNHde2M7RRMltoK8WLLhQA
w/P3u8YW0QJ0ozIywgFFd25TwSeNilbTLGJ101JCPc4LyjeI1qibzU0P4BRAfhHe9ojLktWJBDPL
7iJeLffkdNDjV5TxQQBtOD6ghP5lHZ4FlwcIegnyw6DI/1sqi83TbdPaiVNTTA3FYoRdHJhcAbtv
LM8bcCUezKyhWnTLEZcTSELOyELpd7Kje+LkhtVGamBI0Em+Kso8mCr9JYHkKl9tpkwBDau8YHxI
He9WnHvFmNLoE7E+7z4tl7pChj06iUCHrzmhNrolt8KL8VnFWL5d8uTkCO6TBDCFPB4dZG70N7SZ
PRyPIYnZt1Kad2zdlrYSDmzDYaDx8qzI2BWhQQnbAN+1MW17XjR0dNk2nk6ZFBG1KyYEimZVwUKv
4Yz0+QaefdsoQpPfLsL6LOSF9GhVDmxgtGOgc4oWtqbwJ6sRbOcwaMsOEQnRoCgRyJ6NzWPTYbnZ
543CrdLqaOfUq2kLP+1nJAGkosxuRRN5MBQCNJ4088U3sH8qi8iDS6gzc5wnDAZ/Yo2ju1xsTCdn
8ejI14g6GteiQFVWXyPImWxTghVVKk4Ctwg4eZjEJrKqoePWucjwSv3bz9o5Af7tWwbVWpcIukBB
slz+KXttxFW46EWt/GDf9VTuTr/ieboFg8unaEAMgYftSeq0SCbkqwWAn7Q4Ubo0Yywk48DzTEmi
us1HOHVPnzI0Eowd8gFY0Xo3U6DQrpUlZnliU8af0uLyWZagPSsIQpQnZ9S38RRxFtI9cnXRfAk2
qmGi/gsdlHevsboXQRCu9xb5vyx/8vu02gwJy4NpBWAWulCpDWe6IAGWFya0rwWdBVgZTROk3Jye
mpCsYt0oPqj8o/qSaXacPWxucKapa6pLw+hbrK2Qrp9IFaC4iEcP0HbySq52qCONlbPC5sH3dsWf
GQS8pdFBjg5VqyoeKqYIcfwHS7SryD4HhYSzSR6ngeozBt5DfsfZ3EJKtQRTXrdQoQ7ujGn3ezq5
1uDV9wdK0E4AkpERiZqDaAiHQBOf9ZkMEm9BxwZHuEcBdvbuW1d4OlU5ImKv27HhLqmcBASltd0r
zTrd0Vez1KE73aeHxEuaTR9JMgLKe5HMU9rFRkStEl5UyeA/R0ZkDMsyaekPyMYDlOw+LKHWkeT7
0FouoWDPTzYGUfGBNuRN1UiVfkp+2XMJyVrCzOERYODR65KWGycqKnhPUANNKP49Whc/YUG81IQa
xuKJjE3Kgun9VrKYP41mZxKdUsvSvzHht5SO3a1XrnwjtfSDZ44eErQkJ8scIjZ9y1e9BTmwh3SE
38rm8ekN7pPcrTBvcGFvv8wMWbWXoe49mwuw3QqJkp7j9v8JPudBtjoaYnpH7f82zQwNIZzB+fXu
j4i1uXL58pnuZqvTDqX8lZ3KqQsxuIzqoYPBFx7cUndL1fMePzctbu/fMaKJMaIRwMTmfZ2lpct0
tUSXmFy6VRsY9g/i/V495gG7LNFHIzASY4SvqF/PoLHKXfokxfoxRg7kGygYrpqhyTCVw7az48Ci
oRXdbW5Y8gGbzE1EhbI/226YE/YhyJB4Ndn8i27H5DZ7XzxaZfU4wOt/dchmc8caP1BSeVV8YFDP
a4WKAAD1ILcBdE0UcXIWMKETWq6CBfnkSkLcHacj00csk52OUkAlrfxl8CqptSvzoBxxCoOwAh4w
rkuf4hH6hy6qfGjFRsJihkd6dGuAr6bbn7NuvMB6kk0qPUWbliOM8pLM0kO8WdrhPM/ZpkortO5F
TywLLzLujK6QQLK4IFMZC3mnwSKruCIS3oCDy+54tIKk3emJuN6v0ElUwxDxzQrPlE1aOfSQ5zio
ztFerc06v9OcKPosPbyifjZbxSlmmXltclpPRuu6LME8uGmdmZT2w3slorZrmomzaB01yB9B3QEZ
3Wg9DQm+GewMqfSdFR6tOiucsOqdFgbW5p0YKwKaqGJ+gVfLA+9WVeuUc5oUqy8eS62py6u9w6BW
MZmOQZ8sOwYIINm2rromNIU06PG23oZMxlt0a6zQljUoZBi8h9YcWhOk/3wSe8BMwxn6k9B94lPU
k3UbF1SZdoty0oxciyUwWSmQNvdCoItu+K7mLehg6ozyUv9ocMoyeWLLHMqhVuTB+LWXJgFEfEsN
VL7TeyiHfzLlgHzWYesxd+8WDvB1LOac5xYB44hPGWvBddO6bQapvfYpj5JH7AiFod4Ax9fcJhyS
4BwV/Nfbo6kND3xP6tzfrrsVC8lDT7LRyys7yN4tyawKn5HkUTukH3u35SUwabPFAmL2tcksVVot
Bef4fCQqiFLGkUd1Zy0x1eP6LKTTwA4FVmbqCxiIDQMsepQK31bvumTGb4cZSWLNsPLkJQdJQpqH
XGOFiNKAEfL4IczZYB/rLFHb7VgwYS6b8AjndcWqZKZu5e012TjzLprtmYXZ7kJZpc++xJFz7yjD
aehqVqXHu1Be2R+6XFiz7M5OyfWDjIfU0AL/ft673IR2SqG89/Lf+3Xnnw7z3UM052pwy62m3qxi
7QGkq+e5VNCcna2z1MLi/nCbANmnCPL6atDr2W+g685dibaaN3QRfUikY9S83PMmVw3AZpB5wZFj
Ng1SKZ3x5S5G0P7Ts0lH188dQ0/AEmGbdrme63gkeUpK+W0UwID0pJwet0Ls87fUoDbsOrqSAVcK
dHWW7cvKD75p6sps0CHENhUr63c7UTt40miu8e1uS+kcPbbDHT9jZfRCmpBESHXZWptD08LBOCFU
dZxFmaIRKMa91ffBpMF44gOcMs/J3s3TbN12V8KSpAcZLcQXuqPB08L/nl9BAfdXlsO3qfHSIoeq
Gfu3je3ZHEDKV0MNb+O1TqZTNWzHDg5mtJ0THcAZixtV4oWtTc9O87WSxvbcGhqlM13CyQh2S41Z
IxZw4Lb1O9gnIxnuYlpQLlZvqe+53II6kCpxDthdV8zXzecUtkxNpPTAR3sqHmgkrsIEoOFUqtx1
1C+C+/xyl849vJYvc4hPGeJ2CC2j2dxWNDrTn9eKY8Sxl7WV9qbYtqNRBf1pDjRXhAc4RJEn2RTi
AK3KaHlSSv+Dda6nr4AxcDOhn+B+47zbkZZWyxxX1gOcer/sx3VTd0ABmlxjlGlA8YVD+vx1uDVt
Dl9x9R+kku3ALGywOY7c1a36MPBsOuSI+lxwV7UWmweO1+SZ+KjbEJ5KA7XvBUQWfbdbh6+0806f
dPK6LMFeFfJTYhBpQw+fpUeEtqT71CiVZAnMoXXgKhVIkWYsRgbj3PyWY9xJMUSrsYcxRnFozG6q
snmwqscmktpEZlamdAlKJi1Zg+56Y1GHyu7n/2efb4NBJBC5rqvS9DaYu7rBPh2gcf6B+NKdjMKg
oVkDrjcoae8ZsQlohGiw2wRkkQp72pYhxZ3urE9kRWyK4l51vj7EHTB1yVMjWKG1ewX3VZYCccSI
qTSSIQJEjEM+Ffs+o7/sl8LkA07/ZgxGOXg8+9H6FGQi82FGeEizJVfQb1Fw2IfovBMqlYXPeRuM
nBOK+KNYGxsHo/RVSg3AfStA+HAB3JLpLiUZlm8Ud1iWH74+WAhJxse29AuDxr8zmi42FkhaVKm1
J+3CbjoGB/ruQQkw7AUOR1yaZEW5ZZEBau/mTqeGMNW5oDOwZAWhFk6hHJT57Ie64Uwn9rNgwvDz
uuM+I3rS5401qPzi0IUF89C51Dn5ryDHl/0I4+gkwRmYg7hiQ21jRP+wM4pDTmf+88vtDIGeGpBt
yBZJk+JsLVkNkmkI2vFAI1oh5glIT0/tuYRH7QKpdiFV0yFWoe7+QHu/zpp5gPioiRbPWm+NDx30
M3ew3BbUL+pkGdq45TZIzqDiomtW+KPXvB4dzQQ4SnDHQtdv/2xlTdiTIemnGXKK4CCKuHDjRlTG
Mq4up0o70wyY/+EDbWpVNh7MA6v2xmeGGZeqLEhBn+4IYF+h4Alq5jbENC6JnB5acsOtr/zeoSjf
ev7aLKEK/W7sEqqJBidD5KzwC+3jn45QYUvloFy0IMD/Ht0ROKe6Mp4+OyCYaP65un7aSjgJzO/J
4/TD0SJHm05Ol5N+57aLICl3HmuYngtA+O3hR7GnVpTHL8UINhD5R9keVUdzQkOPLpRD2I2E7cTi
TnOCz1LV4nd6Kj0LHxiXTKGQRmQtQXWmdeTlkqYJkMZGgji/TLlBwtLlObPFREoNzFPIGSl7zVQ1
/EadgpScXaaef6MUDRLfRPdih7wVARqzvy3/tMagL8A3vwWKLeQ9x+oV9IGuopfmz1XAV45e8fbZ
OJ/tvpzKskuX0RPmu/Yd3vojoXVW1tr8lWze2eLV6fQKVgcXBL9frdA+zv/xtOyidPwll6IU1utr
vP1XnmN3D41e5IYk9w3j84U9nIiFyYhdSoImmGx7wwThHxPsMmvW7y5WoWGrPf5TtcD4npuwHm4W
6W5d4V7FLN1cMNuaMyaExP+n18gBM2dGy+C0hbJD7dKfu1xgPjrNrfH7x6KMaeRDSAmH4blMp0st
4l2ok3QejOk6F+KLwc52UAJ5hVMtKlMI781hj1pq13MY92xzN0vyOo2hOXGSmkqHe4aiG+PdaS3R
aa9VONgdJS4XrtG9Awj1oK+KkDwIezsYNvRL73qZxE9tOlnWS7baA3W26Z7rMac5nFfmvpacYhdU
mvYZrmz9tCLNgXUMwI8u2il84Z1v/pab6hoIqCH11EBILveHpp27T07x2FK/GVGCQzyygMTQJMFP
eoZp7lyyuoXsav1kBY/e7Ee50110kn7mWEU5bGkIAofzh550GY4lav2DAoCtNYfIo8DVjBvhJ1Tr
SBkrQENWawjiTotK9oTTjzqSHVZy4P+N9EAnxU9g+I39okt4mDlEXamdhLBXwIYlvryEZGMji2nn
2K56ARH8j4eV4ngyTzlJWWy9gFB/pFvNf9bVYdMuOIgvmN2yKU5dBymEmz+pVmPKiL79qtH9ybfJ
UO7/nW7VF44uD1vE2Hc2yswQzWE05UQCfKeSzavAN4EjHxr7anMs5Avl/5ECIUi2N/HdbT5lCgmP
vlTcVDJDQC4ldZUa+LK8Eh0VZ+VQ7Q/7KOycuH+2yQZRXvGycc2edP1Yku7HTy2Zcs9x2CNCIuJa
BLLPO2aN19D3aNlz9h6ea+bd6YymHQ9Yfh4RDDJ9iMLwbEZzCDsUBKDlofz25Nk/XfyMHLV4eE7D
7sJp4q5Y0K6a/9SpGWpug1HgzzUu+1Y3es3K4r8Lrryv/Wh36hYmtvYqXmGawgO0geLzUduWzD5Q
cHRc5ws1jbAuZbYUzV+1i2iuEW8GInnBrK6wyMKr8f2ZIPgJ2H5jNyPjzn9CnIMBkxIuJxmPdB4y
XRDwqWmP4pzW+mWmA4RWF9ArMcX3tmhxXv4nv3Uf6Jtr4OZLUK0sfT5SzOkxLUnIEvQ541ZAh6fl
8Z13+3lFA6najYKEJbCWv8+BhnJpsdqFebeVavXATcGZ1x90REd2XoANjozRxGORs//cA9JogFQk
ZNK9/Ay3OkocBD0RdbF8HdQMehEpV6G6qyxPWqUv8VWucp3CpP8XQGYdXF9hD0xbnhzpsRO5/CK3
+/w0Dr94UskWKnf8FUXvm+ZboJUdx4yMeQ37l6x3QuWzxqB+ztX2XISea+CIf1qDtnxdEppQerzU
fvTjqWz+rskB/kfkERW2dquFHxQSZSSWVGfp9kA1cp2M6+42f9Zv3xghS27bWPoxmQn7YeT9Nl8c
u7SCTvSzaNR7rO8028kV6Fh11eBRUT7gI2NlUMaJiHpYIgVyzPfi3betBZe2qXtFixRyCcu3emjR
7cOR5etp1FbJu2FnLyP7K4WtUAUptWSenstBccKRnHi5CObogSA43WgitGezdRFfP2GIL5bj+vm2
PDVsKKCZKPs53SwRLAWNqTKNESmsoCIWmtMJhXkPji3rsrWk4BeIC454i23x0GYBHF/76EOl9zsG
UTKBTSSDfE8nZ/w//H+naEH6We0nWX/zHn9bOWqxcDePVk8NXz00iTmxT5BDmt+OlC1xQeTBmJYU
OYjmwaS5uaS5Xy2/aBjgls/uDtCCMyfbGf8tXp3HUvaWktgGLCklODv/g0t1pODQAYMdjpSB28Hf
eZPBhBd6PCd/ePAUK2tEdKwQ9BzMmc0lbvQ4ZrKClvYgmeGqbHVWSnW57+b2vXbO+P2nrEAgZaSR
/6sjY35r3xv+vIea3komxWoTRGx2mAvDhSvjWqmxxeeI5WoqH+qV+xAtQ4/QSq8xXL4FxHOfsXfp
9twDiKyiffgPLDbY6Mijtzbmu94OyoeGxbkI6VpmG3YpNImAk1APRUa8Mttx8hZlLE/5okrJLNic
seK5dukkdlDMrjzZpXnAwaq8IElk213rOrPt3NedItPDtrWeBWv3y7JQI3qzW3meg7OpEAmCF39E
7jAlqqL5CIIx0eqHjywM2Cxia92744ng1/lEdrjqwWhhSxHxhXynxIYKmBkBZKIs7HpRUjwAlLqG
TEEvi3O+UIIdeWvfODqFU1Zm5pZM7GWz5sw08ty7UByI6kqbRZ45oHFwq4BhYYUXNHkxcM6B8iJB
QXZcdN0ipZBLAedsgdteB5yVYJP0oV1K0tvlh+m5WlCWNMQWHCbQ8M6LzmJ/Is8bK4rKNsFOcgOX
gVupkVgu3fY93smnqotFQarV+DlYdGYSZaOBe60+LYQMs7psOyjqNu3nKpxObDK3HxWD/5rg2isQ
Hjzv0YG45getu3ZvJp015FNcXdC6AaLqRoNN+a98pau+xMhl4XYw0ikgXoZgxXbvdZnfwg9FvZ1R
vNNvTiaQVAlMBmvj09zFetabe5wfQu5vLh5mBU7uxTxZ2ePfnrq3cbilNw289V3cldG9GpiUPgmc
ftGKm5ZI8HKnAI3wa8ywZontNjTbmT5pHhfTcSSAT3H3s+5l/+JVmMCrinea3KX2N4PYzcTAwBeU
SOQtFAnK+qNh/B/4jzY42I7LP+/xq1H5MAi1f+O/QPgBWpMqXcNU6wtgU4s0amjEcSsNEi0rclmz
VQqkR7H8WQkiL7Q3A4La85QoaVcj70xpMT7ceXuLXPUO8gWx0q/w6Lcm1MArMs8iMdo5ZUmCDZlb
tkQeLPnNeHDL8b2UeA97+CV/hDt1+yd47qFneMRSAQPozXnw/IQ1nky0hkunBUuPrCL84Sgx6tQR
bpahGSRsk13qPW/3aZRWIJFMuoVYsOePQqovJzzqflqwk9OCMqKqlzIWo31vAu6KkQuM2+wrlP4U
WmRPHfJaHmOeewvk0BfvTiYYxjiUPP5yWgkES2OT14UlIw/ig/BiPa/JOVKb5ubjclcAGychB84A
/e+o1Pi5oDDVQuT9p4D7FYjRR2zXc0qVGd+tmgGlZXF2Qem6gzE7RToA8RWjsiXWcFvqaVJc2dWz
//agwcdTluAu4dkCwhlG2LAYrVZh+FwtKQVTgAzik2xSF46bBaq0IwdvhA1PrV4sCN85qNei30gn
MpMSkj8nKQrLSMcArXWL40qcrRULycrg54i6B+shlIJtcWX/GK++35ea7k+GWlj2r2McrHgfJHmJ
u+1CSNs1ddsCToS31/W9wRySxfUPGbdAbN5+Q8rC7gP/6FXO1daZByOwmbWbUsbPq5pTCAFDF1tn
aNlC4ZxHx+Hn5YA8QuIxrdaf5lBTu7n3eocX5ACmlMBNwgsJxsd+Uh8hl69GxmB1+C+0DwWsnWvB
1w585sYVGDAR6DMtdCgfQi5LCg4scNbRhERngAe6begnxM25278jenwxaJpdiy8Ei/RPMGti0cuB
aM1w4r+uD1VrCK0DAdINdBuZxuyPRu8OtVLMg5IWS0tptD7NetF6D+ZPk9DebJ/444XDrQlT6wLM
5XnBME6Xc52qEeCFs+hoTBnfCO8smwZ65tMH2YThnI1QYMBILPizN+5+vFI3nu5t11Wn9t3tJhqI
9NZMqXBH+xO5cPpEHhTqUnICcQuxtoLyAkJOery8zZWTMXK2hAWQNvsK/W7p/bvwYe0Ax9TAD9HA
nexbd69F7DiDB4LhjsmBRV6YRyTHdIGjeuHEh+kMAZ6YecMj44YrNnkj4syfH61ea3FmII3FA7ag
EgICRe+0FbmFIYTQVxkQLuwINuIGCZyQjs8tKgnkH+Mtu26dK9Agsto6Z2m0gSvXFEWRJJn1h935
QAyMCWVXj+UMvmGPWH5yCz9DvcAXZ2oi0w9p8q94hrvryjAWXDl9yyFa6GNqDqi9jwuvYclEhHX3
MCi2EpZxNu5Azde/DrWFFz26VGERbn11W2p/UkfgE67G/DXWUTZwpruvsHHS5t0/OyfDLBqFyGis
Iu6GqculT7B+85KZ1B+sV4pBJ6le76bM69MRlefnfeBuAt0fmvSXuzd6hZKiQb5WXlrKPN/P3ySA
enaiotHnhFl3tn70gm8YoN8b/PZaX6GThx1Wt/lXH47nTC0IDZGWJ74lQSCXf9KXTNvNTvNUGIS8
NJgopMUy57qRdWXiMSUpMxd+p5/SMqIlp3QdAxI8i1eJWEFQuPBw03qTjGkNBHDY0bNWYcE5tDY4
1ai2k06p5Ac48PN4wRxb9rjStjNOcV2oZEPexVvNgjnG69BegWTUHt8Y1ENHwqs1rJb1+KiNFhNw
Y6yQu5973kAW7cEpALpWl7z9zOnVLA6Yb85UIpmgL747vMZjY/pRwLcEStjwkL5mg1m5n6q8GdRm
gfo6O2g9Kb3UBQkd1NNpfNmyxDaTDKgiXDxtJIz97/PYB6weUfDRsQ+gALt28ogvvzuIwCU0DaBy
4DRnMBls35FxaKvIOm9JHFnM/UP3PGzJFdwwxqr+RpcS2EqjYe2Tr13dy75ITTvQyD2reS+fzfNY
GbBoItp4J5q1/fLSbCNL2Hi4DZ5eUskFdx5ZIcSdC5tWBWrNJkwayCjJl2MM83z3k6bQDMhcRUI4
jlJQy71lGf7OfAEY74HqP6WyuEhsbeLFMOgCi3eqGyGVFRL79Aab1s6l0MZ5G/OSP7QuqnHlEkmT
2CawdelVXIOK/2stOWZzsiJS2g0ZwFsOlXlkeE5GPyUi45cf/vt24AHMmv0ex48J5OhNNBfEDpxV
bKBduZ3juWNPo3HB18LezoSCwP1e+jmqAE+HHkcP9DP1W1l1Hak5jNVyoC8na7AZHbxsOkxnfM3w
BmzxfoiD612yXyJe+TfMsIW1FPRZqhlHCZvvTknTdGLje6t+rjACnavOqLZohYF6SzKIe7H48Q41
NaEpnrnvo+pihw9irplQgi6KndAesLdkVi+w0LqLCGgKTYwn4DmKFvE4e045U/em+iNAaCbrSZp4
8+UgFkTvBRcenMalIqd1M+l5vfjovK54mDqpJOyZ8dCx7ISGrwEhNrzt5MkHkTnEQxZW10SY4OWk
gLp7630O21aNE2zOfXYByLvw88AtF35xrKluyeJJX5+r5P/PLDCRdzmY4JIQ3PCDljCHjI+4H/Mu
2ejgE+XY+50yv84L+dv9U1lFOonMcf5ybI+LOPdExVkORwpoeeyZadoI4WGKisaoUPGJaTDNbt/Y
Nbvi7aiJprXpsL8fGonDPjaOeNXsiTL20FTadYHWVmxK6bhnKzOUJPUN7hhCKqqb9VCKzOrY9L3A
AIJJHuxNq7lpqRpT1WNf1CnaqlzO+jMETVJaWclX/4pVJKzIjE4IbZL1dQRUW7kDh8wDlZjjTKzq
BJpwdWfP7Pcamp/0tQ04L6HihlKxjF6WZxu7KodpJH8w8IHzJxQ3Vn48mFOZp/1xPBSs8pgWSK6u
UM+/e4dneomuJnzoIQ7wol7pseG2LTGbqTb9hZeB+4wHi8Ya0MqfsOTQavrQSvy7+aDUtBjpoUEb
nXr3bCdcoa6k+bjRwlBgDTPxNDd6I+p9OBQTKJ9EBdPG3NBTuWTSB5rw8He5xKqPNheyruEC1T3U
KNz/kq+7w8y/NfkrAJ3EbQZZL0Uw/L54hOsxA6gzm45xPFKcUBMvi2hM5vkQ2O59m7IUi8Kde0t3
Fz9sZMrKZIMgzA3yfxuMQjetfBKdxTGLKRkUJvdyOn+vOEBlii+1LHQyNZ7Y0FqR8WTsDFb3fzDp
Sj2eV7hqi0qaq3g3WorZzu0WxirJWLaN+/fH30zm+hlUJN78x0LaeTl1u31+ivgX3ZxB8J/H22SW
AgIlCyMEtCofXZkgmLgVABsa4gkpZ+Z6++19RHvQ7CkhPB2LKYIwPpbPGqj5afQ3joZgsC3rcK6+
wQc/jRPyt8PFuJoct8LtTS+6/klraxiwY5SSj+DMC1HMHKmxtYfmoKdIlXI2MPUoOy5Xijk9rvyb
GUrDtDNu2IO6NYBOCo7GIn9h+l1GUQQHugHVW7m9fF77XMw0Vq2++UZieptG3d2iXnm33610/z5A
dPiY+p8xbB4iUlSGdItPNbTw0vtPewk18WUlXhYcUPO+h7e/QlAZaVRoHx1+tctbCUwJPal41Q8g
aM83Nr1ZsZnZMwk8K1o4FhCOHhkaXEiSaWNHJ2EcsOz1guv236Vi0iSTCKGvZTEv101C4Gxr5tpK
5bq3AmCujbmVeFs1v2MPKea9hbYEbojgUqOTIETnxr+s5X2sNbXF08R6D/NYbUMfCrgWKC7UqZRa
jnygRsqf0nVrufJKJvY/qrivLvnkUGV7B4TJYbGnptG8wa1aPgSAQV7OYj1chjlh8Ny1VxNOeqU3
y9Kj/Y3DCTSi1DX2hPS1g1nDsg8wyt3Rce28c7Hm+Ja/5Mv6CazjxNXFfl/zyXV3uDgtVcoBWMHa
87atQNa0OeeDin/ucIZlDl+AAOOhV0EtxsQ8Pa7N6zfZvrEokZahc2GEsQOsFXRoW2VFpxEGoKsT
0WQdxi3HfFbmhe6SIg6u8DGqx7fhG6kB70vPdX1CeaHWXS73Ji0bthnKg9eSMxoOeI9iQd9aTg86
8530MkWkI+ODZqPfDfyDNJhsDZUoKe72cNtXflm/WS0GabUUY+NCRpPhaaOpGK5hphP8W1uOoI3o
cB4FOgG8yeswUkb7zsmTLc8KyG8+T0dqqvI0+v727kapIHFWrAGNSFjhf5NaxyRd0xMG6cfzVLbp
wIrRUD8gkiEddG6iWOVnketIdARkzR9hlFlDoeYQamCZWg2mMMQ4DXCKG0Ho4/ohAEkW0RhEq/4p
HPZYD63bHKV/U8MLPwOVSKg+sotel1V/oBQuWsANXFaL1KCKqcXXSCPaZ45lFjuGpDlHyoH0HRZj
BBWHVVROcF4LkysUrTbfnFMJFHbIhD4Mu2WCOKxPYmy1EvA8F04iNISnBwyXuhI1xrdBMTqf6gh2
RPI20jSbfZ+PvlQkzGnk5UbUwoGsAs2LXvvST8I5+wNnUDSctnykrjPR3xScpMdFlwEXS9nDMQK4
F0NqzvH745h78wgKEMwQXHShwc6nubOzynnkYIdH5mt1cWBHHfY/1xp6F5whhbSOfnz0s1jW2a5S
wrcLxzvcCGb0t6JmG4xv+elEjbFfo57UYa0BIn71A+8buL5G7prPqSBKhDNF4M1WRsPMdzyMZgXl
An2GlmkW3J73bfTQaZnHvgSbDyVH7du6G6MoS1nCKACxu8Dj+xsQ0zHMM9EBZSxwUsL28zIKOUw8
uKKbfJkIbDZoQ/0GywdF/KkLeyyWeataRs6Yh1XPypcgWU+OeKwK+efiO20MF+rsGvt8c11mX0ll
4mUql+rq2ycg/c+UspDN+TMRKIEs3dh0/o32m2xmEn4cPUvsa4JslMQGiubVFJEBpO8cvUd9/cwK
TG77khemOZSUan2caHOvQxm7ldmTo/FSkXGCO6QHvXWYF9I1WldSZGeKPwIrZuMhk9JnYuYup1uT
uZxHrKzio9KUCdlfJfgjAQEO8AnjjH0HMH8eVY0YPeojlneYNC0QfSRP8ccEwB6SuxPG50SUCPN/
rk1rXwpjG+vlaNKTe8Srh4qkexjsfXPv8REu69JN1pcmT8+SX6XGNw7lTuE4Dfj1TWeo6H/ioJ3i
fLQOA342sv3gAR3pvf8Fhtqhlhz6TBpOkBNhtcecilZVWaAK90IhM+EQDALNtDzaXyVIurL2+sqc
Gjc5eqxpi2FLyMcKKnq8IPaJM6ZEM+k6bxM/u3IaYyJBsliPQ/OLvQ3xD+oLqcfN+Nq/AFQYmRGl
Y2w+Z+zbpH/w/G/Kz0iXPu9osPW1ENKXwk3Bk8AhhwScW0tj+44npxVW2mE02wCoOiBmdcxw7KUx
gnXbi75XnJh2BkKL1CeHHEecpKg1D6USxd4Z6iwJ3uieNK8adma/DcXsBCGRmt5sOuJL8tQYY7AX
x4vCd2oacmyrjBfP2Fk35y1+X6LNT7GaTs2DzW42XMZ9ZJs0CBlC5Bxo71EdjHkOuzrtUKSZ09mo
tsWOVU5jdgr+/ro8lg3CYI8F30VuapGzLtrmJIdQUr4tu3JCUcUeH9v3PcVqFDqQ7Rz8HOy3flao
v7uTYx3PiiDn3mw86YXlJvLntRDVDeHveX9JPFzTtmAMYHBt/MB+R8fzI1KMUogKyf0CKvpYu5Wn
0crM3RO5XXGKXswUVQaLrS6NW1QKuPfotAncvLyndyrnJ2gnXNrNAXSZv33Bq2mOH/7s30L39XWj
OcBZOYz0PXT45fLOqjUqR5Ut8KxmCGYqXHoEqy6rnWubfp5X75eyrdyxC8xo7ADeOYKuRhouk4dr
8hPA7GzrFEKZFC8vSFYyWrq9NhaW0bcrSDtJPLrxt9QEaZBgu8Ec+qSHLJBkwEgjADoOr7qVSGry
VSf0CoP11jaFIzeNwkQT8wjWrsQrM2Ssy1+HEYnRuU4fHmtw//PHjNYd+QiUVbtXW6NvYC7Z7lWr
5rsrZ0P15CYQBJPFkOvAORqbqo7kttVlVZFSUtF2a4sxukT0e0iWK62QIsWmgSCNVjY+YvTn0aDX
tSFbuqdTjv+xdiaAiRZVDr/7mMAkwmG+L0lZk1hAeo7K4NcPHSr21tyvU54NksJ5G7i1rSxkhv8x
DMeOL+LvDL5JHltP0GzPyVPyDr6cYqaGcs9NzjR4zYcqt24qYHwipb5wwXwTFyMfKwZ4TEvsBlAQ
RTQbrYpwhW2pfszDagq5aOaAxAhmuF73yOzAMJXIEeHQeRLlrcImGYStoTwTwzvSzjFch8JZKl1O
vn5q2A6AyF6/v7s2bAP0jZ0ySwcSS/zkWY/CxTjNuYrn3ekFQSPQUyOjgckB11dF5tZVCDuzxFgD
/uBtnIKdvWC/Xql40qWxVkl22gPVJ2mB3x7k7s18azW87NqRpICeGesw9SnEW+qeAE2/lp77NbfJ
6+wBvyH7n8hN/OtIzEkPKcJJV5F7IZtfP17oF8ZlcEg13O/YE6eAGIvsTRozhi1lEkd1l9uie1b4
r+xyLaxCqGJM0JZjn017hODbwKKZiJadA+ABwWnDlmcf4yVYitIIbWJ61ATFDvIFBbyX52gUCUm+
+xkttD/Q/I7XbWOY9TaR9hdkWDugCGCiDB7zBnziDjyBfYP9MH2NYwkEdAu013xwgh15BoEFbUy+
6OQldOKheyFoH7/XBIAdgOtDntBv7L+6Yvi9c/MKDtFez7Ziy7pXY9nAVelGal93DoDFQEcVm45O
wDcKqlRqXDkAVsIMPvzGsRsK9JOEJfMHjJME6VXSKoDKT31ZbsvsyKAhkGtpBANrimgvu32hbRNN
1Tjb0Ss6c41c4SOqFQpCssr3u5zPhedR3PWDPtjILNyBYD1PX/nzuIKBaH4RV7rOI5k+1lreaZ1d
dbtw3IdhN1v8p4qFCgkdq41ajXk2EaJ26ST3Mi64s5Sl0w4x9SBD3Gv+iY0t06T0zTpl1LhLv1y/
QsU8PdVW0z8Ku5SWRoakVLkUdnFYw4JvBy3V81poJuVEotewppd4s/hqq9d3YD+zgvuHpOHd1Kxs
YLEjeHO8E4zJczq/F7ZJypR66Vdv19Ayv1JqP6skh4K/UcwNM2LYtEiFWLhiExuvvCc9m3bQlovV
7RvPnG0udZtxZ7qhZG4R9D8EySS2XufQNYLnbcjbkzMAk+WZTzdM/p5dVF0acQgjDU2oOx8+FCxQ
Q2cmP9aipF2CrB/B99Jii8gF6qyYKTrRIhV19TwC2NeZzZrt3cWJc5Kqe1yc55kAMBpGEAotHOZx
dl2xqSkTdmXg7c/74wpAwqEPmt/wjZr+7BAAL5B0s5T+ZwsJv8Obg4fcAED78RYxn1+cPd3P0WfY
iFkakpPNQhy6+x1EXaDnZ8RaG2ktXhwutP1DG3av2wKbHGKE3yvLktbPeP2H5tvxyk90NK/Ba+LZ
XQJnCyFaemOY/7VMpWXugvLLTjx2MkusRwZsuVQHktqCybwYu05IwCAp2mQt1hqRiYs56MemfND8
D5zYG1mWfQKWdUvagWR6R540+weUMDertZlH7KS15UHgNjJoIAkaoReEtmbpkjv8+kyTzSx4M7WY
Pnr0zLAwGnoxi8cmDO4UD+MWDXz2zkDOnRoVapDBTpgvJB21Y+gzWzeKdLnWdCtPkxpX4c+Q02Rp
83lAx7cQNZXX2chmjUomOq/ErjHkeuW6H9kwcjXVyczFCaqX0FGgJ29OhPExlVynOmqehYLSw5Cs
HsAqxu/aeBuVSuQekHAaifc2uWO5j3stKSWO0X9bvcun8RlyH5msLnmC2jcf1RWmdF71qDU4W0WC
twR0UyhbEcpqJRfaILxHiGlZq3Zwa+2TotU8esbJPVb2ZvSdVHuBVuVhlX9wCoAnATOJ4aKVlMTy
6qm8xeWBX3/sFrWZPs+8hLSdr8PtUTFZX4P8z7eLP+0lE9qOhcVjoZVo+coVpAiyOUVb5Sw6ZfCW
h28p+qlsQFAYhN9ewpb1WHEJv0erjIARUq7Aba3uvqnZY8LHWN27qXyojp08l3rjDhS0WYp2VXft
bz1tVT9ySn1hrnQMgry1YhtGwlfASKFRw+aDm1R3cldtwNVDLwCCaCDDTqRWV8cyAGsRmSsNLx1W
2qSnru5IcISAu+LWstsdMXiQuL8jou1b11Ycal7LauVdWg9v0MSKnf8ViH896+CMV+HrW2chU+iZ
GjvrVa7YqH/BfWGeI1VpZ3MsSzXaOVmwt3dvqaw5FyHX4+KB/KswIjVnPyDjj5nkKgvYs0buA+cp
4PuCXKcRTfd1g6xzcwVh8Sbr3U6DpQ2UC8qbvieOOvlTC8RnDQ4gKzwwZ3lEiXb5HKWYFhkvhHkW
wKUsH+NCzd+0ddtWICz+8Mo35/P4pb+Z16yAzwGNNgW55eUk9AGvv/aOOMJnqLS+IyOnk2QTexw8
9tp5j3/xSHRLPuq+pzTY7696X3z2YDCZkx90aLAmzgl+09BqXfnLPvx5/m+NyJTJrHRxFsMNC8wl
/2T4cY9n67Zb+qP/4i7Az7VB2uJXpUiaN0ZoBY32eVZiPOZqorfo+A7fQSD8XrkGsKphr/lc/Ims
1T+D6jVk5LTy+1gz7LUXS4ga2xLO+Pg38HSlVhfWLH6SyytfMvEp2PIab7igl9QEG88G8Ug4J2UN
3vf+ZYraEkaj8MFOIpd050HSxIN4rnMKPUJ3/ZrtMlRoJVpr/TlSh+8TApdp0WbYqdRqQXDq7cvS
N0rVK5WKxkBeA1ltd71qH9wAFLXQuZWJGesihGnLClQUwSff2TGCHgKTuGgt+C+u7tWksmVqbrpc
eSZNc41Mw05JkoQPrvCA/720z8zxUIkEmWsgzO6LVrCFY5AB58T9Om6svyHtOdzWUEyuNmNHMATa
7Qe431cff2lQ80iZULP+CZwIEVgyB9csd4P4O8i91pH8Khs3ZCXZwW47foaoH9nzjKCFgoQYm/0h
ezk4PylBenhZAT6JzhAUOp40qo0dBXcPDpeztAJJPphr9b/8p0I+q9BzuRS8MsFTSDJ5XeyS8nuf
BO/F+8RxQOFOhzK9A8OE18/vbLPxbQm51o/VyHw++TM+jXb8Gl2ecU0VLxXrEZQQK3Z6I6kxo/2H
ClIK/qUNEUQHLdlpkMnpdbmxtxc4paWrliFro9gO92SkD9vdKdZVLgZSU+hWaSusD9ZNHY4WUy4z
y1Liqf1owFOMLALofn8CX8gGsXRMMt65NMd+ZgsKNZHrlZ4mcigf1B5otlX1FOcj+nh/+jrvACR0
J7Anqincj9ctYQmTcty2x+l6yP4oeMUBEAcV8axIxAd5poVhtQzuO30wgebR5aY/DWPIjq8tvqBB
lZxVZky+UOnczFjNHF9m+L7WDT2hzmlAecUNNVYafQmnlkS8i4dWMMNY7IlX2HAK0fQwziRFL1db
+K2RAJFdEseocfZp/d9tXVcDstDafY0X4lII+dzlfl02lTJI3Y3WDIuyW4UNYDY74QNzKLT2NjRv
3EeGXikYdFUWJvKo3myWD5Q1TYrsYDhiDnmj7QG8qBeXzuYAnUcK0Lsa2w9OLNAEcgTHTmsQxJLu
QAP9n7B5Ml+dt9Zxtw2h6xJWLiss9zhIMNKMOy38SPzAxong+NDDf3esL5kNkCwkRf6gTeNCv8KK
LWExSueMaTwBszINy3WZ5hoop3f9JR9zzup0sH4vSaGUkAXrqYHy/UTKFJXnCSc8Vi6rcNSz28/h
Fe0gqpI+mnH5K36BM7nOkDnGkzg3JHEuXZglv1BpOwqrGA9mTnd3LavNM498HYYphY1unCEn6Mkx
jRA680ZRHRejhObK4KsCgf7ZHmACCWVWapj236b/kqpRUtaYvyn/l7YIlqssW2qG46fmudXAHM5o
RKet6v/Rpx09bVKeH2icII09wguQ32ibYyIl2QIvQr06T2WQR8K2SbhDCeRtY96daqGZE0bW0qo3
wowNox+a1TvP6eyzRITgqrsKDHz6Ms/qDiGHT/0O7loBaJd8k61dl1k6ie72lDMvVpq2v2NGB7YZ
4a6LJkFhbPCe0DNY7m8+eoF2HOBYjOHl8ASIUAqfr/ITSGR9FumJ36e20oONaDzsb3Pc0/iqY6+w
qANUYBGbAZi1iIWrUkT0bk2r/owCj2Vs/1zhGJBREiK3LQ0Nf83h8qf2MRtq88ixGUbWeABkRW8n
w3Pl08K1GnV3G3TT/A4eOyUbaa4IUDLTVlHYIlPDrNVrwL6bZsSXCbFcMG/ugaTQbdUDbAm2G+Nn
W8aOUfZ5T8SVgcOj35vPQPQuOvbu++d1U4nz5nPpyTObAMQ4LAqUs6XyFHTfTijk60uc3haOvk0n
6VXlFQKPvmG1OdD5GEkBcHz26oXybXlUpfPH5P0W8DRTyQ8vtPlM1cXwsOCk0DOCO/YCe8nk/mbA
bzpnqxKj3DfjsuaZhPazVR1zd1gIToFiIOEwvT2GwWa2y+/gA0y4Vt15H237o8skVT7ZdH/iwhSC
haUCZ5qsJ3wSAJz/LMZCcZqhfALgYijsgHEHiH6sZh31vt0Sid9m5aGzr3JwHabNx2129Ty1MMSY
DeEWnB4waKFEtvQ+jUL7o86T2FPoWhaDRUz0xaHA1AQsEhi352tv/MLW2cANY7u6QRqm85CvOZC5
K+qlKwrjmeIuwjvRXGHxzK2q9FEVsnz0IfURRs+1vhSpzGEbfyUjnpJAo6bkBrIFJddkqQnuJRiL
E9JVjuzKVAZrSg2CpOLtMIfE3YFF8Le4WPMqLcyUcCpeUfOpk9BV4m7hfnJMcDUR+jt+baKJ+X70
582uW8jiLX++7ESNwq/icGTnViuiqGyUvRUa96LPn38CrV1UzzmGdjIyebz6JRLImvQjl66kBvaR
KHXUfpZLY1H1QYMXnziLUfh4dob5oDXIziV67kFqPS6JCjbcwiCn5S7cudU85W6LSu/Zh9BFl8UZ
4aaZ5/TxeO5L7AmrRCG181GuTgic6tGmRgBZLoR3jVJ0T27yfSa5ryCalIHkRMUlbk5O85I2VMxj
v0uoFdWu/VKCWYR6EYqEon92KQvuXEn648bM1/slso13OsTcmz6gxFjfMSoO639ZCSRyiOEJOIsQ
8o+EJRmqrUuhftq07ys3p0uK4LlJv92JGXOBjgy7Kp2KGfC/cUN13hbrzIYCtVbB0iL6Cjn6Qey+
veyQ6xLQVwKgwDvTomY9uxO4NTrnLVSVwopY3S2f0BrVbkR15t7FGYav9jvHREMKoyJeZitOhdmz
0MP3tyWu4a6pemdmQXt75n8bu1mmPQo0XpItklx/2kFn00B6tMWXLwviJmIkoU5pa50/I00Rgsn6
7wk7oEvIlqaVDzjoUKCsyC5kyiNTIVrr3Q7j2Jgk2yKw7tePOgZb5n2TmaO6DRHGViN5r9bYMeOQ
1Mw80Hs49XZjof9C0QfRTJtfQbi+NsfLp43ipdaP3M+LmNaaCNWCF06VTGPJA8/fULT82majFvAd
FgWyyImO0fEMky35EFa7usX1fLWVKTi5oDIZo7S6InYRn9n0wo3tAGMXFDZRHgiqRUV7hhO7oLMd
3vUF9MciyMBf7g41dwpocE76bCWad9AZHQ/QWKQZdk6Q7QsRycffw26TSRn+sUGi448DMuL7quns
Ihc5zzKy3u7lzcwQawXDG+KzQk7K2hnRFAL+fKVghArDIlQu+6y9LBk8lO/aOL+O4/F/pb0i/Plu
3K6aPepIBf/odi26bwjBUZ1LK0etieNvnGdJSH0aI+Bai/qNGMJsomBRmqnsqiA70hBWJ+BfSXxQ
fch9c/VdDlwvri6YAXn4CoowAGHEPwKNmlRXX3gcqLY4HplaXqBSL7ur6wauWdKGR0k9wfGtuhWQ
Jih+W7itByxoYRdQbInTG6piyJnwYZuza7LEYPaGgdiw5/n9JZkR3fdtndeOoyqizcA4ciwYtq2V
8fnz2HXL6r3n8NkZ0DLD3SC6hdlWlVtpB9SZXQaYgk4myH9okMGfUNobHMDqs/mlOyA7FOMhU/ps
apgppuGouq5J4LTVScbuMTO3z3xBykuhO91qkuf48fzxJJx6WhYm0Nvdq0GmM+Lk51UU2Xn0NfQx
FmgY6kdqkmgbHyr5yHbUYfSI7bNRQTigNEuDE+zgcQB7lz/1kgwqhL/I1D4VOLOgdeOf1X2NAxvq
09T5zOR5WshW+A0O68Y/rHovJHoqHAIKn0rzhlalci2ztv1bX2S4FgLK1Th0CjBbK934UM5WSyo/
zipG2BPTtjGbTbxI/9SE+/bGzLl6Sjhx3CkWwFKU35+SoWfj71FPUYf8aRjjoC8TllvEuKNgI4Ox
/W7cuYuyorS7RpaasZo1gkOB5ktulsiPape594aVZImzUe/ynVpJHP43IAopqPAYipSNZq0lM7MI
foFJGHCIu3RhHwhIlpwWl/ZR0pmPacxSoG/CkwVbu05I3nuEd1y5JFi34XvoHddUw/ScoYbxtA+w
0NRatcexPtR644xzOhenSOIsa89qlsDHSbJuaPloankLmdTOcdAovEf1A8rhinbvdyEafXES4pUT
HcYhmw26dKyZQxtrpHZFdy9cUF2nPzm0q6NoAhNmq5d46tA/PdLF0v20XAu6FvezM4dK7eWWR6yR
hbonFpfH/sSs7qk5rMF+kstKsN92Qqe+PiYyjcN52fC/fNSGOB2WhqYkF1f1NuezpSFS54wP8t0h
SedMwNy/olp0WbIPecfWEPlaatXuGacOpnJg2OmiaPiGCn/FBRhHxl5k0u8YS4yMcwMB6Bc/3CbM
I6KhcCLgXRE9C1oGTV2KrunMX8hNBaQMzaiL2n824q7wfDb9W/eibBq4jTP8AGhVb/KOKibdvVAa
Jw5fC3Z2cSbQD23/4NGk6uorLzwiQ4D+JamuPM8mXV/M2vSImDsVm77fDdHr7+scACbUlnWJsDVi
pYNH2pWIc2Ys0lGpGP8IJ3egROODX+cbDxcuEK0ATDKvGnqJbl8K/5MPUUcCa9MGEs9226wgCCML
mbi2NJcPpyU/+IFZWlvw2OkNRX6Jg/BpeRmwg5f3v2+vmeRBTGBb2+Xuh4b+EQgXtxrsEgxaIc5l
F+71ZbAHUYdEXKo/Uw3Gj1VyfNP7M2Z8Cv2RNPbG/a2ffeaBH9nhAzwR+xFm6EoklkV7khvk6iSa
wA7dr3XlW6dnlPodIZaSMKrvqRUieY36YIYKZztmDcxyO1DETOTaghQxfJP4V2wOtO1nlXQIDvLK
sBPEZ/HDjM0VU47XRgXplCZzFXeiW3UA1pd8pcEykbPPFNEWWCaYODT0zVOmKbzXET9ypjPl/tvZ
71LcVXiCa13xRt51eOSQmlGbnsLj9FYidK+5nYccWXvx6ekm5GvtdllTrISJI8d6IbfhMjKNqqge
wQUR/iuXh0POG0+kERZzl+36Oh2vEFOaXsGOHjci8iPNLxyRxeAx2d6rQ5MvGC+ofGRLFCUNxJaK
nXrMIa9fsiVadiV65ZwuYSfiZ/IYlyy20J5XB2P+PLYKY2Cp9lt1KQvPOTFV8Ul80TvnyosIF+Jq
+CFbeu6/OtyDKbgE+LNPLAcF7oKfBtoORw4qHatH82ANzym7d5IenCc+IFhQX/lwmd+Zbg7S8NJg
CCHRSHqx3b0GM0V3/oJQB3BHGS6CZhvOEu+Vq+64as3h7umDU4QcDWNjdOd9snY5hkQtIn9KyYs9
OAS3XNdCwIRWV7RIcpv0VB6jk0pEl/Pb70sZ4bZ1Cv5GzyVuvXyo/awNqisoM13m9IdtJICu7u43
5JmblVepWsShaC4FkqkAJrEbWOx7ehq024YN35udbrONO1YSMxBU1BKeAswaBgBi9kIXE4UBh8eh
MGniykphcrnjRTIv1aC6zc/Vel+dzxC3erCRjjEp09k67Vc8uggQ/YXXzS4ZhSnhIOLIhFB2Gcjb
M/aS2teSVq5WDdpjqn0+nIrGFQq85iZChwkz/3vLl2lKvLwqF73d/W5982bTf5oDtU5+i1o0CJzq
4yn7Wd8EvBLTtYKfp9dr8f/782V4Row54IgLhbDTGe8FuDNyoCGK0Bo2UIFHGY70LxDhPGkiS3f0
YwqHwt3b5vt+jrAO06zVILRwa+6rOJR+M1m+79b7K5RkFSSmZMNj94jFYvbSRM2vreKthtxKcrz+
OEK/6dLJixQrJ4ilBXfemg526SUC//CO1FjCTegkrNro2RvtwSgyMK+zrjgZ6o5VBz+A6hwd7uGU
5Agnx1D9mApXpJYs0yqMdAYNdFEeg24+CPFboGHH+7VL9BYnjRQdqC2lE3QgRaI0jUSm3mlXE/bK
zgcdnrJh+rQMlF36eIu9zVxDmXcAIFNmY3Xrj3b68FK9AUqvsY+XN9vmgL6gsxloJkog7d4HUky+
W4Kmsalaz7wO/ZYDF1NNSAAaDfv9gNyWNwNcuT65Ner/FLEZUAyA7iCP/ag9QWcUD1ZI4OS2FiB8
/fSquOrJBdWtCrQ6+0XG1CesdeDZS/5PlpvScIcenhoQVUEI8MntBpYaU44s1O0rJg/WKeJDFxr5
P7SYlUIMhT9YaATZbTdifbjvhULg0KeDyW1wPrFidEo1fxRwktyKRd4+kjE7LTl7Sl1WTPF9W8cF
90OacY+lN+8fCLUG5di4asEZ9XhgN252MYBsSVisiDck5796UfBh2NBfhXMCp3C20QFIuNAQIvPd
H4fPdYg0PopNK8Rlq2cXnN7EkPhYEdNBnJtL8d0jy9GveiOiXb38FT+E8H/4/VHTWzwYnd2q9as+
Ah5wVQVzsFxNUv2ikNBcpQ9cQi5DkxHI0xlMwuzX99z14zzzhVT5emZUUc5HfUvwVNv9I49+FieC
mdkriwjC501YpKcNgci+hVPovhEaBT/9xosk1xWFkXRePP4Z0KqTbsWDvSiocWJPcrufpyPCI2u1
IqBbSj9YwsSo//jlC4dEiPAn5RhNTPi+xcjqY+q41+zu+lUze3p1udzJRh7aEh5+iPxM38o/o2ph
rrzpD9uEoi1eshyTRYPPx8m0jdXWrOD2a1r/UhAjSGl97wwQ28feu9RRYOceL4+/dOarar1Jf11n
Nqs7+i8sZ5L5Rx6QgUl4LkJ+BSKNAf9+aG5b0AL6DyS0B4OMXRqauy4d7yUHjjyaj1F/sX6+cXEL
jeg/hQpKYrbrN3yw+HWHQ6/RYJbUEuhMlKS+XlvBMplGCP/ciz30uJlfqmZ+g5iOegPPtQVYJzgD
quLshS/ulwStBmdtQ0uY7zVNuBdx36EulUSW3p0mJUbnyoS0DskvkR+m4oL6b6z46UTL4T0QT/Qc
r421EB97vp+4Arf9aH7piQYt4NG+skzdctAbtU6oeMWOVZS+ittVQyt0usXr6OCnJFhKi560lN5T
Xfz4K+WH4KfLLyHh7tUoU5KwxhSi6/fOwRST728YGS+4kyGMKXT16RbzchCGqA2K4KRKfQlYImJ6
2rI5j+RxmuNa3DruoFgizGJp4P9SYdcMZITlLJ1WGKP2sW+XaZ45GaluGtE+Pqf5JlPlzX8ElFfC
dsHJvCl+bOWUorNuNN2WNkDFYtq1lhs00rmC5niKbkOZj5kv6fASo77NSLtZjMFs81vuugCP7EUj
GtKFBlGLlV9Rl9NtOhgnUSHNQbwBYgA4BiXiVbhbEEvxfa34PBf/c/8qIiEv8YD9zpWtcsGjgtvN
TK4cXFPlRjbgRRU11k9q/V8VWjf+kTj5ee5PIva728fBBSi1LA/2yRU8DkqC8RwlfzDZoyRn8BeW
yiA+RfgJ8d+Qu74hYXhpEYrEwp/JHAEdOoFbe7dZNGP3fsIGX7vEP76YxAmBdXb8JoJ3XUtPk0pq
8Yh3iHNJ5g1Kiz1E/YviJ3WUCkd09XT51aN8CTSLf67gKvy4ns1wM5qy3syYtk6nayivr++WWG/b
nC629Zy/lkftT+80HedHa4JGEPakMCy7emYPk0SkIGkbt8+o6XeyMMzKtbvVcbzTPydiOig55iKn
CvAyhA6tdB5JnYHVmU3ivAhK2HJh6kj+qDX+Hji9C11Q/PVS8E0X7EXGITWM+p4719XLF+mLXCwO
khqocYAFJt+VqetNNIoilhHw1VonGNBV3HEQy9i20+qfldPve/U5Y5H8UICVaC4izWPnFAlLK3E1
TSA5K/oP3SuP2F71r7Bncvm5jzxIYyxDBVOtx3s1oi24n9D7O7hibPdR3acdlmJWjZWGElmiR9+b
Lkc0wkbBegowAzqNRxaUqpPvX4oABJfoP4HRZJED7wknc49SeLW3TjQWIPzK0/JedMjxXkHGX1nH
I+4QumvOe3ree4+iSxx4XDvFILCCXbOvtAOfo5PjpILqCI5cmxjSuTraa8OKibQNR/VyRX2YYAQg
ZNGOr7cTP1sjASyLiRto947o+iciYin4znv1MaY07gzyGhXfSLcfvobf5D4CPXO9qhKrr8uba3n1
WhBBXmAaPCBLKYJGjPTfx+OeDXNOCbKGVRDz1O6aJf2kJBJrEkUpD3+Vo/8NuIV0bcL1ZS7DRl+X
Wk53JaO6+kBEp12xQ1QPkm4ILQyI+MCA7IfFv7yzeqgqaI5WnxLJ/P3ksPI9q6lYTxAM0kEXO8Bn
5xM0BAOi2OmAeDI2GwlfvJQWYMxpCJyYsjOn87ejCAXPenkhgsk7YOb00JTh4MPquKF7FE6wcDqI
pov8A2T1GE0rXDwc/rGvudjVWLgl/NRNS/xkPRFu3yjb2NAFilXozLRaUtG4otQFpkTDBl+n8VR4
ke3y6gM1RTcAmECaoUnDrirKc/s5iJreh9K5hfxLae+G3rBX7GU1xWOafbcLGlLOSp4OjPIbcR8n
DEP5niEPgI4OWKYMmUhczxhasgzkNusj0+GLcCWuNCuCYYDeyRcVkDwB6JBKH+fltVGOuifAeu/z
n5rZOP1KDuIO5zogvc3lVitPG5zy+5V0yrnodZKivxE2KoV55YOlS/23MkkEW5txALdWH0FhEW6T
wngLz6iUv1cdF9QH131CFkPFDuj9GNo0DYFjJKdALyf90QoPgDshDtxkD97Ta5GMQkYfJstD+28g
MVQPyKYMnoDm2Vf/qkPBTf2ykilM2uKU88zWVjj9tMo2abxNWp2mukKq/yfgUMqwS79D6ZOQbZ24
1q2AvCYyYjg4dNEMbd94rMyXhj6f38svUJy+8wSsizoh5Zfc9ze9eagHAzvi3jJXdkay5cY7Nf+h
4diOUkHe87JLuMJsTET0yrcDNG/zE4mxxru134SkiHmN6aGNwCza/304oG5uQTA7hpIC2byBZgTM
cXFLOm6BJm+7GN7Op7VnWtTmhZl79IPTgpyPdRrJeDVAXxnFvYKYJ5lsi4jTzqt7pi1BFwe9Gvyt
ijAnCh3p49InsFG4tLUVx8tcNIFv+Iw5uSaPlDUNyU2hoSyd55iTTbF+Hld0bgA81hKrPKqon/kR
jSV86gP+Fd3l1q6iSn3c5SgIpuDi+pxNt87lEXzbfcXpUf5bNaGvqYNMT4GBm1KbTAwUjdirff03
Mq8wpUdrW2y/Fg2Bxj3bXk+1IPPf+tD1nGePaMP7XRjXOwQB2Nj4/t43BLXzZcN4uAGnXPWVPmtu
afLvLGtSiYnLJIgqBygNYdCO3eM3BinWnzhH6FQv1LLQ5R8dWzXbAaEmbB1l0/0uN0fItOrhAbAo
LJEtDEB8qWvVRPTub4A0a7/SWDwRXkbdesiOlIolDZP/BRrF3ebERiuG3ZhtLskz/ZC+/8ooizXg
YlTIOm6INvFlXTeiWvTQMJcht8P/8V0XeUi6jOw0iU2v0xCVFXNNeuonVCpj/VsFe99uHF8IgkhS
cl6o+pAudxYaLyv0OEQ2kRsD7ehjp5pdIGGapE2Y5JFXFS3C1FpgRSghL7PoIkMDq4m7QsdoNg8L
S59eyZlHd7Rf8SUbhsvV9zkFVC42gUUhdKS5c3n+BY+iPYA51AiSbaUGr2Racrvsswo2OJaFQa3B
TDXx5UK32YMy6OL4d4JdYKvgGp2JNXvSI600LIshPdTati9ydkPOEZMfmmwlTjxmfICKMLdujG2K
Ey2XuY9jGoiA4ESUCUeQVf2I/cXMDSSCsrSLqe9e36WOveonTXWBjk1HVAg70LC/TUT1ulruQ8C6
D3DO6UNcPXiEoiZJjRACnJi7A+Zu9g9fKNrQsU6TIlziTDwzT2I6jRDbhQAguQbGbEaJSv+G8Omb
1+mq2ilcDoM2EJ2C2KaZck6V7pNt6h1TV5ptC7c8Z4Tw6E2Wv5P4ofs8dH5TW61vjON/ysiGVD1I
VmdyUh7kTKPk21iAy/ayGhh9JWYm/f+kcvBiN1bW+0QGNL3Tbb7TwPI/+VkXF9FJSGN03RY3KeE7
LaMdEIDfiE5UEbCjLZTzPzoh60S1gwZUXUh9ormd7K1D9ZJZJgmxdRx+JJ8Rgh4//pxTJO0NkUPf
1ErktCKVEm5xE6dEpoS0hrcEBcOA6dO2qSNqkM/LwoU2NXHoMBR7jz0sNSOXLDbtdgfCcY7EMclo
BgfRV4L4CI2yE9//hvF8QfhS403qlHe1Wz+4VszD8Djj8DYDpT+lig1Er7pTRYEPMu1oMlhvXpEU
3oDQXWFf3tQ4w/u87TAReqyH7jDYdHebgMNjBmhr2RsbXczVHIsBUKacLTWhuwU0gr8GTXCJx0qA
x91DsATHlHobA/dVrASKdSORiSiGMmYL0jpAqCLpS0gyycuZkn/ijt+wNidamtK2OPhYy3rosSAO
rZ7nph18xwoGFF9GzcFWN9s9lAJw9mlbhNsFclb/Yvk1//+zbdVmrQItbwGhRJWEqJtaSAgsxRdc
nk3CQ7X/ZzDSod82x3TgsfVB/Y1/NzFlVh1mblXJbzXu1MWxdO8/W3NDC0BKMasyIvSAHgiIJHUt
NVXHMZCnwwQRYp2jMi4qLZW+eXuYam52hKz8xfRWZB1j46gt/TlK7hgtdRCh70L1sTaeghQG7lG8
cPmjOxe3SUFOpNsJZTtGeI6xiQUMagUezc5QNo5NwGFHPlaBWZw3IidTdSDQJjjWZQjRIVQvM85n
wX75941HHNzPCThyVP3EIMoQ2+pPO1GQKuIqlM7tBBdLOZWSxGKOX57ZgCDrMCk9PVtaHBfvICF8
sjphyLSwTFouKW6/8kcMETWFLPytf7hLr1HaEyRiDeAoTIwXE1eJIW9DebHfcGiDRSAi2UHzrExx
LSqSiF7q8yZFOfF4zp01jRFvc94rYCJfZ14ERXIajrHlRv/mjJ4Vs3mTKnlgazYVNcrPrryXy/uU
MWd/ByraObRIzlhxivmeCRmW3ojBvIIDQPhC+JGd/605sAoMqX/3n1I3m56GwYHOhvZhekcTXel6
6LAgPFPGsOTWHyhGegorcs3dc0zEP0cQ7G97jBXfGG4OZyKGo9VPnJYPTt/1LNhC28bf/aQusFKL
nmjbUjxvJCKJUqPra+MTaw9vO14YH3rEvdH1PbRfym2GLlI0O0oEn9IArxjINfsKCxPnxuJdxWiM
tEObqys/d0y5qpGJs2LdSR4xXtYJ609yryGe3+iH90lrV9P+QqjMumbto/Wv2InDrtV40tBngQax
Myt4Pz+/2BH8DgaOyhopr58Ouws+q9EnYbcHNBYx/6Td8bzF6EZsjmCLC3kHyeor0Lukhp9dTOmw
C+jCyuJrzWNGpS4/AheCfaGtSCPUpIy+ABU8h55wPnFHqcrdne+clphe61EB3sQuq5eb07BpVN2G
/SYyPOOedbIyzedAbJA4M9Y5HaBPItCf5gzs9a1HEc9p4w1i8m8JW8Z9r+Tr1gCsuTdtBEByNzJI
VWmirapFuj7n/8EQL+l6qf35j4WV207QBGU+mtvr6KyLqezmoz5W/AxnOOUevenRIfdk7bk0B0ZI
Ny1h/duGffFpeSvGC2fmiNxNvktwomFTbPGMchruyBGnObncIX9pbvenkMgz1RsG5v2cTZ/KoCHl
bxnaEMoJWNwExNAaRS6exilFcigykgjaVoBrQVhahhSPlrxNREarOXvog40Y6pay4joi4BhLSHv6
BLD2VRFqw0+o78uZFiVmlOdrxz++oYAfDnW/0dnEbBKgxLMIIoQXKa+t5tAvh6tIRLscbidodVYc
vCDhagYNw0PWhTSnNXuexrcpl7M8Ih7lq3KEPlhWQENljh1fkhl5t3+kda2T6m7BfBZU8O5ySopX
K8sgFQVLTuJVt9RVsxnSLl9XBnTZS65WZyW/k9zk/VX7phgehmwQ0eDgX5gDI05VbIG4lOJ/JLf1
GtmmJ8biZeBmNa98BESOPHxbNRF/s/5c9br3dhxJpU+8yDx3XQEeFv09XM0WIPsqwuoqjT69+eiT
1awYAyaDeKCkkn3IfQy6C2SrVbrl3lURVYlbnJu4KMfKw4a5KPL3pVQbVNWahOpSSjYXoMuC4Vsu
KgPGNunnSCPVr+FcKs2csBhYKB3h8hIV47GF/RuCQgz+Q+Fv2u1AgUlWGZdf2/Jk/Nqa/nReSsTU
eQghaHikIXczgEu7dSstC85DNTSwvSA0GcXBMr8Lwq2j7hdw9iBYT5U7U9UJgvrlVEriVHiLAMe9
clwYPCtzZA/I7tXQdmEBZWbEXjARR+ojG4LlcdVAf6mZGtxaHvwywxGgEmnyI5eJJ82lIsZpSTp8
vEXqq01pW6Kc2SLMnQqCkNZDQnRuBhJmEKTW2x01/hYPGFPs4zUnZUI/x9ywq279vGQ8GYM9ZTZU
8Ij8elE1qXmTe68T7F2y7ZJoUHBVLUzQxy+fyizeYRF2sdSB+FMyYqt9/PxKANeI8RkEEuzV02yK
gnFp9iiPgoZ8E1D01oM5KTZkdg6Q1H2avTDtYUyLjPXrmOJXV9xUIzEMjoMhlHi3mU5c3cVUH9tF
2eoClO3xmLAu8f/ID2M0yW2aozN3wSeTaXCGPWFMrfR59XZSolX28kFVNbqAXOdSVBOom/Om3nLp
6Tnbky7+jd5PG57Fypuci/cgTVH0bS+PUKwIayi+vzjyahCFo5E8hqKQ7+sOd1tIgwyhIKGGVy1x
b5Sk16B7INy553bAWIDZBJacBHs+UKPOJidblmc6LHgHUlQBKYRXEZprg2Sc61rhvjiESSBhru40
VIs66vBB/Mgd5SLaO5kDRbYClChxhlYa4D+emte1z6OHvogBoGZPXeQ9h6nliiQWfD91Qn6aJO7S
fnl2uDy/iuT7/S3BL1uLVnbLcBlydJ0pBngen65XzoI/6trfepHmq4/PvFdY+kY1Lp3SWrR48loC
HJBfY9Vwg2vY6C0VHhr9HWFF+wePI4tMZ9PSLnLZcETFqkLt4RWe043l7bKLoV38m7p7Qgz3i68s
nkhA0wq+QmOm7u9PSkfllyiVcVDo5Q86pKwFtVgJ7vdbmF5OwUivL/h4BXtalNlORv0oOwcqjRcs
4rStVWZf/Gr0OgKEXCgFr90zYd7J7becYVtW8ll+jZOXYUh89HnxB82DUJYuqpYXZN/hBNQ9ff1l
FfYOfglEK+Fo6kJ+HfSRbvrBYZoYHCMV6LYP4Flm5A6OSgAZSfdCAc5jcrHXoTfhS/E8yNNbzIf/
P5oh8Fb3ml3T0W2PCVwa+E2E4/py+HStgv5vn1MuqPON6tyFw/M4YpbK7Km5+8ZYqRNfjgGNqhef
ilhFIitmBawv3vJ0fctpYHgdD2gNOmwMrKf4UY0x4fRlcvgaU6jb3vARmF/66XUdID3yEjwpw93p
6aKnCZ/NBkAoq7+6dqFQMpqlZpDWSOjk2dftzOBMT8z6pWrjl9ImyaXLlsXyDtGQXCaU6IHF713S
JVrt9Y+rYIyCkRXg0KYGL+qf8FsDMrvHpfrBZTGIKejqKHuVVKxBZaOPfe/9hUxs+7nYd2d+DHqU
RBEZmlqEWGRnEqnpSe9rIg/tNWtyZTlVUmLfTx/N57B4heVuC9r+UaWv1+HnPkJbZNJQdc3RUQfI
Py5TbVNdjQ9LL9CHq0z6GXwt3j1kwjh5t0Sn6dFRt1vvEnBNhgo4+Yzqnd3umQPcdDLUuQPBoqzI
mdZQnYcH2Vuz88xmWsa2xhaQvRPQZVxbd4heGGhWiuEGAzahG2vWREL6ENsnWhYCho7eupyH5PTe
trMF/hX7XXbXFiN/GffIddRjk5upPBYCAbnkAL5ZfX2UWjDE/XKExcSsI5N8qn29BMUWdOX9rB9k
IxIKK19auWwaogkOymWTJSKfWCxJ002kLvg+1rhvUGbroJep0ZGDL3YVheFf0iSousXmBt2jt0zQ
Y+4RtwV9Csiu/68hMZMgaocWQZDLctsYlq/qK5VuuDLgFEVkXVS+A9Wnh9HfObGOea0xeTcUcklY
fetRfW8BRQqD/ivlwiegSmaRFaDTiXRx2b0USSf37r7mDdMBCDZvsH5uTyeQbgJ57TVS8JVhvlAD
pH550FSJmlY3QTzNE5a1vlYRzJp5+QFM6tm5uY1JqnDjwfLxBBnysgf/BIS4LBLKiRR12bde/DtS
x5pXCaLPqV39S+khBa7JS/s0iiAO+LT6r8cppxXDDDfI7fsYrQsJtwUauXwFGeTCfom30jdbadcR
Y/6NL+Wz/NxtSQfNHdbS6co1Sy8ec2XD0lSWDkmZ9FsQreOJWRHcvw6A1S0Axmeq7VmCLF0zA3BR
wX3VHRUo846RVe2BXwVqe/phggwZB+pXw53tc6EeTs7DD6q6ltHgBfuDdPfv5xdOjN8lco5VuuEx
P7U4r4qoQKyRqmpqyV4VEgIxmVycTW4CNr24mIvm/3V62dTazYIXTvS7WCHz8+C/PXtgsexO65Wm
MCsXe/bfjYK8eXE4S3MHjjh6hK7hgdeDJhVOWaZ3t16yITz2KZS5ZmaYHKfwA7Bvs72ojSH2Jw+6
I6+fymPZUHXxIwBqJRtITuwGsgZ0Aq+LBn4RYuHA9hJKcA29ZuVspKP+XjbB7rACYILb3x+lWau8
2LP0xxOj51eS6uYPUsyjMzNQiYww03PSJ2o7Txp5bKu6O5lMwXxCUH7XPyOoeyWpZWQjVzgScsyN
PMJNBxm4Y5ERvoaF07+FJ9FuJ1b/PYemZ7w/dneTjtD17j9RpD34nt8MDxaPDhMPEaRaZ+WNbfJs
an+IzfC3dkiQN8AsPhu5Obi4drqVAVkOtJAm1aqBAgwE941mBVbsC5nK8uMLRdWnJvze7JTf0ycg
BgfsRd7hCCmuH99nqm3eiZgR3eOml68hLCmA9p94Pae/vy65DNpacbtI864cSGjIXVeRgDoV5Q7O
CTUDVAxfGk+X0GjP85u7Ae0c2aoOIon4aEFg5INQ257+Y3qGEpuNtvTlW6OrCYDB9eoEpPnxOYaZ
32QNCE/gEA5b4qqW5YzjQPSczRVLkDLr8owwFf/qrQWU+cBZXVPSvc8GZ6bifC4u1M9Icn3oZ4eQ
YfLsPrFo+klVdJCjKsZtO4W+ZRpiTuCrZsgI+5wa6i8n4n5tv7SKf/wQU6blj+IBc0sBWIzE80xC
9QWv2hj6rYz5Qu21cn/udAtAhNDFUlFFgzOXU9//b4OFH88iTmrDx+qTkoXqY5wPZaj286+CdAGp
C8SKlQX2L2A0ufa08S65VP4fU02x23P167RULfo2iHSYhguINg/a0sZxXXVglaNxV9xIuIPIu05P
XgKzKjc/DRT+h9lvMkx1OGMXhXQz0ieuM41zVuAxvPkMB9OJCzhU9JjAs4IHRjxgtHC6yk5Kc8Ac
6FXwZxRLUD4oWK2hzEqZUzkmLkzET+gjhshfML8q9jzV2b5TasTHrFSPqvZko7RLjp5QYJ7D6V0y
qJNxx2zOqXoP4apQIpjK6OmdlpyU/lQ/Iyn+Gny4kP6zc4jQcgZFwCj2hbuwJZNJvuTWZj0epwNn
8ssP/WCYikmCC4uMmze1PgYm+ts51ZN4wpRJswL3uBiPDyMhL8rCSSXQPtMYuUiNlyBSiWtzQVoC
i6Ie8Sf3QCzuoGkx2cF/RMl097qoRrPNO2CKWNVGdOwe44Dwje5hYywrwpvOtDrhnZDLZNPkHgmg
GfaCslQBnh2a/JXzdrtTHK5BNx70rq/ooIf+L7No3Hgk5epKzqkGCJUP25mlHjqkvb1z3Ccc4KgN
5pgv9qIWtK7zB7DG+QYSovu+Y4b3Iv7ffs1lXFZeMBPfvWFBcmuKC1C1oIhF1Z615bXfKXBIrsHo
+HqZB+0kyeYURqZZrLWfgyWtl6u+/xS2gLK10fHpismMnsG9lScugyABBtHPsDsvBM/DRIPjT7Hq
zXyMLLCgn+GPloIHM79TNf3TnQbKiilVHOsG+rTDVxGP/n4l8mspmU6hCa054h6vBL3FxRPhnfs7
JFG4mpwRR+cL2DAyaEBrdlTSyz73SBMzUoBwzsAQlFCHRcaA6R8yw15nihpK2TSxtyWVCzEOAmQ/
BRjXUwodQXSjcvnhl70b4urZ6HZc8xLX6/mqqFTZfduaoXoThWHAlh8q506bbVjnzKe/djmR1ZFM
yxNMaApakFwhtaCJ5FFfugbT55VzEpCf8pnwFZN0kqbHy9JmlDDQ12CTj7KvNRW94JHUKuKpuqcF
9f66hox7P1vTuPlVD8+4Tb0i+01p5oGWgYlNaNGvTghKMePpOjxtZ+kwhftupBSfa9I9PwyqLZoD
O6v45oC5d+aWBtmerWHyeOZ2nPJt9iJVfV2BW4cSDg5cpBH+EkaYA+OiWrRM2v/Ghp8U5E19wPuF
Mu9hWxt/fA7Q5HLOUTObhNmK6JMyOzlfFohUvTyMNYsYcd8oscUMCXxadeiN/BokfdytaEUJr8qa
xDbgjYxmWLPg9SsvjiJHj/j61xq4UD9lrPjtY41UWoPUM5T/tGiZvaqpGHCuwm66Rg96zAFLRR7K
Q/yAZtCMx04YhQObCZxbnMcFU3LGnQ61NAkvt3t2cwEKYjTzencjglpYI/u9g069eFWDX9F0bYEy
eTRESR0eEXtESxetRQuJUFHRJoZYKbRMX2RS5LsXycy75a/UGx+RP9MnFJTOxOezffatrl0gQB7H
12nLpDd9lXa6Norl99unGPW2ZuXY9QAXsgPjHmXbYConx5gZGuNIkMYFPo6gJd/jy+6wcUvmQkQh
9xkacToTv5Q9zuHM7Rqh5RcepgBWAhb50NgavhJ1hogqn3wxIsNke4GXiFeBeXeh41vQecXqPNnh
S2+DvIs820fbtXmnoEUXS2qfQCbfkJA62uJ7qSZWovSoPsukTJZvuvmmYvnIHYCbUuSjgpT/nV68
D2puz9030ZZLIG2IfBGphrzXY7RKCB03vIsoPvWTP1fOMNNmjvg45Xx/bRAHdDxLm8a+LMVdHjgI
1WaWS16IOoEp8+33xz8LHgFtOqEfLG4Tv+PbTHftFT8x41GTfIe5gs3C93AmjkarrdB2wir44ujI
1AO5Dw1sTziyeSVSSL/rs05j7p7xwMCYuJwuP1hINB6RaRINk0Gv+qHm82+TzXrq91E+KAz+/JN+
uEPyTN5t4W0VJ7Wtwsei0Bmc/QwyL8w+foGjQVhFb4b14Lu8BPol3R9WdW6+1ffGaLg/Q48qtJ06
ITPPdn6xi0rd0he6hrIugv7SKWaNs22AHHpQ29Ne25lB48Je5B0jvLmjzItDQ196wKON9GFHyYVW
AuSmGSn24zul5Iaze8wBXbE7hcvzc5LbFCYKvjdyvZ75Cav/PXm/DvB56m3OgSNSbc17oulQSOjK
pxQg9x73QNJsVp+Eeqrn4y5jhXny7wi8s7ksgj9jwZwrVVk2Kkh8I0aj/GX3n6XPvXrCdFrQWakQ
pET1rjZbiEYpp1DHfQkMrsYvwgjWAXP5LSF7uBQmXjr0dHCzP6LAG2SFQE3nXl3QAlqC5olzNa/w
hZXyc1Ab3JjXoMNvYho4cW+ACzk4DKECnjEX4TKc+uu7Yh6/+asljBLj2mvIAKsW00MAuHn2u68g
8ByNCr3HhwIFD6Hj3EpYykyhRK0uj/8EgMFRF1tX4lri13/oUT9veK5ZqNwwCNz+MHUTx7D9jazE
+9AEK16mW+cCOKED7sigbdCBffKHDGTeqtKb3ZLU2S043KRYaJhRaHkJqXG9wDR4ozdXLilSlO/+
Wp+OrmRsiZdNleekPxsi1ty9OuIOt6jniIMSZdoM0Bk0t9m4qaTXXMZSc920DEhkm/yXfYKOQZw+
7lrRO9TzxxMWXz9eg23fHeLLW+f5upY85WJG4/qc1f4nYTP+e9C8slpuILc+/0WfnCKdhUvN+s2A
O2UWdVLj4IA7qY9CSsmQufttLHvaAd3WSlzWmW7LjpPDxXgUX1zOlCzM3U7BioCF8fEJsGqHOmYe
NUG17ygJvKCZLPQpEmRLb4gIUgLer5uqI1r5BXz/oBkrmKzFKVwNIYbI6xXU5+IWEI9CErs9IFd7
aQDf2G5Ba66z6+gMF9kIp2mTaWcpp29sPVumcshMymkXjATiNJtD05sdUaC81+mxDm+q84N94rGx
vuzGqCj0NC2S1/rVT/wMIYbAKyuOUwllX2sCY5oLlYAnqekNbqHM//Xi3PnCtVwh5MpXNc0fnFSa
7yjXI9u1KChmAHAhs+b8n8o20mdEVtLBmgeVJMyYr5GBf53ER1mzXxU2KLLV/ZKs051PVHB+ndcR
HqIo1zoXrrIXfVGmEr7oqjqIswSXLMR95PZVlVpfwmI/Djp0rId5HcjrLClrsqrJ/Iwg6oBw9Zue
tCyEN9872JnPXfleR7UpbrrwhSFY9FPSt6q2rSKeknpam3uBzVkargCw13+eK6YqSUDu2pMjJ0Bp
Bhs8DFfGhvw1uDhTPOk1/ccrc9PMh3BlEWC0+XwyquEGEI8Mt2+EFIGgSRI5L+ZZrQvI7rFW63d3
cVPdKgQ5dryI+9C98LCK91DCoWXn0Eg4gwTDYgq4DTO1KltJu780CvemRfMQgcF63A2wHF4pQW3q
mQ2+6b4+M93GUAAyNWC5tVYcKJ0D/O2mflEKjiPDmyw1/nrKG7RpKMb1za+r57s5vRQI19SXR2CP
A5bPIk/B5FgU6k58E+NnPw1MvEk66zjF6tpx0LigvAV4aGDmOd7s5rFGAonvgSC1ZKR/W8kbgIBQ
3EBdxp4uEh18Wc18JhoPHRT8SwrCvhbxuZBSDqR4dCVLLIBBraF7HgypTDhkU9653mff9MQkQ4Or
ey8thFS7VDcOE7hzzGPIkHp4FOtJmKyD1+B5Ew7jPBXVhoOmqA0GxgFVSw6iv6JOK8B821J5H+EJ
QUHEuupicgDKTL3m7sXbuBPF4BXowEPilrZAVZ3npIpP4jE9OwNJJOlNX4YSG04Fjy39Rft9URp9
XTAS9fe7DuT8RdYJr2sbnIwn3GVkMaplazUFSvAXGoXOCrxJ+w4YX9f2ycXlF4pFrE7RdUIGawei
S3XjEEYfQt0puSiJ6jgzGKnrkhNY4SrQp0JBcwaNhyhpmU9pXBphi9YmAkMJF1MUcTWr9b1NPExW
YedqzjaCvZptvhoLFa8rItdqCkLTEScCQDHiY9uD3sGkjUMMUTgSBRAdtVNEiMFqt4bLseVIQ2rV
ENzA+rzf2cMfmDIesToCccl2gt204X5nN5bcrRLtXAGGebUfyJOwL4V3kY0hKb/IS7YEpNtskps1
NBEvG75IfHxuVJ10Akwwp74h6q48MIgdU85zHWFpb+qC9X3pCQ5/pljRsdv1Xolr7r/ti1TeK17V
YCUN0R7+q3es3xnhsLyJEgY6J4QS2LQ3J/TDBJrBoFgVGw1cOoPkTK4RZh/VvYZDPNxJVH3V2Am4
zP6A5Cj1ZdYco6hAzJDN087CEvXocTpWMEzzMHamriqSN8fr87YlxM5HHDRnBqfUUDL5GB1KJT1j
ihgnSTM0G1tmtiH1WO75xDw505W20jkFeEsPtkg0U2DviDZCUE9X4GlI0KjEeSBTG39NVysWedWi
TgnrAlrkvLji9CbtvLDnQFhiwXflFIvn1gq23+hxTpoSwHzBnzP1sdd998uWlVChUzofzIbuQh3i
pQyWqkOcV7tMUcsH6n7SWIfzi6Pcs/Ultxss6eP6FSFI4xnJj9Cbwu5oLDqVY0Lw4jo5ZfTz41HJ
yb4HsXYu81KOFiIVA1EL5PwBGNFE2bHGEDIMc4hJIJZkj16eSFBb+D186kLAbTIVeGODi07Tzo0j
Ll/qFnMbgH5nvELJv97tzLuwPkgbgmMBlqZ2qL2FlKRa+VC5oF4rF8YLUEltrfekocHclTw036W/
+yUjR8kuXHKwidpiwGT5/c6l/TN8TxfEQJFEYBhJBbYA+9IW4CpDW6mlELuClcEME3JF1zRpPVrd
0MclpDynQujyntBK01mtq8viXR/f0RWbAk+gI1HNUh1fJvGuIUiIi36byX3Beo5D0k9Vnf5WQZ2S
s1i443C6n64gOEP/ZFfSD8cGPI5oLqcRnFGnIt4P8vKSYAJhRpbbWgXO0To5Q12SZlVRnct+IPzL
KCoaW+eCP8wJACsKLyi7k91fFSzF11MsEWwg2MRFGpr6TJmbQ+Z5ooVZ56xhkb8z1dVpiGN2bVto
zz5DefgODi0ddR8HZHZio3/HGJXW/Jqr87fVBv50IJenqpyW7IFzXCL34ZV+n8JKIA3JeihnDy5+
BXPvdWT+UVv+fgKx5cjAmEG4utDxSAHTklYASqderRNbHOpfYnVkwoees3WuqPj0oVuZlndE8u5Q
djk3btLd4q0BhmHuwZWY/UmvvAnqCa45IbMAjb0BAimRr0px5vqTHCJA3LtZ2v+Wd63hHO4iqtjv
9tsvbVh4M4Z7oxoMDBq1acl/6rRwQaa4/t0huMRNqkEpKgzmdVOAfS37a4qre1P9naNAUhWiI+J1
sHG3QWZmJdHvS8YEXM7BGc608J5ppRQJL+KCFqTmOUVuzUQp60UZHUGHUm6PzQbxxeAAD5PBO/aX
LxUjUB+V+w716fJWEBSqXjJqx/JXAi/fjkZfm7ckr+zrmNfPpufgxW1d17q8NegtEnlEXZRMLww3
ryqj8ugOD3uAVxmBibDewutZoQ2vg75j0O9GsSSllBM/3Xj/0HhO36slbpyo+F12mTC4EGZq9mY9
OYLXaVPXna1TRHlAbh+cLypJo7IiTV4gY70YuQPT/VMe7w/mSEvsZlHvD6o5t9JfQW4zbQrTRIZb
ASgFjK/LI8e+4NqzkgVvfe8P0MwLHrbYsOl3bpv8p6lsMWlM1j7rwz1fjwQnAAreEtUS3wOqzMf6
T36DMIuDd8JoPU6a03MrEFdQ9xODwUCD739HQwH2ubwTzBJ3OR5IMVf8iXUoo2+8FLv7CVrK5Zik
2BqZyA3OepcidtH1bNPUjW7rOOKZvt5Vxr+WcEj0fL7o46OGkHmwlDfek3ymuAGmljfjsYSqEj5s
5w3gnRZxYS0eaoNPzEHvdEQrDJ/LdpR71y6vLMMKhi9ihesMMClHs9GSkx5O2252X30Yau4DPkfe
MccC7BNnjwGrDsq7aFut6RPByJKd/wJ3XT0WP4pgmY+DWGdgC7Ja4fE7kdz4NTloR/lGbW1BMEzm
4vWd6rZi7LhllhnApGec0Wynf4+A5RRAlZRVb9wb2WGMNewOO6GaEVTfcvCP/HFiotyjGn4eojhL
9906dVNXYPLHWv3PlPT5Xmj01GG3NvgDWOD5d749l33Z/coT5hLAGcsTgfFtkDAjH2vR9Dh44/Ub
Dm+aWbQ5QgVoHwL6j4i/a9iNMB8Kxz7YaA6WgybQBgHm3ase+rpl1RshzlwQniFRE8iMyQ7M5VYr
p/cNSZvwMhC7L5z593fljURBmU8MyKI2/8qoYhJiShSucJGucUvkWS77DRdr05PEEfo15D4PGs4K
SrRbe31EponUCVlz6z2P1XR17Kwe3lz3uRGDwV2cscHYfa6uwIpIyp+hLBJ075DYBdUi3OCBK3Lh
pnJVeH/Cnb2bSTi0cF62I3G/hMbeYVXbga2M3Sq6y9HZKyGPpZAfSTurhMI7GuiW150WjEEEaIt0
2KGHG261FkbITHAAnqGBBPTGR3hM04dYB7KBkVrbP8SShRTcQaTF8mUC/VSj3u7qrynLGE7CQ3RG
E3DcnOKqRFStM/Q5FfLTAkOdmxcGOcJjCebxcrBlFUhwjWL9lUwTHgeCrQXeW97JMSIaD4ZXzwVi
YbWrPwtNLswLKvrBv2mvdLnjQ51Ktsa8fl2JGoh9XLipNJfq+ggGbd60uZhvUvyC/JBNNA2DDVgY
wLAyiOFtYLxP971jnF/i9f+DJzquooZ2EalUbxJRWVOXXgW6qKvWF9qoMiOuUPhzAsoEglBodzdn
gP5xXLB7Jyf9BRLDeWfHOo5aptHl/KBjlY7JB8XNFAh2HTScNMpLleNavf+9MEEzZvzI22OHV8q0
LNyf6a6nBYx1BNnsTH5czHLrDdRizfxIPtlNFuZyk5VVNuAHlTQpNXZsNPx3qa+MmfYq8zK3KtP9
e3uyAnAG1QsmltYRhn3rsNthst/CpUgpwkezNQUvW84kRCAL+sjseo75SnGwcuUt6vLNLOK8iE1F
9IlF/RNTTaY3zuCWHiQ2AZVDvTao+GLeFXcL/Oh/zGyEtlZq++bTo6IDZ4Yjzbg6VWzOjApSAT9b
il+RolCYWUeffc1l6DyWDJHhPAfdDxZg5tLXbxf9OfppYbd0UIvy03PV8XdA8OcbuK716AVYVWTq
w+aIx+lv2Zxb5Iz8x+kP0hSn/QMCCaT0J0pridk8pCkVTbYbG4By05LW8xNGAw4OC5ApPMU5lV6x
iEcoNzieIUTgY5/TeDsB3sx/ILygE7R732Uq04PNDk0ImyboH2zzmRw7CBjspgQNiw0AjoqVg8sZ
BzfOnTe4tTEozOoAGq4mapO+Rwkw2MRdlNPX0+jQGfRLZ/SxUty75+wV9tbwPelWKF06mGvlSago
bR/h+OVxXNILy5on9adxjGmuf1IeA9PN8wKs8OGxZuUXTOTgBBbBIGpJ+x+dMt4+PIyCM/VapVeR
Kk2u3c2JYDAVavVLYiM3YOj3HfRZbL6nd7v0jJfgvuFAYR4oRn8b8hMQy6IfFX3VjvgwXks1ommm
c8EM7JtUbeTFEcGval6xlfEIM72EKa3Qd2cajP0yzV85+AIk2yi3hcJ88bAvGzCWk7XMGfT7NC/w
un3fke3+IP8rVdIG9JjHLQLno1FxhHohIKPcKMfaaIE64llRU1A67n1pBc2Qg1wnkFczizETm7Pn
jUNQ1iApG796URL2WacPURbeiTLNVf4H6w2NRRoEJ8xM4lTaJ2ktnrrXhsHoKL3eeS6ylNLisEKb
TqpGIqJ91JQ6XWpkAAMbQjAyUWCQ4/LQ8e9yZC0lhQJvm/dbkGKuTxTzhlrrYx/UQI0TultZZLqR
yuRAgV//TYovv1Nr2A/Locih4KZVAkdMoNjLoQCVEBf6nEOdFU2OcPDR1M6TrpmN0sZjxudnmZJU
grOmMxGArhkwBHlvFDkFQhgeZj6MbHOsAmUE2q7HrPiu2Zc/TDF6s0ol9jHPSHEP7GNk8l/Fq7bC
coKk0C4bJfxnuCt5CaCO6Dh3HchzqX9TPDXT9NAWA2RlBfLDxLxKeVHnB/IREAl+7fETeGma+VCS
Q1qlIfGZiRkB5Q8wtcONCbtUpMTZHz5Y/WO0/vFUppb4ZS57ldV6y/63lq8THiayZqDAN9yOqGa8
VDselkS6tpPyzj2lAbnomUbkARG6wQT2tlLDzuRFHTwWxZvt4juXiwdfXus/UW8tuWlsFtw261TH
acVTYDc/0wwVPHcP4Qqho+hiLeQP8mb9XZmXGvirnAwJQWK1MPbKrqkgg9PT9zZJba9db1YqAp97
6NOwBgatg8m3RX77CPzGNnhrseZ92si0ZNIAvAxpa+mLY2iLvUUc7SYbY8Ymef91ZvgEua4q8wiS
PyNeNxVlCi6Mo21dJU3NbNv7xSqmC7DYsLeROC/wsZ4wZuDdsXJxbMpCHtyKcASldU3hPEXaJEML
vCri9AOnxrArfPvf0ZPDdSfFT2jwbgg2RiO2YWhTijXtYWQLckoyLDjoHlED2DY3Nt9aIw+WMblR
jIGvV7eU+08wjuaLgXuNTd7qErmFA2HcObMaDwKZuFK33BG74lRQGV4j6K7YV7QxqvD1YT0k9+rj
2jvWO8Fl9U5NQ30MgqtZe7J/+ZdTxHdmOe2bPw4/yOrHB2JMLFuWVqJXZeytppZoY84JdQ8zltQX
qrDkR/ziR1BuHpB7Oh89dBmFbPxRFNwy0FwNbBY1GMAxQINrFKXsPV/xlfWAIDf5QD/wJTX2i/+u
yjDO22x+Bayb17naHbrE1uOAP/gBHqS9YoKrX8Oat7kAuHdIBsin49csyu/0dqa+tj9ew36StCxF
WniW08pjN1QS8vZ56sae191qT6u/DtQXIjfF2pSlDMZ3U6bXZv0cdgSWnTncsbiJ72IP1XMOBS3y
/9/S1wL1R3lRhCk6Dg9R0Y4h/rMEwwo1tfRjwOurs4jsjFI2dwBT7BfuCXmVsgW9Se92AKjFm2PP
9oCjCk/f7dKJMpCu7Wz177I6lFotAuQuraW8DRpDPkV7QpuxIPM4PYFm3liwmYx26YIWasJ937fZ
N2/Eb0C/9HoBDRRYfOpNa5uR/F6eTpK7Z3Pep5Tu85FOHs4yhIYfQr0C5lOVwtZUu3dfZzQC7GvB
eDmON7ZmvjQ/q/T3Vu6ZGbnHWb0AWuhJNuXO1kMZc234tp6yOhl+rwpzHvRRmcmbvoMQKUKDCtgT
RXkhhRPTZRXPZmu8hl1WC0N2pzspBLn3Xmx+7Y41DDRyRSgxhHZx5Hstd3ffkyre2ue5hHLJkwZc
QDIECsLpZN8DwbUCyCYBR2gLc/5fXChTwZa9gcdJewg0wwL3OWZejdapSXT2milhFZt6k35UOqet
Z1Db3YGLbdrtuKWr9MdvHhXi5IlHiN0GmWAqcZfLM6BaCkVA6MF+vGzF8WxeTb+EZK4vPK9PtZHE
X5wBNEQEtjtYbnzIqPlEMPXrvawkngde6TJdxMwAXNY0CZpEvmj+CkuhNl/8J3kdPAlh/7ynWOfx
i3UTLwgshC/mX492t8unktOL59X/5rxcQAKE40dxkoVxfW72GVIfRfxLTAqVoVw6eC4bLkzz5DVt
PZIEdi85JxiJ+lR31hi0v/4uLBVnG32q3qa+lbivLjnkXk2jEdPCqtji9+ihUkPyDhPqtCk8YMT4
A+2ZzbXHpfqZXtxnf/YOE1Ib40km1YHaCVXRhMbC+C82zQn+/EXHAkNiAPkOXfK29KSC2nWbDjEq
x/GyU2P63qECh6mux16zaJ2MeZ1DPbDasdnNzO7g4m8nfK59NqIaltf843XHqFfPpsEqmItn0nl0
CNrpU0rB0VrUMxmu+857AIvNLie4ge+XV0UT2T/u2eD+cY9ho2y7pWz5dNMwdBbHjMNln1Z3umj/
xkKfVnWc8erZ0b+zmjUAijpHhe8VNo4OBVssp8cFVuzx17mThz55w25cBMeDmzy9uq58KqaWNOSc
68m7L9xqmNaSGNBX9hptmAO14CXB86dr7rmei5C8h2Aren7Y2wUpBOdDkbSmUWa4tVYR6AFJjqhX
Nd92dJ3ZdTO7nSFqbVX9m7oNu27hNXA8gKFvY31C4FiiPB+IWhxmKIy5dPi9ejSql5HSdFbtANGr
x4d3xhALMfG9pGBYG+vd8yMMf9S6nrEhpJlKXWS1y3j5cNlGlDRXc+skPacViL51GqHPf8gla/pj
brLUFRfAXO0SqAEMbp9oyd4sFqzlRHWEGIQLbBQywRwBLN1VKZXlqrsM2IkpRWoioe21aR3zRs2E
atBbGJf3A9DUT2Ft6udkx8pxbMcZumL5fHCcItqJ3GvSLLqK7R/4MoucYVs10r/qo4ta0AC3f+3C
3wVrorW1W5OO3fkNU3+JWVtfBTPRTFy1p88BnxaKhtq02Wr+cAZoOW2XCw61f14dtBr0VFlD6VHq
FNNu0B/D7bwZzaq+4aYwZyiXLTbmTaAg58OXFSB1xdh65j/rIsKVTgyXBTmWbT5NH0yXHb2nD7Tt
o7Mpihp7ii2XnneCWDOPHl9u/xrMun8NJUpMCL4FZW3LlEphlL6xNztVEvQmh3hrpkoxbZQktgfF
L06yyE0OaZVVdiTMnAyebC73YBi5spK/qsOU6cdF6IiL6RIf7MFuUQAOkQeljq5wrlAboMN/O4y0
R5ou2rVFLO8BLlaLSY4ePojtbvPhovVGFN5z1FMKnwc7FBnfrkKMI5ESYcQeqFfne0pB0ndESJyP
aszOQdoE1d1sWO4o9NapqSVuU6YXb9g12Bw6j9XRkdWfNesiKIgFtv5MGIF42B7o/WAN8eOjc7hW
SE8M9aO5LvSVldMPPCkhhlJcEOmxaQTkYl9G5xy9WGJ6xk6iMv++6aAv81NwpXIjTCjvvv7dLbpD
6w5ia3GUezAZ4NX2pzpkZyKIJTmQSh618M4rDIHyyyarudvgdKUgP3dd+1lm5C2ungucRZ7lW8c/
iu9pdFQGuf8jNukwv8KK3bBvf4XwJGAz1BBcZZkRF4bCTEPG7TG8RaUv6r7tIEOczdgbNupSesrC
QIKA/Z0KRLIiYPOSwhVrpmE+RHVog8uYSIX5JRYu2+NqFK1H8H9Ga4oyEqpGzgR7zRSAKdmxfHuA
uk3eACS0TC2eLRStek5EqhusbfNro23sTnAW6XF7KOzVvHKsY3QLcx7Y+rPZmW3C+XJ0xRuVeYLr
8Rty+PXOsdFqkeZDalPA6GEAjrjo7YQmTANuFHimaiEo6UqHjXg75SM+0r6h2pfWD8eIEE2Pa2GF
5k2GRONzd3TIbaahuodOwkaW5qGRDB9aX5Ljm4xaHZz4EaH4hUyVNA4NTJMO5Py5K0tMO8D39Zy7
1lXitfjHkZaubqJyneSjyrrkKc6QxncseXgbI+Araq8E3TXW24BtxAfHVGS5smybHQiE38QgNDnK
/bpczUwYGGiF7j4FM+6WnZU7AayVSivKpn8BcipjX9pe9NUwVVZxg6uXXX1F7ArzNCG/o5aGBKTO
h7H/8DJcAhUnOXMuW36IQ1CXMUBUzo78ZP55BEnbtN5NnZ7Ng1TlE9SKMYCBb20l9CYSPwGSo14h
7rnR09N+/BdLQPidLpopkz/3sxyP9rtfMSUWFfXNHVdCjel9K8Bpy2aiNwBW8sy5VVeA6ILbSaEg
7a5NMizbke1kMPdXnFv5lAr9rzjcTV+MAT1VCRNVaBrsItcJgSKDu42ObNw1l3ZBQ7daCfZy/mao
uLxoqYvbng/Cc773ZRrc6foe8mGU77W/qUV038HL15AWg8pgsYTk1mSYUgeMZzsQpSnpxvKXKyrg
K+OhACtteoaoJEwhqZ6IBnhrT81Vo53es93GHfs38D1nPXsl2NjMUCEdhDsAliNHNV8sIgJydPjc
bzsbVSYPcCMy7psgMP+jSRt668G0N0AmnFXTg/Hrzw2lLTM8H9ENdgybqowBVOirpaEtgzMCBy3x
pU7C79U3bTduoA/WozFeg+GHifjk29vCcvfs0j2pnsZdMqbbQvQNyQtzeVeZ5XZa/9pGa0FHJ41F
YN8k2jwVOWXVqEU0ZyOxlDI4gIUyx8dXUZb5RQF8cw38MzmeUrKs9tc0QfrLaW1WJ5doWPF6ZUDP
coENuasi5Mx5lCaS3nZU2HOpn6h5951ArbjBeGFh/W95QmfOPBfgFEiNIArmZBrePhAImguUVkUC
+7/+phY59N2UQznLnumrGgKo73hf/vN6LRPayvofEVk7Kr52kX54kByFaXjpHf8f5BIofZCCjil4
YyHKv+eR0XB/NVYXe2dGfzHXBagzExmipHqazQxUbswhpKBqUwWtDf3KTf3USjuVkzrhUBh6x4FD
0tlsguOuNNHJxR5aA7JkxLbLzmjQv0jGl+1Dbl86ha+08/r45/6Myr/3+r153YvzQf+mmtZWcrYG
unMUsJDNBP2ZHxptNyTLVmEKEnQ9lqUmvW9PRyjqqGDkywxjMT67DERpV1ivfZfA7ZW44WqsZbbC
KdVoLBTnR3f9Qm+vSCh4rxUIdqvhZCnhqZC/WADhLFKm1BkKTcaTOI9KXDmihv8ZHLiV989qOjEu
OYiMpx6j0hCVLnmHpOvVQv+Jrokw6CvLqe0ABMm52ACfjIGPFUMcOgmQ4jpnnzKBT16FDHXxFf+E
GR189Wfz4QSokvHUx8P20tOMDjbg3Xy9hcZvXsh69SdSv4jO7OFBMAEPGSPr+uOOy7yWucbbQK6O
wGh3JoH1fgQlPRFnEA+/x9dQn0FSuLUg2zvRaBiMO5GXIMzn3QAp2DQXMkPPxlXLvc6aF4lt692V
XvEXZjdnIUU1/fnSYDNi1AlXjX8UE/WTTgqV0v4WmGjsYPOtUBEZC43+6UDoehvRBo7Puv8aO47b
m9JA3YMISxc54PMJ5E2AafiIjxAyE2DjKIrAJHzJEYkIdZ34yfpZNidXXEt8DHjgIVFS53SOoI2E
xdLXe8jLchdphCUkH8y70nOrMwlj1QD9LDNJ6aHQsp2k2Rt5h9Wry6hrgJcyD2mUVp3puVDfqIRC
Vr7F9zVE9DVYJ2RY4ZMAs+kaJuka1viuI+UVJEghMLR0Iw3fqleR163DIWaa+gapTlppF/gskpkG
el+kcs6rBhb9O/omtylypSTRsZJ3nkYvKG3jpmC2xs1w79WbLY006cgw7GlcEpEkHY2ogg1Wm5rj
EezHwZfaS3cxJcI4DvEHZgsfE32wDH1i1tqXgV1/vOIHw9q0IdXxRi2SGQZAuIYZ8uRsZiJ5HUUE
5vR2mnKsqQF7KKc8TDyWQ76eA6p7aPmWCoot2NxYrZONsErLFZEdW2XETl5z52G9rTM7hAQ6RC3/
IiJziXygRaSv5l3zKDWA/i7ntoKCwvRKDgPNufNxOul3hZPHhlDRjUSkaTXDd4mon0No0h55eGVg
7KJBkNcUa//IxNaghB9eqMBsVMUbxMvN9BJCs4MWNjGS9Uk/1EqVwCR6eDyfx7hTwOfiHXYxX5ZL
jxBIBmK23vo/RUQZ3lxpjz8TwMjlXEB2yMSQdutyLCFEOO+kICddsI4cNCVJqY1O6yh7QqbnVi2D
lZR35r76VbQgFTtGVtuBf2GTFr5De5af3Gjlg4Lx7gqB4mNa+lqHHVFvtw8I8aEejfqD69fQsLW6
IRmI+Ql8PJy7dm9X3yyXwkBEqgT/k0wRGx4ZoUNlRZbfKrKyT54YE/U1xbaYHmO99ILnPr6Tl0sm
S2lGeFH9OMjeFMvu2oJqxdSBu23hJZ4CFrXMrrCphxydhg0MpZl3yuiTYPfKPd/pYoXxj1eoRlEJ
weLGSmz7uyq9+bNb8GomunaX7zOLsbRUR9T3/A+dBxAwK9M8VYh38FMpmjo3ocgGGnKeGH1G5wRD
RDKKoHyxpdeiRV7XwxRbHT6R2aNfbEqFp/nqg/FX2KwjkPWjni9JJ5FYcapbwyGrxq74qMJENcd8
v0qaJdGR9xT74xdXnf7mgIGYtxjl1WXFRDylf3U/gwUWAWPRqj+VnDWJzstu17ax9PJMyOED+cuR
0TMTsCXMKQiPK8SZvC/YxHV9ji2LwdeC7G5aOJvtfjgcuG/4LiKb6CnE6ONnarnO9I23i5gnkTx6
YB87bDwNMbfuXk+VKFoFds06FUO9EhVVI5Ee6pnqnULFhyGGh7MR1QUxQnyebxXen/+F4pz3Duyx
weYVODkJJTkLwrX1yxoR0xbGOL81vJ/cT+i9cnDXpACMnJu8DIytusHz+lzLbqQmzuoCBbhRilR2
kf2B/ghDk48p1JsqhgWrICSf+eJyPlbh1NN186kCTil0eDPrPaoWJiYb3BXJcUKVIyD95vSOj0+K
AeglBL2xyaNph1yaSMcSW4ECQdP6RHycxoKm0dSiDnuzbbuQBIaYtUZmuzyrrviwdfXi7Q580rEy
RMsCNq/momb6HxkqzCJqxUT75Vwih9kIaMVnblXL+OYR+OqAvInjPe366K4kSzUso9ydiQ0OQ1aR
fCI/1cMThkKLAmfQDcJuB8uqvzeLAjdSOZYAeGtjk0Y12+Fa7UqUQU74O7RCMoRkS4y1t74e3055
EWg4uydlgrrJwodGx9pfZr6mmAdc6SzJXFPzyR+77f33RyP+bm996Rrl7IZACC0BNSjrZ8qoRB0L
YHmi3KZBN7OsoZuYzcCP2mvByelLHoOsApWsSnUFUK9ZtU63AZVHNGSpVCGIeA9dUKtqC7htW0Yh
7AoxFe8HoYAnxG4Lc5D2NfwHJ8ftOrpUO1LAE/ubP3b2GGjFgcpPHRNwePypeV6bHCRv75VeJzWR
cXsqw49HRMEK5BkQe1TN2VDYKD7Dg/kyRetGQqAyrWQsX8tyMJzPxil9ZCS/1a0Mb9NKbk3dsyq1
HRTStKDAroyLQVn0sTtU2FMJ/+VfnRTRxFoTBReuHhoIKZNgdo1U5DHXco7yC7h7hhkx51jg5g5p
CTN9rKDxWZMOEF80X4tjzWQJ6yrYYwMELg/2SXG1aoAMYorL0rDTY0arcUErCFb2iAG05C5s7rFe
Oxp276NqbRJv+y+BTG1bMaGXYswT5e92Gp4g+sjXmryiD6bkwCjJ40RcPVLN18ZFOJkTx7vjTJpB
gec+GJnNS5vhJ4CbpOaTMf8tWr89VyKYbEwRY/lazMY0vN7+VRWLU+QMb7IZ23nB8QBaPeNH8JeC
gRagt9WGRRCgIUI3vtV74QBFfw3UXWTFk48s5kl/IBwWoJo/Kvb91YPZ5+otmGmlKS/TEg6RRxzw
KIEBZftslRFxjj3CFyHDOaqCt+g7PKB7Iag8TVezDKPCb5CLYhcRCDhnnmZlX7G3sJCNgJNRmsfI
NzkcMioB4MU3XLaylQmhdD5TCOvwv1YEvDkh2JcN/zKjo+ecy0pue/1Ij76YL0Xz9dRjX5soRxYf
8x1LvwAmpfzFlfDzJ/Qz6Hp/ClBEEpk9gGvr7Uymt3MZqNsKQ59t7Xeb/sPgUbwfnHYXMY4dTbWG
ZN/+dbbSiJYe4iFbK7GNLY8YiMHVrjTOazrAOlSWXbYbFzeKUCaCVC98nrJa1GOMYGCkMOnXzNTY
HyMPH8r5KgFumGUYIe78J6RmrhLBo2jsNKr5GruTqzcwgKQCc3iQkWlsgJlXXo7hxNXruuTtvc59
aEANCUHLkhF9rdOdE8xQcedmIZRGXImc1j/TBheOiKL0Y2VU5ItV8DeWzIyx0X2Bcw+hE8HYVGzU
aGRJfoHOwzjV/eQifgrvDJELgRUJOw8eSNf1dO1MFmfhSuJihdsmndYAIVT+WPWFuA0dVdyV0G/e
OTLxljFG2FiQ9piKxDGKZbzxvbrW9a/XAGaOacK3Y8JW+zfgf75Des8WSpZgZT5ozvbt36Ah7s25
WYk5wyOsHO3ACeqiHfviB1znZYueXiaK360BJz5XjAHjr4V8ckD8Dvg6o48C5bSGRdSwb32vePEM
dp3zcLWOV+WbJ09BNp51I6hC/ndOViNzRvmxIBZCYzO5RcnOn8mzYOooPj2sHimvdBn+iapwb1KG
LOiCq54AdO9ZdBRJp89Ikb26XCOnce2/QAocdmNSmNclQUmPwcPD7CdOcHWD5AGeqOt6H4Xvd/f/
htyBTtg3LkrCH6TEOhqE1CafRcJY5z3YG2XUqyHxRYobgdVcR0gut2oEP5z5AfkMard2dEGSzOx0
TCyloLkHEx9UUkB/7rd/gxcRvrsi8+hVqnm/eP3U2BE+/qOetHC1X8CnrdpqxAOL5iqlba2/CGKc
TwxZOopYK8XWE2HY18Ci75D2cI5L17Y4oQ+C+7h6iPtWeekkRMGo8j2ygrTL+azYL2upiTfmuAKe
bz5JncvM4ngceakxENDrlBmyhcldkOyMXAxAUxTiwNa8kiBhvqowtQyx5AQN5yFToCg7hEmj+mwT
YwZ66n+nZnri2gbvvjeNGGzLqySRNftAnq8i9mjPZzx5Cgm4h2bOhJzN4F+lyKh4KCWX1K5Px5VH
mSYYLUAClw/ON6azbW7g3Se3NIlaJGLhQ/oCqr0UATHFt4c47H7ifFalZwT86uYDFlRYGsu30yO0
C8N8It/HDR8Cq6xUe0TmSmviDjmBYbEoLYj/lMxvP4jcRcHBOZLLdBbJtOTN4bmbzIO3Nf22H7h7
XLg7C++3+XjAuJBPXe3AOFYklQivXcUIz5gKy7S2q3WMnpbenXG2a29W8aT2bfuOWt3/0s7MCAYb
Z6FQ7EdCU+fSOgMD2dUar/J84xjb2Gg6TH9pNLOExI5Tt360/gW5DoRDLCJeyCQG/SJ6kwM0s28m
vJp9ZXSs4r3dzkL4u1FHGYXkqt7bbtl3E93WxnPnoCJSRmksRKCnefb1l2MzoEA/E+N5gAL3pgv9
IyYHCdcEkrhqk3EWxoC2YG1qDBzrnibnOS9e/urIIV5lP8RMi8M9mEY6EJcpM6Aht7iXiyBgDhpJ
MYF+TVwoNSJLAmVRBu2AR+ANfrvrYYBb5RQeeV1TUUoV3TEH9EOlo9O1+j6YgQ99ROAZXeIRdojG
WWYS7OxKO0FKVod8NlSpk0I1S0Am4/27bTwK75MFRUy3LGE836Ya4yIAnUPLP7MBtqdfnQuZqAiV
CY8ITfuUr7uVr/QY1j15ivHuP4emEoduqEM2tTq7KxTBkVFPnQUEaPQoEVOLCIrY31y/7NnlG6jL
4cEHEpStTAcUzb+Npd/2li6s4ED0gFMD8sA8EJy9/FqH89/sG+PKkCepBzExk5Lv28043n/34yGx
6yQGwu6bFFh5x2amtq1EkvgTM8xQJ8Ting1yyaeUxOFGGxBQbKJ3bbEVwyQqx7NEJnPjwHhg7pZo
ZyfeVZnq8ASpz2Mgufm45r38BXI5orcOy1TmKr0g9xsrAnOKvzjeVe7t0+oLwqPetLn3jrAkDQUX
J+6AehzitJhCz57fIxB3fFL0K7czZHqq4QfTb/KKRMGne1lbxvuFXIClFS73Vl8uT+DCEkPKo6W/
BL6GoG8jdhcYbNHas30nvFq7k7ElyomyPMQ3dpdrC6DAWlfCgf9F2qFnDgrJFlmzdrHA5ul/t0+e
ZlnBaz0hyJIHRg61FnnO9+Sq50JGZMlMDppvtfHnSWTIYUSys83UN5KZjdsuid0RJBsLX1c0/dcP
3iVXCjenGYnQTu5alc/8fSIiujde7YRGeokcw1JIsAuPEb38frfsIa7KWniubZN/WMRekMFrTTpe
pdXwPt2qfRQ8NOkwYmvh81vH/dQsMbim+YgwP2KS9eh2m9WeIJVWMpvkPYRVlsCLZHjwYl+e3oRw
xPe5SdOhf2L4AI2mCpIkCA30Ql9WssDhH3m1zTK+6Cqq5W2FckqK42Rb90teUH/cBWNaWUS2NjeL
5J6zqEfLkNGiDJ9qp2iS4ytjL7Ifb8TuMMjDqt2730qUWMEYCm5pkPq/SuAHKnC1UNINHLq+YuOc
22R0C2oVyxiOSlpRhMEisHsB8sVzTckac+iPXypdHjP9qXod75p7syi465usNNSHxeNSw+pok0g1
pe7YzJMvTGMi3/jYtNT5Xquc3ZpO7Ex7PfsvRwK+O2pau7aeRt+uHCU6yGuHCQVCSrZ6p8fsJP7l
FmfT3qgv40OAd7e1XdJQFy/j8vX7rD6kNLDUCMTD2nuCa5LJg6pcvkTugA0rO/1S31IWqHChl5L4
xNQAhs6/GgsaE+9J9iPDR81OxG1nJGpz/T1qo2hyj80yNQ1UHnC4YomgfbRHCYKmPloYPdFF8XCk
R39I0Cm43F2qZ1WHWRMhnQYgeMC6wpBRVSD7uPXXbS+Ay23Ql9tp2Njjv+o5fz/IQGnqBErfxpGe
ToAtYtJd2IM50x34MyYmsp5n5i9CfOv2Eb+krynphKcsRUKICaYd77tf54q19fM1sPUY3JHXiVFp
8G6hTNLQb0KF5GjD+M+IsLRN6a6dBMJ2HO5IKuZ4p2K7aEqzZ+TAlB9xTi35cP7mx3QElkljNbOm
RH8iXlZFmYyJ2K+L42JzT0yQ1MDAHsSnOpylkvDTSFSE69OaBuqyEMWI7ppPl5W8jgu15nL+slER
2qNEeY1vaCtH7NhimxaCPnMVH8zwkcSnq5ptCK/1rcDRQJdBu3cfaUC9vWgM59FNSXI1hiofaWNZ
LQ1rXdx27NqgDTPWSG1PLzGS4K8vBj2Z7zMAALmPcH3VPPrj15mbCPKcIL6ANwMw3G+KXL/puXbM
AEsLehGq0OmO2R/9mPNWh6bmZBvt9cf6Nb20rprpksGIzYkWWy40HYwH6mEzr2o+dUc02haEEisK
auXza+fwLGTjLEtzYn+xgGd/z9D+giAwV8T/J7KkNvw2O0fEqREi3kzyHOGd/WL7CHEGxNWsNP2V
HJRKZnhjYC+whx4UY6bK/IgzbnFcblWc3ZUr9HEs98uaRBpISQPVrb43/ESytVyNoefVSaoHacsg
zEpDsSUxNfqRLIaopii2kLO4t18X6xsJRbh5z4hHWjZeSvczkRweNDhC0pQ1liSD5M+B6/eP9dzi
8wcvvdPvXnXZ7r6mDMHKEir589aV6LhbnKr1rt/O5yxZyMCcTu0q3SR5EKRgrAq02oMNyiUQr/us
CP1iVfDBUAu4lJFPdK7qYK1/iX8WhhZHWehhjEAzeEdCgJB5/NcJn7VDeBEjVzpwPDGF6LpAN7UY
HYvNxnAx3HyrKUIfxxL/Bh1INyjACj+wxcutTwm+YExyAfE6LXkjL3LQ5IGqS0HPhB3ZB8xWRAR1
d+vstpS/fZNsMgJarzQMT64cECpEEDEScBdULN/JEp7HhAqFDRo86XAbznsQEtJ0fk69YCEfHmiQ
1tpF10G8Y5g3OFYtotu/9qPwPpqKa5/N7b+q1LuZLzSXA4I9ujzoRdKkUe7Y/TJMKmBV1gZ3X6xj
mQhBsLpZzlVD6EUFiuVZo3ZdahuwGrl+YcnfC22pOYqa9NQEOXjxyPSnDjMReBwnwoEvwSS0OATy
V+crNZyEIML6TX5jZ5SJg+BlLf+Pr3wz9Kz+VSiEXwpXIPU54RQQlB+MZXs57mVDJLL/3sxUozuB
nvYd5Vl/Om2s+azCGKG4fQwHwm/ZXNlGOG+0WwTAMSHzpSfkyTG13+2EdJXpc+t4Te6vZ/qC/KJl
Ayjdq0IrJsig5FSzQAC0iSWX7hDdNg4qPTsx48NbRtRxoqwS3Dmn3HxfszU21FHIouwH/+QZiEy3
hVq4zvBkW2QggIAmQrkWHkb3QEfdrglunBZxZ848PVkEC4dHdFWtZmTc0LO1GmKocnQWfetwtGol
4kcv2Fiw+JyVI15yUuXQZMF3LO7Ifwd4n1kIDzBw50glh0VHZ2CDXnKr2npFbZfiUJSRx9eduImA
KUO/K8uRHLV6OjbWFqN8dms8LBv74DKRTc8zuCPIZR+2D/gQEA8QHDVcGwVY2knCxuN8hVgM47bl
VS/o21aGTbef5erWzRlVGwpa3UGgjsoi/eDtBRGCmFareViiAdPfFjGIim+pQxE9tzi8dtOPoSec
PXjpOgRAd+VXLXLZSp4xLS+Xe59KsWorxWqifUqa+K8fpo9JSlVAIMC+urAraKqdqFwariy/EHMj
8Ztq1EoO7pk5QNDh6JM9ePWLmU4jTOXzYqQCJ/BTkuoJpkq6q+llxD7UxlkcyRjrm4Cm9pv4IpJO
SiY1s6wFhcIJIG4Hp2cKZRv0+/QdCt4OCtG74JbXHobtQydflbDi8S7qp/rMacXWcg1AL0ZMU3DE
96Mug0eDhvSVmd9bsNBWjd1VxEY89GnijeXbfS+4gR7f4C2hznkEuIPKhpnS4col/AZuZtfMSaOh
nidhC+9vh5RT6qmlN1N6z+Uesrs9Hnz56Bt1rgwGnuS5jterp1nzO7NODMhdbGtoO6aUGltlPVvU
t4/l71di3CWayVJEQeu1ruE5FmuyyhnikAHbTw2AGdBkJDLfL05yydV/xA1hguYNCWCF697udBhG
CiwLrhxyo1tQq5VojxNYWxzpaA0fawFVTDVzDSfKp0pqQd3JzY8tVcWdA3x4ZpHe+MmUoJaAB2V9
fTL0ocv6c1Tn0XZUGICFgTGFaoo1jTkB/PdN6LmHy2466PUSVgnfu/yyEOcvn8MDwkeY4YNp170C
pIThm5mj96QgSK5BKkUFqNVBaFxByZQfp6Kn7SPTksCEGmPZ5LC7hfupBlgmac73uQXmHfJZB2EE
Dp7E5gl0Pt4Olf6NZRFwssOmyvSprCGldTPTnAMBiLiVTy5h037EZoq+G35JQNvKiqofGb6Vh0fr
XZ82VnkEuLiCX+XGrGy33fGt3En+6pII8WD3TrMVb6VU2WsURTeuPaNCpzIxzNnQZrENCQbC0Ovk
RrHwOAC0sjZnjk+Oz19QyKmu2476vw/PRwkHvt3FkG+a+yXqur3mpACnVL04URHAXPWDrbibEb11
3yTVeHP8TrRJKX7j39EyhNobcTaFDS7PaObO/gXpFD1NFIRXSpUP6jcDiuwxd03atMbOINyCNaKI
OUGnZx7hiRf4Tba9JEW3DLydFlDuslvkl0ZwJ8o0N04VC/WaRo9DzPAMa+H40zjBriG3wDAsFQLV
wpl6+NLC3cQGzU7HdoMx7RREC4lEu638IRBtnELyPfrqMvOvIrTB7xxFGkvu8CpGB7ERt9alB5eJ
8EPUdNNtYZK274S1ljfLwuTPbDeAGa+nCLJIsD8PsGUYpTDvaHkJQ+llp49MJJwNHeTzBdygnI4K
+ABRtC2eGYitEs3OVIgvOLZ4OMAs+StAzwyqNBIT2l1MrvaBxlbHigPNf1we6jPLjS93Y+Bm2Yfh
R+uhY/Ock5lvsR74nLNVtyQ5tG3x1dQAOnr3jyZyw5cExUgLP0Z5/I9d7w2Mg9V1YqTrMm2MihYC
Shf0ZuLe3D81JFQrmFacjNOljSAlSZ9LQ5uZUm0UJcXcRJjl/PDvLiD1I1zTz3rZnbcHP47n06R8
GR4w4ZnJElKx16sL8r6UPv6o/jDsIkD10p298+xZaa+ETUDBrXem3ZBWI10ycklEWol/XnBRGZov
8wXZpBdhUWSXOUxCnXJQZMtuVm1pOQhuaEdlpkl+Q8CFTLMijHr/uCGa3QTLqcLghsNd4+RypfCF
nlPELc8wM8kyo2buduKAErVyBa/2N/oATUawKczX6oUGMJYV/vlBot8wvV7S9TxOe9nDsMLINExD
+uJPYUIjf1ekB78nyueAtUmMhGpKZH2qB7jfIsP/4S9MEK9ranC7W+ZJ0aFQHE58Bp85BixXggcH
oGwaWA3gFI4klRLqyaWW8UVyDhIoBIFjnUMcy0EIFbXQd9tO6dfwRIcfPp+acKA9bKCJWm/vRgc3
IWO80Mpb3cCk5ZApk+Vr9oZhpD3wDuUu7rqgBMkgxtmUTuSjeUVU96KJ8DEwpA0z5WrkhBXH4rMq
iJBwXRa6xZAG3drHKQDyorSCLk/I2ODW4Pvjd65K8pgG2gttV5I2jlbwr3J5yhdOoqt/WVZSTs1l
5oIT22edNcvcGXGyMQHByPKwbzkz2PmH/UJ3AFBTeZHgfC+XqMLB2cXH7Bcas4fnAVqnZKm7hqi/
ckpwyPW85mxdHi5Q9m6kc3+DvW5012iUL4oN+Uz7vor/FuMmZnmctdWNzhYZ5v/uZ/9LMdPAStA/
6lkWRAMzaux7jHPIrNHobaDr4pQ8M8BQjPlJonEUxZJOcXJxJT0FBpoUJk8MqDBXa8JWJcwoD6Tp
H7TvqJXmUz/h0oc5KMg2KJ0Adq1RZ7I0QgQ/qDAgWSiV5PRCPqtuCA++G9swlluHcbk60dm5D+lC
h0p1s2/284GUz1rSAP+ApXzD7ngklYBv6C1wK9xO/uPPoUMu9eGus8j4wSrepKbFGdvMdoG6LMRJ
Y47tt9yA413FhvFDL/D5t15MJZD/Lplna+cQI6suemc77aXxsHt1ScpNQtNPdYfoLHhYzNJro7nN
KADHIx7KO7ouO6VJlikt67xdKGLI/jfOz3KjKn6FcSOXN+G36WTsVkAc7Nmi7scUKrxYZ9Hn/w5p
GF240h98FazY1QSgqvXpyeGCEpXoAro/ASVwv4zzXDpmip5vpjq7ZsUwIm1X11nat1430Qj3H2Ew
COWbha0KJm+8KuutY0jUMU2azA8cpZ1X2ozaMlcfpHur/JR1+XlVCJCFIeAoYf/DfrY/bcJBl/eC
7TnfCRl2QHIdDf6qjz7rXZbcDgrQ5eqKFlkhCvzc7dOOAxPTpYwP8av2j/ctUBFMJQldVpV0cCv0
IYRn4jbD5nP8pVDoAKP5/H9p7KfIBRF6MXm3JKZy9K4u1uIJX/Btzph0qGxpUzZWFJXkiTOiEMLX
wvhNEd9KSP5YBTIfy+/SsWjt+vO94fNi8jhCb1HF0FaeQQyE39lSvDJRHTWJzrzR2b7CHYgCaEQG
1NNb8IZVZP7hxzzNnuZ1emyTO3bV5tj90i4bCdAYvDZiWrfU98TIlmJyoKKHFNVMNkZdAJZLucgf
RuYY3pSwI/k4Bp8yWmcRtoccqDS9wrVmfPzSImzgxWm/RfvxfopU5Sf9wLQKo6mzzzi3/6dlAcbV
CqDCJDhiCQKA8K7lQKzamlm09x8qsiwD2sK+Kd7zyp+902icarBsSGsu0AWDhQXy+bq9DLpEAm6I
lfa5MPpqWS4STctX5QEhcjHUAAwZC/ke21QSVdEV3Rfy8HWdPX/tFwlvUlQKA1iiDMMuvssVrjJW
620HxxSoUE+Jk8zrfjjgEIPYkLpwsg1SRuUJNRg+AvQ9a1rtXf+ITgUJ0QBUbKBo624ooOILgLzF
+Ees43BHUniVHVg5VtiHM2libC0vwaLqbkeReGvKTDg59c34yPYMUdcHJBNxRvtfnb4+MrQUS0oY
7Q+om3VpPZeY/oabLvLyTk57xQRjubJBOiVfqRpqt+oV8d/56YQ7pN1UQxXkc53LwYiy+PwzGWKs
PbRVBXnAz4ben5JE8rAg+6WRPe/5eAhkPMtEdXGEZ7GdyIPk6OMPhpFFc/1pMjCvZvWU3lYJ5zxk
mlz57ShEvYJ+ql4Qw/nuSCam6WZrMhrZT+hS1BqipcrjweofQwqlNM3Oz3ot9SRbSsdxf1ycgZgE
OcoNYDg+IBWuT9h5UY2xglEVHe2w/jNsrCt2Zx85qlfRPxmkHbxc05WXIfqqqBBppYw9GfTGZM2e
KHtCr1cLUggONpedptsEx0K1aAiZEHQ7gTVhbr7Mh7bcU7p66H7v6HRC+fQezUnM2FU4bqaUbCdO
3rO4lAtYIVpQ/rTCpiqaHB96Q+OayO9kJXx3H1Oi6svN2kGjXMyQIvKN3kFhl6rI2b9SK4nMryCW
XbimMfm7RBRPEC0Q77Q8x3ctRfFF9U8E6zRNJlg7gvte/LTqJg4PepWEQfwarWNFr0r8lwx4UOiX
7a2O0EIwuB0UwLJbyFvOEFAjftl9Um5K6hve22a23FWFFte5/dJpzRBa3IaNPKLUIc3bQUk6umTH
NCsEJXqnWnk2bvyczp4aLc/zokC9FnFYwHUuNGLEwoBMdQ8fQTfu3OnR4xiipOCIAnkSM+1gFiTu
EWYtyxMQkrWGzLwrJ2NtLCcSLKQhYDuyMLe9ev5airy9+JuNfY0PRO9F6m9VSu3KqzeLqMErK1Oy
KOJBj4bxBjWqjHiyXy0RZLhUSuifcAf1nP9G50q+K9FDwpsKOMvNumEez4fGk+HMXNG8r+YWQrKl
Lk0r3fxyLNCaG3QrGAqc9eVcZS9A6BUHbmH8/QTDhkXX5rVTgVDJTbgj/O7SGvGST5ADD50JXlvs
caICuj320c3JiHAFbdaGsnKo6n5+oCOmtKg3ilEXzcVeqQ2D9oAMKPWLt3dNSaec3hOkHGiwIf75
WtMyLpB3dwfrHT55I4ofyN5glxBRLm59qAXjC6R85xk7O5qAezk3J+jnzvkipo1/eAkRMImqd4y/
iC23QNQY1KkBRw7L0KRshmNtW5NjYOiCYP3nNRKEv0kz/E/wuP2hFU6N3mpgl0dmULjp7AQIJ9+3
IGEXXB0LuXaQbP1egGJZrZZP3EGCZjJ9sSbXws/DIWWAagBPiOIJ/wevp5bxDL6Bwke05IcHaXqB
uTQdnCDtELPlCQyaRk7Pg59TwXJ6r+D6Mjk2n0EuEm2cBKU6ub5ZF++DeyNs6kiXppptCkHZtYyC
Hq6kCEK7VYJy0GE+uyT43bAes3POG6G4MPweOGLzHtWUAetU8mLiVRf8NEVHwz5tTZKRgBY2Cizz
kevTyaQJu3NhEUrhT+hOYU2dfc1VgvGy3sP1Fn44jx2mnFAXtc4ziBJneGcqcpE1U3ryNbEx1lGu
2QTGqLRHUSAIDQtgtORB+CPBOQDD/eTZLxYgGZ1DtpJAY/Mq/XgR877iHsa+A162tWX+yQee+FGy
+S18yKfde3vDV/NkfdTNC2Pp3SnCbaSm+4V1hV/kkEJy4X5hAT02HH1ueZJ9C5ymHqHrBiMPaibE
m1X5WY1Bx1mh9WiUKG2fdBrNiXDvayRUJ55e8WUp85EKdTDDVjfE54jATdXAcGsLX6+0tLALO97A
zpgcB5IWi/T+lHzNoZ2NudGE8ILJLncz62ENZ4nOaEs2Mw6vxiZ4Zc3e0IqD2HPImVNLUsJzZcCD
SzK6yRYCC3CDGKMGbUAfpVXsiN2bUxvzfd6AGM838dfyaNZr4o0eFSAsaBgpbsNGvX3B0roEAWYS
RvfhM2/0RAOMm+Wm1MOgbL/GExUm5MnMIg2q6ELR+L9Oyj5H/paevmkLl9k/ZSd2fEUYCq+nkWKU
ADIkobzBViSn1HlXa2kjY7waf6dWN6lJ0qatbSJLvrSdSehF5Q13jVSviCPqI/W/iTL4WnnjPGcO
MfQyoZM9GJI4/f3IGiJSsa6BlV8aVs+dMu72xn14GaYlv8gahLrNWZCcvGRBzbjFjUDVMRigYZMl
Z4/ceewOMatYBym7hvuz14e44ogfHSM2U+PeALGJU2nvSU97Isol6nf1fUL1a439nMq2KsaNlWNM
rkQco1igInqo5Hj9s2pARHn7D4d61lww4yxnKD0w6lIPbIklWARCeKuuqim38wqwC+Wmczvta1OU
dRtRlVse/UznTxaPNntb6kTymd2c06ucJJzC3+UeS+zWSdZgVWt/HbLlT71Z2ydSqgu6u65Tvxu6
7G3+z04xYydun/7maLudZo+kUwgjE+jS/nmj5c1ZZ4ebJUcAyjxvWg/oey3Y+8fBTOH+4FViA3zH
8KiBznrPNjOGbC3fDksmtwM+KKcfok8Hz/d4wUjYqr5QqylB2TXSWIwz59cBR5tIISdWoX/96aSm
dAjJUZ2z6z6BTR4WTbDuFiXD2k1IRSf1orcX95jMU3ASWuy7/eJc1FTzRbZAhqgSXJxvCy6ZmKe2
wbUjPcekMaX9hNgQPoO8P9had/fmCM60oKCB0gkdZe3ORIyDfO3inP6v8owPcNMeEiqXyrifCt2a
mjez+I3YznKhyl8RCvihl/3vFcuQh5bz3zhRC2TXnt7VD8JL+xx08G6sgBw7FSKSdmVNo5i48IJK
9ticlYUQ12g89pvAQO/zxe2TAqgvQPp1AHrcO2/DvLqEQwqfgrJhlkO6DaLD83GFCl4IudwusCHH
M8Uhl2TLbTV7JIxIMBVLeDV/K6nMiZO7mxu7ShDhYZrYQS9oVNfqtYUvLmRLQF1ZeJrBDRLWf2Gv
zCnWw2NblMJdPItzSziCiyJbQDAMXxlanf0rCmtrf+dHoSxkO1tQQx+1dWAIJb1SbKTm6RBW+WFj
6UW+AXsOdZlwFozx7VTEZKhbxmSeKUH7B6kF4kVKOq0CWHLuLWmtIF0YQEGNgKz0bWIFZ/na+oo5
JU+XqUA6cHUPAWa3xemDVi3gubS3BVvw5gR5eW7itj3AhFhdSeQKNocvrrdPVQKVHXynygniDIT1
LL8W5k52oPoC89eWykACd9iNlWyvtKOvvd/PmS4v6NWQaDKckF2cy74Bmrvhm5VkmPVdtReZ5nnJ
3Vqe0fAA2f812BBY7cAjCK+375Dq+iW7eea3AMIukqi9eE5Tc6BuVJpHlXkK81C+xYHyuxV3Lk2C
H2pQvt0K6EUqVfxJrW0HXlzNKGKaSjJtxBazoy4jB9xuMacSTNBdrjdchuyPqR5rHp0S805syZcn
lXEPi54oi4qrm4VMfMTzUzCoCSgM4dHYhcq0vPN6O1zqVG0PJbleW4IWajemtkWax4RxeSoBUleQ
u/pKVXTOBbh4XOrqhp+ubCvRnBfIypitWqWEDJkYWA2poO7I0HzN+W5a2iGTtYXhgI5PV831vD/Q
OA8rUyf+z6ZEug0xRgNs3v2wr4JdKZWX9M0nlKC35N3WFM3fVmXo+Sgt7WfbCCFDgQHR0tlFV8KN
9pk7t/+LOTt94i+SGUrbwHxtD2GZJBz4br3fZuyQKgBu+KTrq8kC+sytknMrX3lchMRAwe4TBwGL
isnjuQJHbyR2ayEl0iIWIR6LmdDiB0Di0yxjjdZ55F7hrIF61fhfgF/DElWBl9gWuLVz+j3cKHYL
jb5kzL/2CNz+uvK8hFJxbkCsb174fYhY+8yHTCgTtFKpV8OtWBu/3hxMqx6LmaUDeGvv4RtJ6z7l
gJqJLdxfHeDBXc6/mMi9JDQEvTFyh3Pi3eC1iFuzcDyMKe7ipUcNkXlqz/sVDQ9fCdXtipChIDUo
6zrN0vC60G4Jaq8l4OLcQHpLWLeVZZPSsC4TQyzpDf91f2zAlB+3jARj+zbl9w4SaDzOzVqO09eV
lxY89aRjl2s18j/cKewdbvI4ZjTb3+06DPYTH33gVYQDNwzTJSO+jyiUZrnus2+yWIu0TX5m5xkT
vKOQtle/ZnQKwxi1HVOk47JtXHEeqaklPG4YxHXdLtZ5pVuslRVCfkuJ1FTGTv5XY3Ahm8DzO0gI
jquwgfx9p7y3+OV8PTtul8N4BsdyFqAmjM2nVIMeY0eXutyJPk8IbkTrU/XLoaRj8hj+CukERl3g
uMnranY6Q2XVnlA2RLdsqn6MJbyTGQQ8urVoMVzM0P3zmHJ3baa+N5ljlzu0fYh7NnoFu/l8Ow5g
a2uYRqv7Xrr4L6R2t5no+k+yu4tcZUQhrS6tQ3ty6sFLXsjHZ2yZMDaVxwskGlgC8PRJvbQZZXal
eMN96OGz9DO15C82d4pVj+ESpu9OFwNIIFMFQVuwiZyUaeFTAEiKysSlZSY1Y4Yejhl+TMK03jz/
J+oW+6rg6hurvB1itouNpna+YxDjWORu/j2NT+ICbjNFqfrd3TriW/9J0OGH7ofDlxlBWp4GLGxT
a/DfNRQk6UcNxhRTvoeP5GSyNVdu4qchSjms9GQSS3+uSB4ldXi1mQ/ARE4ZhAiv8maUyD2LyVgl
jtEXX5fVXSkfq9NPj8f2LjuSy6Lxo0tnT0NjbVTT6ss2/XJaW69J769cCboLbampRheUPlzEFy+5
sRlLtbTsQyUxqlsaDGUhta2rvvl2JGgnOlEVQ18TS/8eHRkumDz5x1IAq7g+tKL7jLnu+2GN0/XN
DVkbySmUvD33izEiehS7aXbQ7ZFA5397HMcAnde1ipxIZ9m4WZkyq22bhhc3IjIBSgM46amu8Q3O
y92qVISJwwuLPYJ6Nk3ixqR0PsxmOmzhIoOuN87TNMDIqLturEE2gstp4s0rzeO9DXZEZ6NUdFyu
sEi+bsIPl/vqSENKA23/AD2olIcM0jx6NCyrpL0l5fMnmE9JBqhqQMCzJEQPZnntT9BdKlydQFJC
GiXbyLFw2grfw6toSwgDcldtCz/4uRgDax+O+5NRf+N5T4/5/uTeqoHYALpZ0Jft9GWIDOzA/7x6
xTY7k06UIeb0M9vMgUPCO4d0EXsDi7A3ne3YQvtAeNxN+UR6vNVlD3KcSgG3lkZQxE2P3DX79AJ8
zL1YB/RLhoYYp8KRJk6lhC1EwU8FxocXKcgt5qoH/AQ4ZH5bVeMYThTt8HKg+yl9VCmX0pvrWb+u
FmwufmctlITWrNXFuJ5pJIScJ9JNa9Yrqi3hq8dW6p/ApHED0ki51NUAt7L+pNOrkJtfGxzs9rRl
UxLuE0h4URM8kG/+UphoBWw1z6SfYBNXqS2Yp/w+P/EAK3anXZ1GlqkrrJinj2AgYqR5s1vMxU47
mSvg8wHEoN08z3Ik4gMwvaP55i2QHJJ7H0tEGS6uhjkbdinZpCrbnt2EUFKmlXwmxyNb+XudPEMW
WtCRPzDpH7KD0hD2GSmXC8n9w9XNx2cMhbW1ituASO9Ao4lvAByRj3jXhaV5vjEYHsuQYiHpdT7H
Tapjny934WUPagD9yC4ixxZ9YNPLwnUNiMCu8cToL+mf1LUh4JsjsC2gqnJP9WBwo7++oqgc3v6n
vyRF/owMhPBuqpV8Zzfm/tkNR26HbKK4i8N1u41STy04lD5GA3uUxwMMRJfwdwYur6y+GhePpcEt
M3aMBMBzg7jWZVAJz3YwCx8eCI5MMTQMYklcfTfETQ30n4g2EGcfO/drEf7vluGvgNM/ElmgLcTr
9f8EmSom3HxEo2HF1ENFu3l1FuddC81NSrIyCMXNxF5ns5I06Km4Nwihj0ivdSy0SxDhdsiGAL42
n/pljgTWvGb1hw/ISMp2DxkYmU2hTcLBk9Tv69LYNRm3JIRyCFYg4ZU0zCcdG4IVL2v+6gwSbz+t
NCb7wd2lNMQqdZP9gSS/ZrMO7l784N/csvlAeMGhenih8zeOXse1kLbm5Z3uZWaw0FxfaV2SBL2e
E4BskQse7pt1jQQ1Ant5KSiL/S42RIe8upguALFRD7bVAk9yrXIIE5SndM0SvGyNTMNxhjYtIseG
ltJR8sBv13/JrQFVS51wk5KX3tZBUrCAONUiHpi7d3qnK9OzLfhSF+O2/seKdoC4LIpxM9lI1lFD
4g7yY/H7D2kJ875APyI1CXtoKyPquV2HafluD7KjDuSiMEjYOmJeifwqInaif5eV8BKgV5D+NNk0
59oUWHyjS4QqN9dxkG5DQCuvGLJcC5uq7tCVs+BvnYEcI285xWAdEVtVvLzeLv2Adi/+jqY4+uUz
b3NfIEuzfg1t8JpNiEtaHjahZf9WpQ5o42CJX6lnrXFJMwapwUn5AyE/MZg5yKvW1zYtspowkCbr
WUM/KppeFO4SWU5fEHV9pIC+zbRdcUvA7NmWI8o4ipgjfIvSG5jeqFkEFOQqPTXY5XN64l7hz8B7
OzvJSX9FhjOLD7oNWLKhtCkGozwRB18FsTeyZWUSA0ieWLRTQu3YymfFVaUmvWzWCZ13KNl48PlD
Xn8JUgfbvyoW0fhM7l6q/mawOwLDzVUy/lIhsdGzkxe5yLNhFQMHqTGT/UyBmS0XaSsP9hyfDuWD
Ny0vlu02JqqxM8pW8MWvNoBkWwt5RD560CkLBrYDUa2mUS8OQHkBg4O5RjLNZ5CqCbXURPLbttRQ
mOsbmBMd+bHCmqyezwq8osQIrQTFFwsLXAjyoEGNx1/YTh0JM7O57Wp9IpiS0F+gQlzEVOHZ97dV
aYKS7JYR5Nk7KUOCfvtiO6/KMo+I7WYv4XN3c60If62pOUz2iDS8QK/IhX/ZRFMY8ManVSJi3/BR
ppDDFsewPYiI3hYf7SscQ/dTEavLFDanLDIwNRaMc8K0KrEtIVcco9ATggnNYbqVAKLWE9k7Bpbv
12orBLMPYRgyfATn4sNvFE3uLzgbYUZGrRfRGOU9vy1IcJ8xoLOt3n7CvG2w3bFnqmCgGp4UQwqO
zjE4Kc3KmG5iul44twEgOwTT8ONLlggG5wPWuBJQe56mvwu7XRHj68OvrA87JHP3FI7Gw/Ns36hW
fOVagtX0bYoq3rg0JXH5QC6bVkKk2oPRAyEsH7VMWK5zr5bFM2a1B0MtEkfYl3lF5AewxLtaDzY+
VdEQ2Syj1p6nplzY2eUtwMr6SgUX/Dn6PsJsF4g7xV9zmsoCdrhbMDbZVmp+vFbX3owahaF5vzg9
DjtAvT0tT6NkQcdNr57oS3pMeiaRyucqLo0hjN+aK41B8VOiapbmYXb9rbvz6yy7RYFI7F0/P/tJ
m0FBGkDJewl5PokwwHTdbqBesimphJxPDv1v3igvVnfrQ99S9zERPTj+KU84hSR0V6E0SsZ2z0Xb
Hg4Zs8HmU3oirOL2BOLPyloUuzILSV7IDg/ByyNxIyOZLiOpmiqYC2BTsp+UihR/vpfuz/dbx3HX
xIGUtVYBV2iX6Fl7+fOB4V0BWUoZWaxl+aGhB77Ud2KJoFTJp0l2oF2T+kgM9XotWZo8uwnQ5Bja
msLz2Gm57mCIuar7mQ7Z91XMx+L0+7dj40pMRbJ5P9tDER++xx8Kg3PLtS7Nr5gHpzxsh7Y9VlTM
+xkDiYqzUiqvC6Vrm2HcUgoP9rYnJVg0Khh9KiqvParsjgJFCO2lvRLaRuMFOykj3LqLnR9cYp1b
3DhXYx3Zpm+1PYQgMS4WiJ+qKY8bd226xdLVPxZlZXhCTvKVe0XPUmGLvaQnBTKa+BPXnXIbhPs0
S9a1t1z8iYubDqMIhlxHm1Y3atT60kQcYRu3kf8o7y5bJuTZgHl6Qn7ZqtbsbakxfOv1GFIJl7YF
QVCPgctZbqS7jW+HuiGuNfmrabYu2gJpZsPqnhfPQ59MG8ai1hA/rlHoEubiPbiobE/n9wZJrSLm
6pZD+m1LFnXN6lzgslyI48K6O3ndYTDPb/cCyKwUICJc5k0Ehm3PSTlRwlvfsKSWHsMAlG5XsFg9
OcmXDdPn7sndR58vdwIFacI+P6r05L32ZZrrh7BINkFZ2H5nd2ao5bi69MZUyQdkllvQhNpB4TIG
jxbj93IXd1OmzktiK7BaCbMon2Odilzxu5wprrYz1vK1tYhOJW203KvkWh2VOWmDiqMNYJxPVRjV
QWGBonwdfYrjIVZjJ1IKH6E9dQhFjrStGRFmLZE4Smd64GnU9LyKNh+JLo7zPDANuauQi78alYeJ
DIoAeiw661WcWBQGzvAaqaEbA8JZytj+oXe9y0zpVI6fSCMNhlc+f84BuhgfClN2EeBht2865Vhr
clP+KtUiT5tYQgUuL/qp0yTPYzsCeVjjSwDRqW7BF1scD2vz+GSwCl6PZvca9mpGi4lycNwmpqJX
Klz71UfCozyF+/gTbkCVq124r9FvUcHI6+iuF33pd+tNGwPYwNS/ec8K+LDKxgpwmQvyDzmaXKgv
2Vo1giKHo4C+PSAH7cuOBg3DZArQn64JogCHlM8pvZyGWyEsBa2nlAb1Pxev30UWVsbstZONTGiw
fd/KPIPykLW01U+ID6Ou2zU58IOZZXR9hTuxYQ+6m3vNWYcv/4WaTq4KDgsNwHN3CYxSKHj6hYqD
UvoszyKKNwwYI3O0fLWKt6iF0QvptECMzDG4Bs7TIb16RxPK4VYZFyg/opZFQLMMfVd95O2lVjgx
G3XiMA7ZflABFJFm+hbFzRtS5h4YGnyyJ/vnu1kgeFBqj/9sEBujDt1b03CHBgJpsnLONOXRv/D+
hn/CIbuz+CQnyl0xBArz1ryagCzEYHiq0jhw3TuKUtHJCZ5WJ9GmUXTO9uz35nCCTjdm05M9R53P
YMFAfDW+0G6MiILSWB1HU5Z2xpGZWmAA12pvKoEDL3UZaMSmjwbFNuN0VD2k+WmM30nZ7GmWBA7v
Dg+rKRlexlP0M3c1mFHEjfT5zSJCvMtwUUpXQ12rP7RPkr9FsrCc2GMa+xrv5pQCkjvRep6Np2gH
MgzXNwkE4U9tigA8jFsAZFL6KEQQQ7CQEJAq9uP5EIIlp3WhNthRsEfBHYejaFKAFUR7/3njtl/e
0epJlJVRRYbKXLWbYjOEP7oHZ1RW1lKUp2sGLsWSkNyEKI46TXI9SDxgQfCNT2uKjlFz8mIkzKWa
bb0m+AD5aF8+cI+n0fMpe0x8u1RsddhC8EcaAcunNJnBdFfzHN8mQjcYoI/jfzr8pue7jTMQXzqW
K8SQmTzX+vQN6lh+0fEFoMAJZvLJ+lvAa26uDefxRf2rASBqLvSsUfzxpbHBXELEVRuKbITZmlka
WRKddM4fDr8BMYLt4BUR/G7IAivU+VBFedMzMSdtln55PcYBjEPEQl01t2IPmy9Y+jF9wMFLvAnv
U2e1qE4cyjRpcKZUp6ynNzr3DnTbiQkVPfW1ovheVZ6UMmf9vKURsN/b9rR9fuVgD7xUHroRrbFK
TucZKKiHRWFjAF6u7DpV74t72wpor7hthitpYL5bncO6+mBd2G+7QaIen9N0estRkVjrgUn+6GmK
tFkoh7Dxy3Ye7VlVu+t25ayclug2Hc+7GzBVRn4OqqtYNWlWBhBWvNO8/W2Aw7Gmxe65XLDOcAIy
C0l2PeACx/9PJZy7zAdXb0XaFT4y1LNbB73zR/20w/fpI84UTHhi9L1wPWmgtEKby8aPRCVHBTu4
8BH2smwgkpCVGfCInqz+HRPGOcG8JWKrzEqysa5VHHGze5Cyk1bEV0Q8v3l/Ry/X4hJuHECDyXJ7
i6gAEBl28b+Xfy1E7jffqezwRNJofsdoUiBSf9UAQs83vBikCyk0zSYQ9b/RugfeBGPStO5KAZj9
h5Vng7vBLe0CNlEKWRCwZ1ZB8td4BlanoG8z+CEVbOPVbrAKfIMT0ONaLEGMLvX6Lw9as31c5bmz
3NJlyq3u0/aCgNXnBYcou7MhEwnB2oUImDutNTuR9OOIfe+vzumKNmOYyc+CIHBkqVKufKGgaiyP
ONRHPXswNYAJOTPhRBt0Z7oBbHEE7hirRdACgy3RKG2ArIxvrC6+aKg2ONwHIAt3KSFzTfdwkwR/
f7a5joFBAvMwu24C/2GnSflSoNdppbV92coexfSqOn61AmgEtvxB5j5PE/dL/M592E7RGIeGXHtB
7iBRtgvCDxd8yusShMqWLfZ4PR3hmjsFMPerbQH+gYNjllGJ9yFj/O3FyFFUBxY9yx8VsHLRh5l8
LwCAwDndjGA+qmKxPMxPAHJOT1ulmuGyWsrB1v/FRGNk4FxpeJEF55ZD2zc2hWgqjmzI6Bb7DRSF
e7NGwTcc/mavaX9GYZCguu21gzcybnX24HbwlF1i0WoBFaW2kfhmJcnNhQAANE37Zh9YwFmXuzir
MjC9F+1BTxooIBBqxggs+SbV1dsoPBZgTU+WSRnUSgc1S2Ty/M7FGiPghUrr7TY1UGhVxdy5RuVx
ZLEOw9+mAZOkQQww++nQ1vd20RFceVSX4W4YWgTZHCAyxk7V9TT8W0w9bHTZAuOml3DA5NxrwRjM
L74f55540uf4DUlmEQ7dtuuFdLx04gSkxk3azjLDHutPO5SVgW37tjwEA5Qnztrvv1wfg/C8p3k+
FcFT92rJB+8KQUrq4sRbzPnEd1yX0wgjinlbwIvuWYbR/9UYbQ23lbD1CRJjFSPNUwwD6ndYOvFk
li5rSC07wGSwq7ln7IdI0vHNZd9oiF3lbQ5ErSUI9E7Hv5N2j+E8TTNuE5g0AiRKoGbakEBCd14O
qvPV3s96UeF+GI+u8QX1xvjLhGOVcCWCrlnSFyvQpgO9YG3vskjVeGhoEC0eyaUR5kuq7tFpXLFM
YRp15OAl+c1VouURqsg5+28j5f8OlKPU28xUxXRSM3kdfTNSYpZka+Rlowj6o4jCWltbeJic29eN
bKSObtynTOUkaQpq5HwPTEldG7AeTHpqbmypovYnOPQosdEUVeFupJCEEKMhCidnUSNsfh38Uft+
H2cOFv8ZqeFabqzhvupzxQlPIn7tpCoqDfM/vTPphIzilqTuj9HqD0EZPlY8YJFWOV3oxZve2/ZQ
4XQKqIunoKEDGLGido5Woap79HIT5pWEJx1LTQzTYGlAATPyZxC4XIiBLvkX12F34zeTHuVCcYig
HqfT2wy3ivwBte7sgrybWBrG/Aj+wbOfh0mABLofkLUa9SWXdY2mDDvJsAwpbV+h0eRKa++2iSt/
ib7JmjxTu70HYELtuLzoYt8F380z6UWWxjFxh0P9yCNzluqHz2hYeJ3sO8P16f0kbOOcC6U4D/uF
jUCwfDRD0V4uEZRU8I8guslXJSSvYAYuTHqUVQ6LXruOcKZGGdy6AQ37MAkE66ASYPHDFi9/+R9/
8OTAE/1s+UsJuTir7Gx52tDBJ7nVWe6vIZhdcPGGFZs+tRkf3WkJ3dr8aXBLUjwSyC1tB/71oey5
qa/nXvRPsHB32qabSSDTLL1xusr+Gi1neoD/XVV0GzzjlYMtjVkjaSwQPgh6tTqSDLfMyeQLSmSR
v3SwOCkr8nuoXxvpfn6CtV5S2ABdU5iR2XEuZKj+8strkrJzxfH/3oH2EDyDikF8gVnIcWAenPiI
Fg3SXBxX6P0GZ20T0dMSI4hSOwBvtYlnKetGauw15CJ/Vbt9anVUQK5RHpGW1FBEpaSed+UwNwEl
r3TBVLlFBHfuVO2yBkear1GJo/m6fQ4C0w8CGrBpQP5dUTGCZJdfgAzs7IW515rOfEMo0TXMip0q
CZbum/Qc31BEtl//uEEXa0F17y8k/nh+QuMAmD75R/qkiiiEyVy30UxyyB2Y/MN4zKoVdCiOMDWe
oV+YZinEiWCO8PhE8fZhPMWaY5D/+oNdfoFm5cvBgiY0gARv6fD03G60dmGAbG9ZCcuHGvTaYjLv
Okb/bBnDzci/DfvZgpqtHxE8F8mOCneIFzXk9CLrNoP5kLbaiRLj3bWz/IIq1FCSs7elX36yXkhD
FIYUAc1j8QgCfI/mt5F0BtR+M1sFHN5ChYl/gQ7jcS/6+9ZcPp0TRyuTUNL3hkw3Og48+svaLDRI
Iy4e0Tc6Bdi15IpS6AF/ah3DTQ6sz2gkeFHJIed9GrTlnIOO6eu5bUv7P7ysWSAFxtqLLoFVIMrn
yExXRPnG9hz6mzAeEAstL6vy6gpiQESt1IGyUiEc2AV3+5kGZse9NXXIu30lzZJ2LruhDbJCRodS
xvAV6ukvw2sA5iUx8Ud3hbtQPhshlquUuK1NJZgBc9pwtNfGFWrlXUUvMQgxLO9MEgBTSiNMZp8h
JI2GrHszCjTE5zLXgumzA+E+Udw86/2N3QijsXE21i4Fmx9BphkNT8VsZJOzet797+FrQj6mK/IF
Z/Evs4Ijn4MOimyx8VkcFHhSOlNhxtJKDBoNS3/lWJtWZ6LANKiH1A/W+/IijZIku7wMJn5ioBeq
5AgZQZCQOuOp5lFFPG08GjKxg9o5cYxjtpwDXQDCuuJ488s+/kvQGGZA/fvy6XgAR6Jma0vxI2k8
6KtN/QgtyonfjSxLTuJDmk3aCZp39rinPTb/UVbo/Ks4u2PmRcn1FSXB7pX3ep34RVdnVQswOrRk
NvcmU6YVr4InAqSM2toMg40HyvCz+1Ba+mAPlgjug5t/tf1M65c28pa78DCrTWfjSDoJphdHtMDR
GGeYttKqmmEGNpDDUMi5C6tZVjemCe6o9xArvYUzlkC6em5bU130apN/03BIP9Y665GnitT5ftpt
NpNgSMdb++4n8aRZLB6jMIMpJIqb9eZq3lZQ9gS3xEdcAlUkN8dSBQ2Kx692nk4UYjaFAObCebKr
3AaF+FqrKm8E5nuw2r8PC7tjtG9SnMulX+oRP2SHT7oyjsoTnzaPpm9JlZqWLEs6xuasoRTNCB03
9Dl67cGFXuoIRKAQnU3gCaxSmVdRM06N3ymZyLCcdKzx0ey5ZtMuKqqzN5nYUMNwDDLu3QI/GznS
Vnlot2HtUe840dFQnRzyb/QUmy/oMj1KB7jYOE4l7ZU41q9LFmPk4prxcKfGFuBlv8WRNTjJrR+B
JCrcfVcXnz/wuJ0XCTcDnE278CqU/iYYRz6fkdXmUqEbBzB/n//Xzx2flSCXnziml8KWVjhuPycU
cc7cxMOIcQ8jhu03Q0VvgyDIEwnP5DorAc9KoqiaTILWv5TlCFTVj/ltdY/4UU/bOnT8CPUr5tLu
KmI3c7bu6wkCRMsID+B8MeOj7aD1q9w+e5O2tFfjyn057LVj0u6twij6S5ILVCW2y++boQ9NUoiE
B3lz53Ysm6eZeUnpWNNVIOAhWPFHiLckEwH20hKL7fsLaaY2KxzGOBHmjN94uWanq0VjmpmTuP+S
1T4nwBkSJPmY9Dk3V9YRNAlRawjQlV7WUB7+4cUy0dS+YPrwOvav8Vv6QNvHsRYrAeaKI3FkxG1B
47Z4JdjuhWaHTbxKts5MvVjdrQtETNpx9EXiEDujM8w8Izmp2QDmXo2DE5ZVBA9SmGPKbKeefYGQ
DFY22SHIZ4ngQQWehtSyPJfTN6pr1kHP0YYa1YmSFi7b03uRyPKSP91zhi/63ORxLLQhBAbP6GHN
qxRl2l+ByIBQovjzhMB/Yy53GgRo4DOfLUB/ffdJ4dHaHY4QdcJtIr2ENYwB5B/yzAVO2lFOcG5K
VzT2La6VgnKuiYysVewf+S/Mem2E+vfrfjySZ2njdt3nFxU6atdIIcfsLvd2KsLMNy18DdJ8fhmx
g9g/hGN7JQz+SlJZZtypbIjx46al4JyQ6a3Yp5Ul+p9e0eeneRDFeGv3z/XInnAsqwaEGJMi+ZaX
zI1xRSxQQLkysb+oLLX4jzclBlViMkyQ7QI+ASahNPiSYXX+xNerXXIVY7PJlolxt14zoPG2X6q3
zx3js0lqWqSrpMGfd9XIk8dvGrZbWaSP2J8cabre3K21ca81dZ516vWaUjIYsEJSKv4RjisjLBtY
Tx56sMrwpwoMRWzw2AYHTG+rxcocKW2d5d8ctgIYONbjv14Vvs7QRwjrI5ffTyNtqZRQBF/VH/7q
/w6GNmLw4Zdf05hgr5iNRac8XWNrfW8SYAWbK18iDFX3JKXm28N7Ax9iK5m2HwKFjWiFZmhr4l4f
lE5HOsCAp3A3CtDDmr9y3VVJJmTV4FUzvDIOHMUQasTmrBCwhOZgoVg0prLzlQkWUicNx8mQyUIr
2gQnh/ZpiFUgH/tsHWy80LKH9ZAN8giL47D2fdgSCB17Gq1hdhxR0qXyUh+Wa3nTDPA/AqFlfGtN
lHdGc75TVjziVIxEm7+ulcLQBOS5eeM2E/GiOUZgc1sdGtlS3rX81mvYsHrD5piyr5EXkOdjHs/b
gp2vzVR/UcznEFTXYCagoNUMkjBb0XFNOGg7RNdexBg7htAxbknyQ5KfybpMx13GYO6AQFPjXqxx
miywxPhNL2qmURb09h3vj4sQ4j9+mL7ID5Ghxs1T/vaHKqzEmETkxTiQdRyldlcAxdAprZEiS9pA
0e9WvP2qAhI0tczQihzBgLNuXgy0CncH9oFlVhf915W46zx0cKYXbuBWO3Zy8S68+HcLVGNlQNLq
aUaL3UT9tbKED0v7NWQ40tXz87fHP3sfe867/KgPucZtLxKYK7nuu9Iym5/G1F8QC5y0lRQWTZDl
18JHqK1BxTiRZxibESiB63RWFtsBO9t/TywIGuBAEVLwIYhafr6SnAsMgmLWouq9CIP+6wwysPCb
OcZQa5liOEaybfc9jAP7EF76MbwuPNPnK0MFolTCXmWulOVB+K7qSuOEngu22s51fgzrFrFai5U0
C3+GrMZNckpJXHsq6BmDrPruUyRMNUtYYaDh47/4snG9MR+H0yBusOVvoyX0dc9zabKrX6c41FFJ
jFlA7UoxPk0HXXBW9rf8ab+3ds3Egs17Ea/6fSGaimpxZfJh3P2+jI3Wtkslp2T8D9n9/zx/vN/Z
+beCHTTxQAkkE1zTlqzTwQiHBCV1t70t/td9FlnspW2HKpUYL0uGHw5ZcyaOi1r4ZBxBidNC6acr
7wMwYUTbcczZZBnseFR3pT6XTbHc6gF4Ib9szH07QfHdf4MaBlzR/hnDjDXRrd55OcxhIWK1d466
L+x21IOntCauJ3NDjyVu21altgNU1FulmB4h27E7hQUejYjm1UEvgfABFkheRX7NobgTyeZw5xh6
Yo0GLbiCo/hDpB5Y4LWXuiOQfMK+tR4Wp7BN8s5nEernLW1ZKpPbCCpUpbXJLXkEQM4PbSsGbyDY
csUTF1ypZ+NjeWZuO37hkgaGFqsO8awTy1cqqOK7cp7470kD4z4rZ3b9FesGjknZZQmmPvwkT6yC
4JSxHwfwVcSHq1y1yGU1YG/n9m2vh3aCAIon+9NYKD1l/cAstnge7FM113wIyNnWaiE44TojVaFI
7bK5OEUESuJfbeNPP3u0oR5DRl1IXP28YEfHh0C8uVPD4Rx8/A0N6sn8hdJMa7fBRovw7g0afUKA
h23DpQKUsfdyFUipxvAmeiWJ6h4+w2fbcHm3MBvhNgpEPfaIezm0dvAQXzGYFiBGBTW1E9HUdz9U
grmwd0whRwFlIYFyT373w70NnaetCPXBWPAH4H0WBHWiX5Fro1zVgvE24X2BVC2IW7Y2nbATcSBT
TFb1Dl2vn9O7K/di5nLMOn+3s3aDvA9qd8u974JB5fk4OulMhUG1KcjR8s4cUCcHJd0F5JcUsk0J
2pdILAppyomN0c3plemJjIB+yBfUzopOszxDbAHLGkH6Si1qaZPU2eM3nbAuX3GsaMktlf54kNL4
ZUy7FFqDZ7WVG3p+1ob4f1R7GV9kP4f7d25PUUPFNRrplF5kioInYFhU70TVvd8/UocRujs+N73b
sC06qAVYrWbY1gAZNiHI4NM1ATunRIsv27WVqxaRciTlzpQe1wzPTZ/DlnwpSQ9pjuzaWmTU9DIG
Vf9qPb1cS+c4ABQlOzgAz9Gd4EqmKqOCX2eNXXPQpZUjqszzcZ+wLVIcMZGUDFC+7A0OPulaPv5v
aVr3NHR/3QgiS5Y1daa8JzaQNTftIJTD4Y9IOtZZkaEh8cGwq0WWGpiGddyuiUP0FEfSTXwBoMIL
Ry5mu0VVdG1JlZTjZd/uNGRUVcTHF5HGPDW0ud8tjaoMBlpelilmyO1pjFadA0pDWrO1+Pg0Y0Bi
M36GuJmPfVQGzL8ZkyBHnT8d05e5H/5yZ6BdRvtxy3RTltNw8S9RY5DeNxe3VLHWcnu+4O+WWIe8
LUeAR5gbs61WB3+RwbFBqvAJd/+ruf2YeF/sj7o32ezuV1/qfKwL0KFdPkojjFK115kqrqRUgVR8
6NWaj4Eca4Tdx8Pm1tlqT9RX44MYmcsa/daD9UsSS6+kpsvpAtS1sOCR+33aKAr4oFVf7f1iaIy8
yLx/ofxK25GvR8ZkT123JpvteU/SVpMd6sxo95FfZKPJUTE4TRj/vjP0iiAXY1myqE4e6/5BQzqI
ISJqwG862VgiLvO6AiDVQqkkSP/LHGYG63ArYJS1wDCKkBrEV33xtP1q6ozODYPYux0kqWNNfb+y
L/uFfF8PUtiD+O+r3V1oGbWE+JYewbkDWFdnHE8Vw95tuxuH7XrrFfzp0DcSekmy8X/F8yRNeXXd
5D03pJctwQGdLJWbgVfCzr/rNckRw4DIjNjKC5L66hmsBrCu0Q5xoSQp6vpO5AMCd9RaR5+NJ034
rr+QrrrLQ9J4GxtCTEeov2RfjD3o5NO0Yv9OSZnU13hVW+/awNLm0VdZXkbDlufOak2UbL76cVFw
jsttM7/+BwWNirj7mkGITe6YdhWnKpA8E2NBM3qWUWIrtiEELhELJOBMDpF01QDLP85jOm+RXxZz
y7Us/ntG8o4zGn/qCz/KptOr52Bt695xaeLeDp06uZuDaO8XjSNrDHzOscy8lIRkKiBek2LyO42O
4nHrc2zPUiPjDNXlXrHnFCPQMwHjxnfQvIiyW3dM7gkSt4Jj1HkbMLzO2Q5dpgkJGwl7sbjuLW1K
Fbkngx4WJA3ZXndZkN+cc+lrqoGpJgI9VrWPV3geho/BhpfBfBVE7pGfxvjrlfhMCO0wmjKtEOvp
CFHvdeBl5FGZfe90m8MXDsWxto0fJ3YU5W8FqlKvpvpFsVk5UvAFXbCeBrSSP5yb7MYED3JiyhLV
/1eFXsaIots/k+s4vaqP4cMKyu85l+k6GuasAaFH9MF+c2fvx/t7Z7YCBqEtqQzmpR+T9SzNhCRr
KGQiaLMd6e1KiyVdfccaD5FdzuYFYYoozqUhiD+ntKXomBpsDGHXpLebHR8NPSfv6ufv6Cey2ysm
SqBxyo/MdvvNERQXAlbwVDtygSxLj4huirSsLCr1seNCGc1xezallobLfEinxSo9mG+Hbdy284u2
fYB4Q/7NFqqzqJfwGFC70hw9LcgVmF1UP9yxUzkTHFV3qrmbXpdoMcDEJlUKuq1r5fT0UQa9RqQu
10DIYuQlHb1G8umM53x4V5beYvQKxKKYlxYqLXq3dKb72e2/BGIYo9UyZ+xl0VnmG6IHsLWtcRG9
a3195RqqPWVl7HTFv8PQc7X0OzREAHbLIAbOpYy51xtAlRTlobjNpKuWtSets57uQ3/u7thD+cvq
06KTy01IB+7jjwhyxZ7QMEKfzIMFwawQKGWvJitfz1rtJuWLkyOMs33iMpn7humxSsuLucouqemr
uoKFB7axNVSFEBJ2I14btxbrS6dkBscAIXKXJHHxmP/BBA62O1b8UcLMeZFT5aGBb1uBVa6sScSM
0uddSlrKTVFhPEvTsLQQ/dimZPtMODe95zOjZm5JUhq7jFas/AnD59Pw0q4wTgeXpHyY0VOHS5rn
7mqJtNGuAXlc7cN5JmBwG/cPjIg99sAvodcIXRTia/b6MCVFZ0yVW998frw7HHqFrjUdwq7H1Dkl
4eGGbPwhuFhgCAlu1Mrx5j6mbRLD2ngg/B4kPaG+bK3P8T3PxeN3w5taC9jcD/1Oryrw33IPP/Cn
iXANuIWZA7Buo2HWbDgHWd1d78FnbaXsZEaBbQvzno3mhAQJeL9COXJz3jQqgN2U/Ujb+gKTEvY/
hW2MTXFQ1TPfnTy93wRoyNoGwxl28lkZK43xL8vsYncaqKurEZRENNC/ck+zgRSfeYNrcreNVHdz
bl0qc6jZA0h8gqsUCwLVNNK7Us/OOSMD1itz1ea7audOz3J/B8avysQWCc9BJ8OBBhoy7tuaqHQJ
42O4FLNZ6NfudaEgBNntMmTiNuFWvIqWkM7U1LRMSrWaCMfMIQ8w3QFmWx1OXJY8hN1OYBet5jEA
wOCknGkgkybswavpeJU/dBI53CowZ31lzIsq2sL2Pel9hIftmnSXlv45VB1Ap0HIWEbG4Dm9TR72
ZESkXYtac75iqcQoiLEaHNfOwbw+UNnYTFKw7/1g/qWC5jLAPEprJH9NJ/NCBSZbsfPokKm0E5JF
561dwVk+dZqcOJBjEyXECYpZ5F9vp8BFn/UuAhDZHm2bCozHpTr4rG3jB5Yz/nzSlI5TDRtMrKiD
Q5XBxTT7b3rQpyIdTy0QuH+8uZJkJQrC7tnqiyWEskyga93YhG8KOOlTClxxT4hKkFi1zr8IEhNd
iTFzs6ri+g+Z45WBxXYGbWlE1NTbWlAEWtQ308hla4DvnTEOQ5iEBvtbNoZJy7hxTExmWLQT2t0o
mIp8VFHShVlBRelMt4LBrGjWElVLaFkiUF6u2ZixBnDyeUI/pseEUckCVDw3NNE27ikkDwuw1baj
GwmsKoYbEtEMRsT3f6SOtp/yP+eRCaEviBPQ/gkXTJAoHNvRDF+iWqab4ScHjb2adXQYXhjb7y2I
ScbwH2jyFBMHzW2U9JGARzehjpNgG2+ygmKEJ3hQvahP8bQgzjQMu/qdgCt+YXtE5XrtgDA4X2wr
jyg+QlE6QCMI0k0PoDVmsFEq9vuYh/fDJul93e1VMDKzMpS9IK+tz9zi0MX5HXJ/T2yRicjcpAct
I1sFpKYBHOzIcWfpY4FI70hVSZ8uSea7R+AoJqMxI8VQdvnNQ2vgq0HqigiIklVRVqKpJ3Jn/VPt
5MlgPLAN+lgA+Ouun3Ik/w53LhiXIxc6xKRV7QYWRTAW6JCXY1Ma2RL56FgkDexIfCs75qr9dHhC
RwLq16GFfbOw1AqNAIs8q2Wjcg8h5DP/mFv5htAD/kcHA56SEhojAnTqf8dL+axf4K3A6xNqIRye
1mNLSWAk9Mtxp4OluiIPBc4txJ3Zq9Xlv2ycs1GIetDsXJOFg4BVOjQU3UcpU+AXeWaZXpOMRx2f
ki+toFn5p/OPglVUneGjIeMwQEX8WZnHV2Uoz64RweFbnGI5krSzajXKNCuhaBXPCGPtkR3QvIdU
t69w4psD2uhhIjwbCS5bU2nt5jLmqwdUu0MSL/dvyzXZvjhs5yJoy/DqwP1AHpyyAjGg2lgkOOQt
9LIQITWbSnAL0h8q1/0zECHi16Kj3z4aaeyuEArEHKYn9J+M0i5QJQA8LlWoJMgLBS37CuAbHfpC
9bGYFzu2jFcMq7fZLQUGEIw5iZc9R+x+MIpWlogfg7Js0gY9FepHl+Y3xatDIrrL5PMGShSZKOK3
yzDBPjLaWvN2Zp+ASrOeQDrWgFcmv7QEwotMrYcwmkSdY3Xjn/SndgmLGHr7g+UsTdtcG2ioqpth
BXYYZw+Xx/gWJBLdFyGIJ44HY6M1nMgT/u91S3hMWZNp1ti9NdIpAiqy+6GxCVPuQtEAxSjN7Oke
ILE23H5QQiybyckvuLngZITtty5LX+xYAi6OmV+39bVoAL3emqGEmDFsQunfmwxwPhKTAUnubGaQ
jcxW+heRn4bRhVjh8lS6gZUa1uiUKCG0RdrNCv52kMcCc3XKB24v/MiWGEZi+QHdnbdjWzQxLa+5
+9lVBaPydmNUmJaEUS3VUtOA3V+naoP2a5hg6t+8uD+1AI6WpjhOnPMnwsDfr7Ej7Q2IZBw7Q3sY
CCyIoR7KjyYC/PCPhWKjY+qNUTIJZyLeS2uFKDeVKTuEq9waoWoN0J6tM1/mhTcRcgB2u0UNI4Od
Q4g+LHSuv9EaGHJKdw1ANdGICvf4JZo0iIqDgxGJD8gNdqDCHVD7WqKTgv5LzXqqd50QYsuOvO26
I9asH3hYJe0eLHSVgY/csC81bmKguQDPuWPhILEhKO/NbICmIbnOSESkFOnTZqXRkXI3iegdrTs8
UqgC96kjAe4AQzOphJFS5FQJBmtAR9CYOaVLb9d5md0dNrHF/CTu5d4dPwx+z8n+KC+qWwIgvxYL
FnqEb2V/9LDVs0CWryAT+qGRgjJoyK0le2P45ZunBXEja2nUiZcV6msAFm9eQ2twzeQx5WUzFRyo
O/8QHMMXx4nl7UegreP4TInFnu7aFEnObjhCIvTB/hIqXHyvE4D+u0aTuGB+jwASez9MTFucHhXa
opccJN/E1bM7ePKIKLwkwvEq0yuOoiXxoJ7og+OgM8qMPefyVbb3zwM34z1YEWDGqnHncW8gZ1MJ
GvVSWVZC6LlnN2LoT47kF7MF9ML1uMODuPKcvq1UdoWJe3uDTmt7gB3+ORzOyYX0dJelSwTNKnXg
QYzV+P8oAiqP5TaJ4AB46liheZ8tO0mAR+/Xnlri1WSDimQJ/t2wrP8/X4r8xC3lHlPofgZcNKqi
SZoFq573eyPR4moiyJPwNDUSmf8G5MRCZASN6klc7nsi5/JEG3BUQHAlh5NhbEb2eHjAzZWHQcfS
03hj3iepRInsphIkjl4Lj2CDtXa4vKX3olTheyG/KEuSJTcR6W6rrVT+bfdokw81I+sYVQPer8VW
S/oAcfEFxg5Ggsjiq7iKiOOLszi21N8u0FFlqU0sSBcIb2c09XpSqqbBCdhSsfImvTvTXLd/wqjW
sE0Oa3oU9x+mD9fKw8DZiOkdyD/gs/0QhqP+K/Wqzgjj0kI5LQHdq6Gxy4j6t2TE8Map3V8K7W0n
RNnfu9FW6yg0zvGZ8O1XKq83zIQ001RSn+uM58kfhJ6jjeZ0Da4ZYLU2bIqvlfb9IinzSS90VqNT
bUiwJmfbk1w9ZNjl03732RqVueTWO58Z5J7ve3qbmExik4k30L6PSrbjEJ7JHEdwFd0qjog3WtSi
MGbVZpEo3zA2JWDvwEr+1D4UrsK9nRQTG08CUV5knqoChPeQ7BScgSLTAEVYUCOgQZpXmkjXvtSp
kJ/B/MuX+bk8wXGnmF5PE8Cjf9zQxOu6TI9GgMkt6uX549Bqz/iCw9Lwdc8wpSZGfTeSPPGLoZSG
AmHH+QDSGkSb6EgIQaFHPGYUOBPjEosmk4FEbIzM0iuUWXwrPdhk84UcUUgJ/ZCjdwP8wb2y8emx
OpA+zuZEDtPTWchOISyxCFLueGMeEzJ/BEdLj0z5RsZA/XbDL2aFV+SS6KOiyeuKC4Gz5DVGqvmb
6FI6mR0XaIb80VXC/KxOkBIKltf2/dUsAjNvLkXSraW30gN7OaopEjgQ6WWkBRXPDeyqJbqIm/X6
CaoODgCCl9bMW+nyE9csfCJTYliOQzYlC5FW8zlakHTEn9iL2U+lJBZ+yE0IQ/1Lqk0TMkmlp9S3
NE4LSWqwdpxFZulIDU6ovxKOsVB9yFSYYix4p4BGsLSFApPEXqCSbxtsboWXXDZuWIQwx0B6l2nA
wkqJSBWlKRljpUu459UxICUOGiGTLgR6uThL3W7ovO9nBYMmqK9hRTTrj+4RewRWQ0A6WdhVN4I5
7Pa6vtb3x6pyZNQHoSpk2R7HubbVieDjY8cEIaXqll2u7Uxn5i5VTXo5h7QdDohc29NLYbTbzyOW
lnnV5CQNQp3gg6or6OzolZ5uV12qRwybdI3kWKSGOhFK5z7maL6EQgcvrzE7cTnPRzKd+mXHHLbN
zue1IHGqfrpY6eU7la3tlfKs/Vv8slann3kaMe9s8psE0Fddj9XqRpVgSx97Cyerrv1nws+h1ic0
NIOj2VCDjwX+uK/tYPIbNh5sbTKGGHKyMD/9gp6X7z7BkZ4T4PtLZi12nk+Z3/HyAxXi/PsIwOKv
aT4/K78Ow/iJZE6/3Mz5jaTDvDYm/ubm2r7YCHbw6CvI4RmcnfoU7tXBrNNzZ3QvcRtZrgW+pG3g
n4+ir6Z0O8LhJteS1bnYhl5RPL1hEu4Em/Ms3sbhuDB1H4OptVB7yUUAsEcuiRXfCgj1lpWd6Gch
PthP1pX1e039Kb+ThZ9E4bjjl3Ebs82mRp+vt64cijjzZ01eF9iMexTOMUbQn0NXqIxb2Axw/p/j
+rI0m5Z/rUXzRCt3acKAu4WgytL0m7ivER3vNXFksL95KiVRdD+zg66aaBHYjtF57ws4En8W0bji
aNaGvGiA597bW66T9/6oXGFZx5MTfYrU2iqv33TlrM+K9Mo5k9HvBfww2u0ztkIsUggtVxgDIvRm
9h/fQgSOu4S0nicbBwmH359Sz8oOw1e6MascYmSZheLyH7KySvMMNgB2r8V5QsTUFw/Vt+esquWo
nOAZHVH4fANaJ+HK/XPLAz5ZTYvanvvaCuQEtX83BIBP8HaOjOwMQIomaOFXBkOtML4DbiTWlAwz
jLVIX+xDaIAl3OM+4xHOXQbLqNluTwArd/cgwGbYXZ4BOIrtxJMSuDbunmVtaFBZoIBT88dQFdy8
Kdf4XNHGXi6CWLnnApnwM5M0ag17hGSAykbm9eVBUiWwgYfnwoYx9O8NhutA9vXV5dtJf4Zw5kU+
YyEsyBudX70Qwl9WuCo3sUeu96lzsz84QDrbPwTH5NZsT+L3rWy1WL5ZsUOMNZ577DHl4gDS45Lu
v/5zLzmxR1VdYkmNpL6KaG3oZjfRS441NVdqkdbgPPfgO4dsKuoOLPkWmpCYqohVHEB+mQm4IPAc
RxiftYco0BmtMTUam5AGFh/WtQl4gtlSkZBm3Peb+S1yZzgNFhbIOUxRsAgERZbyIWSavfFrX0wr
KgjkqHnaOBNZsqKd2n/5EawJIMEUwJJsxCIabAZ6NKsJbhIn7dp82vqln+UFpIxCvQYH9Jh1E4T3
JW2FHLo8W+fZloS4IZ2Irqfu+tflOWQWxUhtV/owtvRhwGoyRmg1ZTzHCOWz+0ynuE8/4uWDkoBz
jmkPUG+ATLaMqp/xeEKIoIWvsZpdWkgDmW7xRTdpPGc19GNxLntFbw7SkFbWCjhQU/Nm47q+2pxw
0Sak2lE+9VFE6bHnQ1FRBoF4rQqud0EsgkN150w/8aMQueaDrMqzFae9hmq0gQvoCvspKCdlC+Au
8voEy2hQvgV6GWa45gD6Lsr8p0n/RkhY6p9MidnFAmq/ak35Xd5p32d1zktAVpz3k9chQfaBx45y
KbC1yaKU3SJAsMA91YKsO2fB8dZFa3lwCdVqkjIQB2jKwTVc4aw6uMW8YQT4M4JaknG1dOlvEE0F
zAJKxGihZYNFl4UU9nGF+vDoilEyahz+8aotcjftN9ZBg30FrwyQ0bnftx1FZSl3Yqa3MYdTY1LL
apC57wvbTbS8SCqr9r+k2fAQZiFmm/1pk7V/dcPnTuZ8UdgvgayL4hbFD72eBmWbwTG9JyXggNkF
EpfLohZI/9jHtN+4Nr2gaKYObLDXfZGH4qaVzn0Jb/IxN+WtcoagXEM/7YYjSCkzSHRnlq7vM01w
9wjMqBiPxvBDqKvNH5oH547FObnMNLpRrRp/46nckaRIrB5fS2EiSQTwKTF7BQ4jKFu7Gg2MujaS
Ydwfdeyo8sv0mTq6yvIvNR/AGOHZC2lRJ23+C3BL4nvLDQhtwJfTgysPDSeapDb/ExZlOtETCudM
zF76N8Rxx31QYDYeMI6WxD68prKEc/SzWuZrdz1v03Q4/QZFz40AIKydKIw5/+wq20z7qDzO/fTi
qS83n9vSvb9npIx9+h2PNC5hK9P2ZLlVlayqgzbq5xQwm1yUP9ELkAtuHwrUk9N9ibgb5V4HVArr
rwbtxRtxy9HV3lu12MA/S1s82siqS1HzyTEqy4JnjCbSSTnz0wM2wFU8fXxRLHFc7qL6vkXRhQzf
jVUr/jvIBuPfrpHvbOU8NRXEa3JpiIu5d13dZTsB5hSy6Ir+WHY1KNq1CMi/BVnBiTQ3tqW+NVQ5
VW8smGFs0IQGlSLkZrppVpSulSzx2w6xTkO0Tr/DX/OMD5uwKrIgJhb47RTjw5OR3FGxV32vCXoq
hPSR9/rllLgi9P78y6qLZ9mLwZwkJBD6+CpOOkjN0166S5LAbEzejjSQsa/XEqHgcllkahYH0/a9
PqyUh3j8eczowv5E2LXRI1XfuPUhtqWpUsaZ1wK0S6tsB/ppbgJ/P1R2olK2rpVOyUUwyR6AYITY
ssk0YS+xCpP09dYckFGzVXq7Gq0HB+vGyiCsjzVTOdc3JOgSB8xkq7wNuu0KqjFX3Db3kxpgrpkt
YhjsC9+qZVxbz5eM4/Ud3U3meFvEtfu5JRVapuo2ptywAlvHzvs8xj08P0vK/SrsL9wy+ijHFTsv
ncpqe8Ml1yoERulmjS5bu/ZrC6o26o8dcWOwV9fjcbDzz3GFu3VGFV7L4uEdO7wOppse/ny8DxeK
ocDE6B99ylEJUHZbF65g6rRTQMB9OYGXoPJYI1P6Z2DoAIvfDm9TphXay/TsiW4v3uc9qVCtl2il
4sdn4BcBZ0+fD47+UNqiQmdipP5n59y2D1gNPErArijEGf+oDw+dm3EmY6vTHFD5e3PpAx1WwBN4
mIJ4+k+q9RJvWfGZMYX+/noMIOQCFfVWPUpnICNHuxWZCdgkD31gullhqSzV19Bpo9qqMnQGR3UF
TMT/UyOylpocP2+z5ll1w4zF8Tj1SbB8FGqtBb4lQKsiaFABupbRvbW6U3wNFzcZL54erLTC29J/
2T4tFTk2k5n2NST20ql+DEjyQHgg3RAlYhUdc1VZo++9PQasG/I3mgoIfvHL16vaHsXC+qD1rjI8
gGq1RWI+knXa2txLRf2QL1OxYcrWYp0tGlgQP3oyaXMRj4EhtBu7GMGJxKWh3BH+IH07BMqc5eA6
rbxhWYHf85epQzJ5vXKJyYWVIsgN/FA1o+Y62MdYVuw9wSlz1x3ZDIf4RKjc99WhMudBoBtKgz64
EP1R/lmWifDiVC06jj8gCZCkgxVRvwEdY//5xeq2ZmZUt9Kuzi0upkCptp2+spzJAWkebG+Turf8
3ajvcOtjPxcHy8DL1H+lWgT3CuVc5s7zEDi5o7FFnKrjZApI+JVbAK+zWZ5tGfcy1VNRIwD4qm2h
zYcqz7gLbuvSYhmNNFnxXbdP0hvKK2GUn6iKNoKOh9h25gcDb/Xh0FwhP9F1UN79/T8BdzAgtXVo
ZEdDxaomV/YNZq76D5l36blVBet7TPVVz2XX6JPZoJi/Kq7tsrmCctfEKUEpiSW183oXoB0eriEu
IatJbMAqFnqIizQdBW+3lEJiG3XZZ439ojCiHrAW86k3Wn88JJBXvvkjhqp+DToCFqQYEefeGsd2
nwXqHAV6x3B8rZuzvlW8gPztH1l40SATacxh7vgukeJE+J77KsOXlv7jiF0IBokPuZL34R5LpM/K
hntBDLFuU+K6VHD2HR5+KVakk8WdCNm1QJSkqPu+KLbpmlUUW/PhdmbjdNorNTZKH0fA9IQQbekb
OnkTEocT8IYvzYa3JT0aXb28VwQO+0KYGLOb5KXWajYXwBLLUFseAt2Xf/vq0LGzcJQyYn/iQ7hd
6F323SgvKR0AS5XzbN/jIDyB8dRYOl+1XJW+vNzhQeUm7BS18nm2IcY0dPXgW1HkMcJAiIw311af
obAYHB7/fKIM04j4nbGdMuion4fDG8d9RppUZCEHOVVkOMF+xNKgrKoiepTgrMqMXRntsQp+zap7
GTSdPHNkcR46k9tWC6YX7Xu5gSQYtcFZioYCIi2bcExWEfk/wCpiZ87qLRDsbOGP+mRdW2ncTDXL
UhEc0mg24kao9PhOwFyoMOy8OfDZza53yxn/uzNx83wV3hJfNrXc1CVlXDUu+7WD1pls6K6maICM
dBqdwhGkhIUbePKrFa/pfZkt9OM4p9DJqrebLoyrrc+EIdwJ4+/8k+uYQC2lzqRiPOPmfDcZ4BOb
odGFk2nqwq5fp0Q/h3o1YMNOwLOTaJ1JlIZjbTt0NEaVtxgyicUFZiUdd88W5tbDS0KS90y1Tn3P
K9OWT433VfrZTQ0ISgxqqDw9MrLklMzNmb9G2+f5Guw7IvhZUJfrWR/RZSibInqqyOwGCHNUuSJv
dvpSIRJxxn3A0NMW16H/USzZHSHEA20c2Nf5+aC5iAdoawkVWI93r1nvsTZgoXA/8h9racxGMp5Z
e6D21/7zyvbyFCZzFdEkhj0fNyQYZelSC93T03VVUK8pse+TGMzuOWnzzPW5WKNe/V6PlHGj0+a5
vwZrySIHg9TeiOhcPr/XWzi1rJkbbyqJZRykHVEB1CrfOIyEMelIcV2d9KOHv0Jo/j+++ZoMr0up
VnTuT+qdgT6fqajPMgyeyzEaFsFVhpiwW1HDtQpQO5P1PsLPbBUBW6ZLzO+5LS8vQCrdFeKIukpL
BBeV7BMmU/3NdX+E3NFN3Q4RtDbMuYrxOY8qO+OuXQ6Rbnzlcb3cxcd7DqSFfUlOYCV8krtyMR+h
+Wfb5wcSSkshVXfactrW058k85F7atsjEebRx+GtBNus4RWW+wbvJ2mLGkbIbXI2vPhTSqcHrWMm
dupCCN/MVHk4lIJdNWYbRcCp5o5VvbvWh6SlgrKQgwdtPqvwb77CAf3/N1J39cYsfJ65xnQHjZ+r
em5yzIn6KA7KK+512cnO3FoDsFrsEu/tS8Gq+7pvcrVN8pi6ezPx6YqOmZq5sr1ivCkVZgO5ZGn5
JzPD3P2wGVaM9BwS6vyQlqvtxQCy3xhhbm7J31zKcU/EbKIdj+b39Se9/4n04tMp4ZtCZ74Jz+U1
OY4xbA1IfVo2RUyhQaT+c9P/q9O683Lu/b3BAQetnfN0ZC4p3wrqIC/mHsGeEA84/Szp16Txw94H
ET/ugHMvqcVLNdyw8cczBH0G/eYod2gDiuHHz70gkMed27BxomM6Ooz8VU0dT8LRQGhZVmd8inIK
3HgWYGvuyII7A8Pqq7cY0Lks/IMmO1Kj6VGHrKxxwTjIDlwKFjqmhGaJnihhwzymapPbMkM1Ss9R
6hyhK7cfVBigxBM0E5Lu6w4vDZY4M2Cb7jmE+5nOvd7pUYRD7xHWPS6+p0Hzsg2OgxMyC4VTf1md
Yu1PbXoMmvBgHU63tPEpTkZXOhr+bDvxQSknxt5Co6uT2X8Q796hP5D6MHloQHnZ+qt9XPP/A8k8
laMCQ4jBwd+Tz9bGpgmiIzOZ/AzASKrV4hTjJFWUTg6OhDFXhtmCjXVARqFaUjYWGUh098LCaTKW
7fp0Zdwypg5TW3V8ICf1KjafHjFDRG5zVjJ5+zXxBCktQmXPmbDcNGzcDSCfMoFaenWPo2KDiuYt
HBYJGHVrAQbV5aAr/Z8hHYw7Pr8qDgmkSiALpqz83kggCbLBTHvUegrbLzVDCd5cYSDx3pNgfFhL
tTygQuU6alZieWI3MaQyXnKke66gRu95mfXrYPMCdmMuE9F/TVxyt6LLm8v1tVfF+uW/vECJDF7k
SP9AGuk9KJJTajMp7QWpAc7cy4MAkx+k4U2aH+xJEfl0KNZGiz20BMWh0VK65AljQDt5RiTunBYN
syffiXlXqmO4mriRveXmo+dU7ksBVX6FL0W9VutNBXcTASZ/onnnD6DFEnDAkdgV+kKnkX9x8ctl
J8SGEiex1Ajr5MovZTLKm0Czdg17AnDsSxupKKdB7mwvELVSc/fnHZnaZyJ1fOTdse2md23DrMiv
3VYtFmNWAl2UhrS8Vqzkp3zqgS3GYRk+bFRZGjmtdD8j5R6b2fc0GCA0Fqz71wT5KNyC1ffW5rsz
gE2Kur3ckBOG0kCdqkd2IxIf5qHo6Vplfqf2svHch5FxtEEP1Stwvte/Vg8bBWqZJZDHXKUICyd0
0ViKylG5oFLNvf5eSFkMWfYL6/VH3HCJzQ6jQWzlf2/hAdPcv4grt4+iD9W5zk265D3QgL896M57
XwnfS+Oox/4IzBNv7rCHCwXDaRbkDcAb7fQuuLWSywyO04gaqmDIWQWvmJKT1NW779JMSSaY5Y2I
CQrk/wBqq3atcmMcDGzUNA3O0qGchsUfeOVC+9g5qMd3V4eKjkMHZxh4HH4LWkxRb6e2dKN8cxoJ
NgNMfROpd80pfJWLyBOSpT1gF3J0HiFHWbMu3i0itOYgndvlQiNvDNoJEV0qap4CpVK9wMHIGg1c
T1p/eGA0QkN47YuxeoN9mp5qnUQNgM/345CMXHNE/RpyNLa2VZmvb8w5DaNR8pbYJtEF45fpopyv
G+IPZ2CxV3A5TXhqxijv0Ia8knRR1E5VR0ljjUPugoOgD9n6CXXaOwimrV0wvVHQLXsG7cl8+jOZ
qmVAvXdeemNg2wGerVDjim62XYf2EOUfrCICMGUkJ5Oh/O0u37p90WmNCHnRkpERPpuBKnVH9Vv6
FQLIxZ1IvtKdzInfg9Pt1OkvmwIcTCfp9wLlRlJjKSG1iab14dNxIgCbiVCipOxaww+3DJJiEJQi
UmaLYj01GGF9/gLcSG5eyIQx3DeDteqDwE+D1ezhx0PcYCDRq49w0Gef6kFF0pIcyNOG8kSI/5ma
Bvz+v5cV1qLlPl+kdwFBcGjkOPmUheez1WTD0e8qC/Rbyx9eB5i6DbUPX1/6XI/tRZLNzaSLlJMv
Mpa2F4VrkdWxM/SCTDH6GQgetOuv8G6YCU9dhr9P3w70JDGoWX3qlJ4rRDE/Fr1DBD031KXceJZp
47QyhmEShCgs3dr1gPoJeECsQGfOCxrfDXTUmXL2EbCxk59BwOc7izAm7YnQmo+nWlfC2FGfhraK
wz1+h0wYW3kwiLyKB8mUdvclq10bSA2hlHB1+hhEoXyJLADpSGaKGuKp+AnUSAZQYtAXJAdyPrqu
vHjjr/YCE6cLy8lBJcoHgf7byF1Mz10anuDlfRCgRuKzIxCOaaLZlvappxwPBUBHlbaPoGmJPStk
nOOI9h4u+9R7wCaBN/MDvm7YZ4svqTLsfpeLcjhBHi6STD3p6K0S3u2CijUD1pIM/LRaxOeJsi1y
kLqKM260RZRLEZ8nrqcF707bYdhNj3yvDS6FI/BvdZNTU//vDpzZHUDFw05u65zN2y1mJCklQEn6
7Ga8cncy0BUaZ68ACJnJCBUjr4DClRNqdIb/YInQCc5/WWcliFBi3cCAy2RyYHVKagJB8lNBmwm3
v3GfVnTRgOiWisJwrohLRDKu1bT2hPRfJ8jRskdvePTTD5+iQYH4moLbng5jPo3VGcTWeD7UGxWs
I663VfO8eIU8PGXzaPcrDdmM0rrQ076znaBEYZn00WsxLqSUhhoXh903R8Y8GZ2lmzzkmQixJDPQ
91jKWO0uxTvXdnEqVX/dmjqhu0LGh3xRKkarx+hZVFVDSa4BEWBBNVEZOBCWJYPPGqGhk1cV+Ctw
u1LhbPUsobQvbEBNaca71LTn+PlIYRMMXtcQrw94x0/Ju/9qfcDHCEwr3Fgm1yj8/X82gkkFPdbK
hCMdLbl5l7Y3nLRdqqeYDis2TpB3Iip6U3txI0m/2w9qSatjexBPUopl9NVFFiXcxJkkZztBNfxq
AGVvzWzzOUA213alw60zufRPJ0PUclkWt9KKD98oIikYdWk/ZCNBg4tTfU0aM551PlekSpNd/91s
dcgMcEfbovlLTeMspJg0ZBgyqko0of9Mb2uf7PuUnoaLDvILD7MRc8OM4wOP9rR/wELgxln6n1db
KdU0L+wARVPqIgLPZKGA8zNU0bF6TGrErltYKQOPOhwd4F/dy81W0hAQtL30UG3Qx6qH5Ya2cqwa
QZEFEQlee0W2n3JVlXAdr15K24RD3tENv0AVxMYU9QsQDrNxx6FMzZ9wFCERqdr313NXbtYmwIGv
xocuU7kxEuSicgUxCz4WG7Y6ZwNnaXY8cWsv9lSP5dYvJbRPBkwjMTebnKkziyEIcObQhjw1aovv
qOrQtKW5+1jd7xcBOr0e1wfmzzDYWYzNNA5LH8wPpe5MzKtPGLn3jhiRJuu4kKzbwfH+GU28k5nT
Oo1Md+3+UFvlCsjgaGUJRTEjghQndKzV8eJ/6NlR8RmVAy/bAsjoSx1oL9ZErjCnT48XwcmO6gfa
PCl35bhXmaET/JPUM+rd0UrHbjwFG5HjjCnmXkBG5Kr3e6iD73xSl535K8360NJp9GrVjytRXBFq
o0yskqIWoUP18cqL0j6KuK3AVPxPOSLUrdYUVcITw1QKM9wETaeqPiLGevLGIumftyQuUUWeZYA0
RWyuAodtM7m16T32kIZEnjYUV9n2CvMAm1LFvzBIY9yONoydHWPsU5uUUTYKa5mJx8EyNaSlv6/j
wcBexniD2JZVtazAjDVR9X37sZQ+MCYCjydIQpy8OT+KMhblbc+8cQMjVWK9xB98s1ErHu38cugp
YpFa8+cclO0BJ+OgTvvB/v876Hmzmd4oqgz3Bt42yvqe9+Jjb0WSZ1kh9VzSNd1D4sgPsDHB8Ufk
aPjRyeYl/+6uOQXO3sXn6qXo5ZAutNvoLRdX2NZ5CyjYHCgPj22KqcnKyBb8TNUsPaUruKHozbZm
YJMaxEn3vDhjkuvoDpUmMZNNdV3he/paj3MTZqHbSGgesE2mLPx4CTryKBKZg0N4SVMsgKE3r9ZC
uR4Rnb7SRGmhT9pJMCXIH7PsN4gk+xC8C72MiNvDwSRTIK5ICwznC5qDPFv8KiXxt4xjPLCgEBiG
IPbGXO1hieToPX1jjyrgEiC6eeoPZhsrNUjBeOXM7ERIorsq8PKBo4Cikq1689KTcQWCTydClsbl
Ud37xOL2v4pXCSYeXpZoqGGYH1VEw+lyE9SYtckgqE6V2ypBEkc7EomoOfw85ysHL+840T42CJ+8
l0Ec2npAfiyBlfhhhekX0rSfY+Jo7xbjybfXvV0jA0V2Z9BB5VtD7c2OQ60KNUjO2qle65Yxlp2j
YfacK3kVb72mnQbYlehz/iUlBQC6dtnDcrR5mhmofqz/H/zPQlMpYcAwDyST3yMkAQe/P0YkT39a
WQraooWExXTpRyO2EanD6bM2GRiDAe1pbacO8wrfxQGsUvmantz803fQrKH6cSeqp5RZ2X2sZwzv
BqB6HSoJ7WYMiKVXCuhWW6ztaOCgfLLmm+A1VNsI7xD6/ZM8MCcI1qrTMUHtc9Ed+hOVpEmtgnQR
vFJpo13lW5e0/n6fzmDs9RvPBFvzQ8qJvYHOtK3Cmdfwiwjn1qS7B7GR//Kj45lzjQuKTKmNAFQN
zbxmlimsOeLW3PQHBc4gzj7meIYSJcnj0Ivq1ehprm9hykp7vnUE5mcNnMJ+3vZptU0E2IE1xyoS
W7YW8lFm0E9xRlEXHcw4NUY3Yox3twSjJm/fGi7sUWCnJA/SbBWT361riPe4uTWZkfRw/539nU2c
fYSkyp45lT0eM3Xum0T1z8uCFOO2ZP4dPmfPkHfDXvOLjhCMk9U6mI+zRI9V8buVedTR7gNqUudn
3Mcvf0C/ShH7wi60i/IB63p0CaNc+pllLDNcNE+5IlFdsfaOFMTonZqLUypLcrFhHqY47yV5BWOh
uhQczeaHfTjRxDy80EP+m9SD8cogIWp9zTK4P0etyqjT2hAYVEzO929azgXTuT+DFIkn0BExSkIC
WyUy1vL3ab8JpTSihVhZgw5J5ikyjnX8u40TavayP2KQwKlSbd8lc+ggyU62yVVDggd47ntiFQ8X
YQyG1Rw69/UEcNUJtri5sRthj1OqtDCCRlP/pCRxn5HEdiXPJfvT8Uo3fkHWLDKJ2jidN323vU/z
Gzq3J/k+NPbfkamveoOyQCMZe9FUiJadmuBPMt6tYgrr1a+/CjV6LJdg9xj6mN2s7EnbtaLxfAQP
4anfRpwxzjfIVXcH8yW9ISGw2W0snNTx6YU52rHS3R5wEDkTNJq2c1hyegDgenR+VAuLbeL6CMgG
U4KCvWU9ULJbGdgEVXuB1laUAOU3Qnr73vqWmVnvfBUBydrQU6WVz02Xhso8M1MfkRTK26R4g37Q
CM7ldcwBYBSC4pTAzx6IzuY4Dm2f0Pf4n/eQXnJrFtdulxLh/m+n8vP80s31JD0LEb3j5AZ/H56A
V7Yi1HxnkdlRiBgOqq6FbcjAprSeB5fDx4arPnkra6BvXkdBV+Dv9IsIwQrMfp1KEMpGs2GsnYDY
O9gzwpnA1XEa3l8kQcaWVv26OhKxg4/KyVVLRt0m30ZwCRkIZvMV2dpTm+2c6kWR6vm4ep5LdGGX
W4DJv/fcWaXhlACTC3yZd3GpFGyHUUQXNkTxDNQukibNLtdmBDv48bVwdVjSpVSrq/Zmi5zY7L30
O4WEne1Uvtx2+zj/hDOj8EzSaTiJjPp7f5ISMaurFxi4jpmffmPGBnsqLGUUpXipVfT3F1gbiErf
0Aj1x1nCPVngJ3U+Dyj5HfvcOD1svKHQIHpWXMy8jPKz8f4ZFrvaEjFHqwQHtouDjA8TvIlwDAqp
DWNfn/7enLvFQxhAQAYE97Kojwks9sJrljaiS97wv87DPkHh93ov8ZV8O8cp3TuZ4xck0HSe40ma
IJvbbowMd9covYtU/3G9/EU1UMV07XrJG3bTorNZcYuYEkpKZ3FQokvMT2M2i5yl13jDRem4M9EX
iVfn7aaWjjpOd3z3JFiBgrKVTFLvFXH7P73/ZFFuGFaskmHZUsi6ophVkPZj4dFWwThVCtqO8RoD
dRma1xsNVhBlzWdXq0JEstEkK+QLovlN4mhdQZ8yDX+2ghOZIZFztVv/NcV7q/fH6j4H2nKK+wgh
apokhngUCm6KJcYiXfQxUnOiQPQwhzHRl8UpNSJ3oEo/ZFLxxjZJ6LZBnELGHrtY7nua70rgWhKE
zH08uRHF5i3wsUB20klINChHKi5c1eHUDKW5Nxwv/VlCXeAhgL3jZ+Vf3GxKZOY8ogvIjcX4pU5q
+wjjnuriYSlz5D6Xb+s1i+EdbtnVYriVp4aDkQar61Xk89sUlYOSMB6+5uewO4DzPgKP/YZWfXyM
1JL+UMsTtUyIcsx3AIYa5uZSpWZxzLBAF9NSeb7k6LpKU5VYuVyqUjwDEJkcNW/FSzQyRRNqkRgQ
U5Ht5pHNBDviv1WWT5gkthqBydRYNS0PMPyZWwlMYiS9vxbhxp/Wfph5z9M05Y0ZPqbmHpmBqi6J
nH64dVpxKFXu+GnHg/MbmFpQPhkZFR/zc2TJBNkwHZY176a+NDK1PgjqJbFy0IvOZEeArDlRb7b7
MOlfrjNd6jBXUXCjZ1B21R+cOa0+BkHYi2odfw6NEeYSmYwDCCOqD+AzQ+cwytO9MEQnZ8YwwGwy
4reHd2PULIyKT6/l/uSEa2/CYKjVgEg871t/8CIqTE7PWDPG3S/Afio4GHNGdX0u/IipJU7no+EU
Dr+PYiXd+1/2Kuo7c7U59fCxAw8hKnMOZWP62ejbt/tG2v3TuEJ6YQTwW7G5+2OeEA3oFTkTE9/m
oYW6w/3urz1CcL2Xuk9cXkNKbZsKuS/ou4OjDF7/gh8+was56tVQirHd9Od3/GRdsOf5+2doWScg
Rsoy4VjpnaS7RLP3xSAHGw28tiK9qykYoM86068pqxCSINA2ORhSz43HgTUhVToCxmPYtmT40faD
KlnNKDcNwBSXgYpsdOp3DV+IZrmKV7d7dDaHSAUhTrMoxAOnPKz+dKJzoaw+9zF0/7y2E/XHPU/C
f+vrj6dPweP2pialmFCVgNcF7pUJlgesgatrIV247anKe1U+yN68oMUzReEpKk4MsVM98vfbZT7q
P+EfNndH/fd8vDVcE4VA7Pzf+gxNKimgojfzemg8PXXl3ZnExMPj/s2ypzKAf/b1Fx8+wfDHyFgR
xWMlRcVFuMScrpql6+17t2X1RLPW0yLeWAJMWsW6AqfcAj7SFbaf/56JyQYofKmFlGjOK778wm24
UWq030GrlW8/C6tlE7KTMbIz0Jho0eYjxZ0uYT1GyeuoVPeevoeWps2n2y/0Jqk6t2eTQleFPnRV
jCgk/unhXDKilWftuq7UI3wbmF2Aq4qsPjVe4F6faE3ZRucI3MLWPXceL3sjd0rUzZxSY/yV60eD
d99ZdJfhXunHu6CYCneCPLmsPaM82MwgjFxzR2ZAEjIh46YdfqcVb2VXDvlJJkwfV/lH0LxRJ48A
GJW/go+oeKVgSyEF7ZSFu1UvgNl0ObCQcrIKLIGX+ZeCh/fBipOZr+Rc4UnZdUwD8lhVnOtk1ivJ
hD1C1kXyi0F/JbMo6XqlLU5Pvc9pATcn/QhRP9F68XbTuTkK9mfNb5hvJ4/zelypqAxRokhldRAo
129mz8W3HiQyT/y9acfCmoJJGS7Bx6XjPqWzBwyYmdDqi8oHpfuX1pRs1NcVXp2KgQ6pkU0W0KZp
iUF/kySVGaXlP76pMxk+bBYktdlOLRB85uNDYsQIIBbfu/PSNKuE8nFvPYmPAqSrq+2vjRQVe9em
OotAn/ukiyTKNwvs69lyhfZHJb0IIRM3f6NoZk+BAkpZPNVa05yr03FQUI4e1BbhAPyB46PcOMYA
5rK/oCnqqS1SzdMLNZncDXk8fI1fBd1M4zALaocuh4fZFrhk/rWdPPv2pyyHciHP8JiYwguuqSaX
+QlDsK5GtAdl+Yt9LPg40Nv1syQkEnJTnFOdaoJ79TEKNrbKTSuhTG8ZZSHukGOrb9CteDkuA3Kn
r1Be6OVqTODinYfYTuvj6VmoveDh2J6XyXERm+FgsxP0zyPEiTV/qLFqotO92C94qJ3/9v1qp6hq
3PkK6FVTdOnftxDWp5g9kyrt9CT0+ozLgk9YncFXx5o0RF9Rx3598QsW3ks7MhjJiTnhofERh86k
OrcT/hxp+qfRl3CD5tF+TqGRlenVeojHZ9gDUZFcL4lWBhf24YEaEHWSvqBX4bDgK5qhz57x+5qK
LBN9thXhp7Krk2oGU1K5AhnA6U05oUJmOMtiGuGHpQ2e+WofFJKAhJ/qNPGLLiGYSWNXE9fG41bj
Iv0rEbA7odPbPMK+Bqd8OkDqTd4JmhxmxB1aIUobD3dMTAKVeHzo/x5AplEx/dz7vQZZoBXxPlSE
Rf5AKV0DZq4UUMJDk9Ya5+WQgmrcP9eO8jj7kqklOLp40J5nE4mA/JEnwvnOnyLf+DcXFaqqexOD
O8SOiIBkOgErvF5BfiSydiIy6lg/WmJsHGwYdmHD1RQB/ALdH6sIDYD91+mTETDYQD9eTl0EKwyL
Ik7yZWRboRnkGK0P0bKOANi9+ey9mF8qXG090Kk8cfLkdV6ej2A5c56qwSFuGEqo8eQKIv0W2/eW
V3sN92/pjRMcQ14YOptNEoV5og0T5Ktxw98g5NhMPR2SGTOdNpZO37Qkx3L6708YTngAU6yjwNxn
K/nwCPmFD8rz+ZCftkBiEk/Y3RPtKa9gCGc6jwCLWSr0y5ZuW4CmOmR+MBEdrfo57+xsOCnNyjcf
/kqg9Mb5rL4yGdJdD2wIO72ImgJhWCb9PlMRNPKpVB/cAkFkZiTA95MPWr4n5bnx75eQo4ugHkPR
8idNnHPay0caGErhQAFS8cBOBcRnz1GN7ytZv7fLwpSaZb1VnkT1usrYm1wPxT4es4YUpOsBmPPO
AXBKd4w1PCZS+ZUE9OHtq0h+lmBTIntIZFVwYv9kMbmiTL7doL6NAp73sjaa70BgkyGCv0KOGQcs
9GvHZgqIf1ZAmduIego6Mm4DBvWTAENtcgkJgnaBqcL9QsUi9gHlgDOthSc1P4FT9EE0r6E2roC2
yoVz3lg6hC65rAIqOf0V+D2x53pIze5ea+sTchQb+lomaafz5Ag0wknt73+lesAB3A4UHZ+G0Q7q
f9VePFBIO/2aFScgixKLzeCMNuJRHgoGJVXAPm3BLNSah+N3unZ/ns/CbY0D4jPQj5lcBAETVddo
Ajzh6pqkm4tx4KskpTMrQyxGrkVXZvKo4hMGASneeDGWmLUvXVBBAb/mgBx7q8dosF4Q1nlVcLgH
x7PeflcIJ+RWoXhcggeXkEb00d8KHRszNLcR1hpCMKHCpS8Pa7lbuijvy79V8Pe9mTGfCn4YIphC
AxH+Vd8SF2zdX4EYrCHtuaVe0yiTKl0LYZX2LByVFoYdwUvcs9qWsEmjiGXZejtzrRzXXiS+/Lcz
2iwAEOVAqLicfyaVpxaLC6t5zRVF7v4ml3AYgX+oivcWikaXa2X9iYGL3gNfvD8sTBFDHywMtBEu
WilUdF7YmfGSe71aJifxklwufeaoMs3qscn9kfKf/rGtfpL7cj5TYQdR9uL/JkErpxJh7ca0EGGc
NkLB+x5oHFp9fRER/k0gnyQuDdTukA4jVnzJ8r8xyjAjkXpQ9Bkv85aY8ZTwIYejxEzhflBoWC+s
LyqIKevGcaW4t+kY/dP14keVB8pyT5AsEamGGT4x+6ZSosHsejvD4mdY5nyJSWR3oDfYC8RYAUU6
V7Zq4J36Eq4Pw+AkZu19T0fMuuoY4+Qp0EztKC4FS/VIEI9FyPnt4nncs/6DhC/MPqOVMEGCARNW
PUeeqsV4Wh6k2f7OEGfYR/CiPG7r4LLGeeZlFBCFvA+fA+PqwEXaGMVuW2mjSfJ2NogeUlzmC2lx
X7bempAVS/cLoPkmACCJbvWbEvb5WenqvOxTpgXdXJuvzmV+wFDs59QHXzRmZMJcqoKgzL0ozbr2
ddQT0F1zgCTiwRD8qaEuCYzSAJbi7xQcUXFVFpE0DWza6aI1EvTfW5eLjUJXsTKAw26QqxlhKBJ9
zc7Z/ySYxvWVAtQ0W6saz5Fg+QLxHB28f0a1XPpWhwkUikfFmPn0Gc2ap8+LDsziNZJCAMQMx4eK
tKeFIGAupNnen9I6co5/WaQV65FfAsWBF5yE1QNxoc6B2iGwYmQAE9qVqpnCbp2cFGJk5bs9cCtz
QYkbQSQ5qCTEWPQFU9/vqAfEKCRRQ+qR/7UFHkh2Z4DOp8oFP41X8/T4wrK+feAf1ABjuEosqVr0
o3W8c5dSluA1U2W6mm6lCEIQ5RwyLNWl5Trx0dpOfP/ZGDxlIBk+8jVpKI493GZpFDr8Nb1honN6
XOOkUttzcwOgYf/qbmOugQV5Q7+R2JvwuI1sMfG1FCQdkEX+zXmq4QdpPU/dMuGyUxU2ve9NDz0g
ItQH6Vs8x7Qkt06/c5ShJlYq1uePyhaN3sq5jaib3EquDbR2T86y1brtZcWyMLXCkhnwxAjoPaKy
CSiMNzHgyxn6NyOg2Yq+K4ezJ3CuXln6oYX6h0rn1OQ8qtQify3NGUZa4mATHfW+mfsVrBcDx9Yy
eKpYbVVG0QllrCJB9i9UgEE1VNGfU1ajdYKFjokwVMPFbOoz41lOjOqUFUeY49JDmuCl+IG73aRy
d0fM5ZKH15Iryx1VHtyAH3jUQulmAkDNAdAVYdJMjuUoi6eUTUFnVWADVDokuq+S9IfCV2bVCNxQ
8ig1OMgAxGbRO9pjdPlkQlTjtpfF+WtfRrF3uf0W1/iLMizSYEeodLv5SizEa8OlFuPseV4qOWqG
Yq/lj1Ll75rwVnQ4mepvvHMr96YNLN11lV9m2EZ6CtzlRovSnXQ7lj/BgeXRKbzimsxE7jqgSsZr
IEWEzZDV7+PVzZAr+jv0oBXmRROLWNJyz5iU3vpcxPBiUro/b13JKql2somGBC2yBy+SNSNeejJr
poOL9Fyw7PTS3wbabBzz6yhB+v9Y3iPrXI4RwGs74OLhzbxX5NIovp/e8MfOqoXGjRswNNhDo0AE
4w8CwrQE8yNGaXjy8pD5vyKBDnfAcCIqpLFXy0OB4UMrJgqg7wrjGZlPaxbRI6fLnJZlhUuCuPPa
QjjZmlhn59u48lRZ3m4YzRUvv3t5OBg8/0j6bHSbt96f8IyFlh3McnS+Cjjm3jymlRm3bsIUGAEZ
fsAcQCYmVc95n671lzGIeisxvWv/HfbsL1Pow4o7YtmbJD/bvl+8/MFkLLw9trgFNhEJeTTGC7RW
fMQ1QWJm/3eJIbj6QFnIlX1t8FxYmYLKh9Paui6/Q7xT0fHMssaT8Pn97z0o9yZ2X4JbgzxX5Y+f
RmM1MZpZAUQ5xhrdhSWbG8MdPVr0vJTQChB5gEXMuiCivsmbRFphbZ5L6EQd6V/p5Pc3V0FIYjGV
KXcCrFKGzkxsIAfRS4seJPBZ6u3lcBwWq35gnXeZ3+5DmbjtUmQilkDhoD68QcdJCQWFdraYKLwW
6QsblK+9TlwQmEDJfg9UAss+Z/70ewpSqRtTYGA8E5Ef7nHRksh3DBpaog1kQ4OXciMc3e+lGSAL
o7hU7yCtWKAIU4Hj7Mz5nt5LlTVkUDuwC0QmJRnfKlHq9wBlYyCNlfazhd17g6754GtaBN9BZUaA
TOzf4F4or2Mmon2H7cVCSx8fMd3xMTRkwlNJuVOBSjqOjJFd/KPADEPzBXrAUcTAw7MPrPGx9uTJ
/3I7Mgzetj5IF6ZyOoILLckxUr/A58LuqN+0t6xmeFKSfr6uqs1bPBc6kCD9wEaND8kWjKn+6qr2
aYwMc/vtn/z7+V3GVcErdcvtzQgSL7Dm5azo4gPtmHOMj172xdb42ivTHnq4SbY6q5nhNzIr3VhC
mQJUPe+UZKvjYxx71CJu9XIWN+5Rkn4oH/vGLD08rqmJHgxjpN4m22j3V9BxIVZU99laYS37AP8u
rGoIOxWiGkyrbVUR0jmQpVm5M8DMbE9Z3hqqajfXyEFMiQN+JWRCXRchSwACOxPQupvx4SiQyh5p
wnQszmnHhjgURf4Drxc7eWbv6b0WUDKZHwLfg91TnYtw87AsZgpmpL0ME3Q0txU4YFNw49cHUNi1
TVQDv54Mw8G32M5LS0Z5aKGGBG+0FN7+kDyP61Su1v4PDZ8U5mCgK6Z7jg8fVrJ9CvZA/YwPxn4y
HqvM+Bb71e+cCU75ld12n913icUMwnaKsfZKbCHWYqnc1Ja8WK2tWQTmT1xrBr6eCuzk9qk6iI+z
nhqhQJizwdhPKVxgs37tL1PLLCio3OnpMljWe+XqtgfAc7GBxoSntYHPEG0zAjFFUlARqRU39Y5a
urhC/scHFBR2dvjsQJUNmDsEWj55lgydhDrMpD4xEUK9mZHRLgxj/Tk8TUar/xuPbbeHhNQ+gmBb
BRnVOpud3tZ2G04ioefGNuxJT8dh/r+UhFQIaelGD+imKrqV44FT8f8cXQVhic6FrFDkKwvTHCXw
YirQ63bDQveNhCiOIpSwecbUotulPZWBE1TdriHdQnoEshcKfBxo3FCEt/jPr5YHNcMMPu0dDcp1
I0eJtY455Fi1nTm6L1vtPlplrUOGRn8fi+mVjh8Phc64w9OCJEDpgPkQQ275x1ktvlY34usw/6/r
O4+iDCRLHYNNwRs8Hrujx2EXWf7d0VEiy48FsDIAa0UOn+PBxSdGKQi5lEKVqwSEp1D/16Fk2tps
ksSHB/Wtn9cljANRHdzMToMsqsuUhmfEov+1YCMPHphR7e9CGqteLLhEAWz3HNN4y7+RYWNplPt5
SAYz8zcQrzmFek/IQp5z02Ljli45ES30QPggt92Th6smjmUBPH6MBJvA6SmyO7j31WofWANZr9TJ
7Kpxdb4l3E0BlQYC5slcFOLwUYtlwLNQpYUUc4jMr+LR0cnh8GY03SyKUSRqsGo8OBudGuqM2/Yr
mmJi30+HWNk6QlnkQJeKtOXbCZ4yUHvumbh9YhVHJnm8k9deY30U7TI+V54zWte1CI1BfGza2YuH
1CJshVwQQnoY4Nj42YuQiJFoxIcLyM/YauEbLsrIpqp/nDXna/v0HgMt5yG2XFnPurYwHqhqBHza
dyQnCBEd65QrxD6E4OJLM5O3A/YMdHNMWZbMlH/7y04ezknUBFC4dakhB4Mpx3KVMX6gmAIZnui5
hW0ADElhdxtMjNniQ87DiIxCG70diMhXeNQYVhb4EA0WpermKCG1GJ3FuN6vTrVYE550AhT/cHs6
8WmUxbZHdZoJfkwihcImQ3Q6LIiYu9Qcf/DTwh3bzmyhlwshO1Ew9zCVMgRycLpnoz+7AwqfQywj
VYs8GfagsWPOgJWihCYVMJMzVDCaohImQtKTJxo4iYp5jMnV4vkEa0ZiDe/jCnJxaXF5l5cjog/6
OTCGXNN4s4KChOqb3DUCaSGt0UYrssLfuZn8gqCFTbAqIUKhscO/XvCO/69IbJJ/3kWXUQgv0CD6
q4w+Mh+s7vvj84U+Rck15upfYyi1YxgBgNSFHjJSiIZuVpPv3qj9gUHLThAQ7wy790+99OTqX/RB
nyDMLmSLgufWpbDCkxO6mgcZPWNBwqwwup7MoaCctSF9rRQFRPIdloJ9m46dgryakGd0AYVv1OCM
+Lol7y+Lxb3yhRXYv6LexQukU8PYYkIgNPR8X4SMm7Ujm9lFYHYi62nSyu9vsZ+yvakg6uaRMdUl
oJugxGR+KOP7Z/y45Lcui5MdKV0L2S/+zaMD8jJ0tvDF4jRiQTLJsvqBebSotVTuTIOKKeFBPBZ+
3d5IHE1oNin3aROoVgDBopWAgyJaFEJrh/6EA/YfKuY59NfoZJ9lq2V0Bzr7rkXzSJdef+Sx1VGx
SRP9NZ3OaJ+RrUc0WHn2FelRS2WPWYim7/Y/zK+PLGd1bkqfvAOrcuek6Ux17CytSI260ze6XUUD
7yVGHrN15cnCZTwUZuj7OoC4bYw9YpI4XdBRH1ObIxiCS9qHgWn2vHU4CN4IR317YXLK2HJqAfs/
FVfYvjFIxQ6xhUGFXjkHJwNWKzQ0wY9dwseyj6QuTFsMCO9cMq9pW/Ubg4PCIenG/F4GnW0mdNVa
nuX+GSrcLF5jMKBXoYPRWAlK6j+cX2jMe+byInDafftoUixZPqrxz5gnkDoM6KOHL14Z9HbILQe2
Q3IeOpQ5lHF6fn7s/nMbOo+S4KTLjJn3ZA1ydh75/SeilyQ+YTXq1CVxHWONjHFcfNrAEVGxPX8d
9F5y1qCPQoSOm989H1k8m7wmxW3hpMbIEyvFSsV6WE4aT5JUcBf17fYOekwCY7FLDMOeQOCqKHCq
c1tz9Sdi1oT7LDVgUAnlwf12Ekh2rm/Bjmb9lZBa/kwDenrKGLpoj+dvGnfRzqt3TtPqNKEnp47O
cvZt5f993tI7WgsRXrBMAIqLQltvFtkjALbeJVeEzMrguw5Ts/pjaUFl+hhbDDU4uKeZRoKxzyfa
SUnydL0+QCQU+WrAwAI/QDNu3ItQYd1qhf/A2FiQ7AL1lQ1K5mlUaT5rSeZPizvGtexX65ONTM0C
Y6m5G4XBlm/52DcL6VMJJkF8UUOvZs8mlDui12vLhgbNSM1JK+OsO+0TGaHWXMXziqRNIkn4thlq
SsnH6YexiXYLRLfXylaHfrknTDjcGgJp1LZ+CoJiy8EVEW9UGfyGD6T9l0zaN5EL/kD3VFyF6GKs
1EnloBHvJxAz4lKb/wxwd5S847CQc5VKn8j85pEmKvwv8c1lCuMkg29jQ1BazFXDvj+OtmDcVwYZ
e3/aMfw7uvROg5WbAdksEsQNycvsJnlTWDWMSRHLkSO4UoUGGLtjJE2VVGh2yJay3xvUrw0wRCLc
zlxWQMWTEytzk7IXPzlIuuA3yo/vACHWw9r94s74ECzCvD3M8LPPS8ge2KbSvuBlpDAwZEqeCXW+
yM+a1nLS3yTMpFgvolUuNEHyussMGdH+wfBxqHB07aPyr7gzKEVtdZcjqS0Y9Qbt9oyImo0Oc80J
XeQIL75wPm15JcyHvUbPxi7URQzBR3m6nEur1SVPGOUeqgfYV0ORq6fT2/Q6GcL+Oi04xcM4ll5m
47han/lAhBYW+ma3WzPBVY7b3Y67LlE7lkNVnTr0yw2y4Yq5cp91fomywYGWfkZUE43XLfMANd64
iFow/5v4JDLwEQg7Q4E5KyK3gN0uQY1M3BZAKW/Fc+5JAPxUmmqoZmY8jZwDdF8uZza64in4Qj1+
9T+3Opl2QAO4Qrx+wJD8Dx+EfVUW1h1uz+gRLp7+iV9Y3XTrRdVG3gbodKL/r8siJz0+zV4BXkiK
HA1/xfglqhXQ6UvP1BX8kk5SE/rh6tm3FmO6Up93KW5752tKayx7gi+SMHxL7AGZFt4Ok3AH4z7b
4a+62frB9oz7Gg03xbwhiJqv1VAq6w+SE3KEl9oiGm+uLV9muFspqbnUbEcw5Rv5sd1coyfvUTR9
0lEC2daWUESgJzVMEYMse/6y/svzM60ZbTKNPIvKHtdsEP6h1fIfnoo6r4b1E1okYOVCVt0Ixucs
/kD+XHWYGTCvAsvi8+6SW11ODiyMF9c2/Xbk/6VnH0tSnK2FjaR//yItn5F/hey6WbyS/q2VmbPe
sXvbk1ndsE1J/qSSnoTFgybdK/1QBDCr2wmd/IarYJ9ZDyuZbPfMNU9ye7SBjshJ9oi5UaDeLL6r
yfeX1zEFphSEknIodiqJH1wDQ5B37tRy7ikeSsTu1Cjn2iGGKbFteIZD8Mp+vXW9mbWSZx2hbuoh
RbTu/AR8Psk4SyXtFl7RE9WCnay5xTTW6VYvnS7EMda7g07n3UQ1BJ23ogHzDG1mbF0z5Ffs70MB
hdfG3xEv6Wq4uH7KOHW6TZ+F4kfsBlsuHEN7yNxGTnKnKGM/APj3NQT3QpiKZau5IO3wtT1KN0wN
iZofelvIhhrMS5lK+YITu7Q52SYuNt/c+1RfrSrqXuvlEAJVgt9OCLVDPQF4dHJ6c9R6cbWvmBkB
+a7dfpHfVamJ/u1SYYYASd627jHZXhvntW07HzjF37QDlC2QrYeD+YirR5l2jfdmKv4h3HlZCTMZ
xq6zhHGxF5S55roT5aHVJbwk87MfP6KqLPsaU+/OTLDosIDizjyTGADoULH0rPXrIYjXvgtof8qc
qzMjpDc+YKIlhGYGMKwD6H8QzlBbhygwdxTYtJrKLpOz4t2RIu+orFzrQ3it/q7SUpMOV79tiTIO
/pM3gxpvD9mY1GVHdl7/Y4V7KW2h1pCBT3FlAbA6SM5/eScXd3oSbKDfBEbpw/DKQaFrQn+I2bbv
1BgYbqZwRLKLsWXf7FOQmcARHWGTz8M9q+vgcb+JkAKEKZ8iVu1cjPEJC3mOX5AukhDlS/TRMhOk
bHa6LptJBsIADFmzC+FMTiHCWVn76QLLwJWGg7gjLlo8zO0EvqDxd5++S1VnP5KEqrkKlogYMgCd
tDbu26hlPaTWRCc4sTMjoF0ztleEvjqaM2vFHlOALLCONeCE/ZID777oG2KXHlB9LIFhgYzYjLp8
+qSUXBK4pW1+ropUGUe2i3JWjFIU9LaEAFMOaP/qBFbvzP5gDNmOTVL1oZlBi3EqSyXYoXhwWuUM
lUZAFUg4aJKweEhilKxj7Bd8mOpgUbN7w1TjAOhVZ9vVFsrq+GOJrcY2cxzvV/rVpGPL4ZTayhQ6
mI4IfdA//i0K6Uz9kEneI8zY9RAIKTvvrbJzM9FxCe2cihzvWkriVYLDsPUA/7Hh8P0WQJNPcMB0
kBBuiyWqo9d9KXkiL05pqzZRCXr4r14IUTojtn4XD3mKD2Zd2P/vZ3eCDk98um6G9Ps7L2zY/6Kl
MGSYqUgkhF/UipVBnchN9DROuzfZk1Ihg+3W85kTNuyGG6NDubzBQZKuUsDUhxcI/de+2Kbxj/Lj
anU8k452ySx4y4Ahl5PYlThC2RYhx0sCjaND9dY0/pD1Gf8p97aYfPHdqeI1rTFdmC/LKUDMO/du
gKYd63Wv8yQH5mOn9ZA6zgC8uklmJjhQMi55QBz+JATg9Fn1auKvvKdodxry0SfRKoInKxPcQs+9
UV0QlQgVmzyTWPTOVMi3pznpo+bYm+QJb+IJToK4Gm6dVAzg91eGt5pWMC5p4F5B5lA61ooUW1Io
/ljS6xV5ugGB5RVmmJjiFfrVGPUYEJNBxGc1gzLQGSyNnAI57efoSh6cAQv3uApzNZBkJCwnAykZ
do4cinpmLfsFu9xiuB8o4uQE4PavqhqO9h1agQEUfebmY+v52IqqbWtzT2Us3ulbl8PqH4GX3LvY
eC8H2a6NkDSzRsgEuIvVGFQEKYa58yzvizUQBiwlGIQs9G/M5dYnNAhfGR2rMOuOrrT38Cvkf6vK
Q5mbp/GmoGkbMBYuxtRfaDXCrmkSavzCABE8HGrqS7iavYVxg/y8Zw6Dul0QEW84Dm5+GzVoW9Rc
AKYoavAz2CiMrmtvw4XFkosf1y0M+ePVQrJoc2IX3CoTxQGLdrxtPbxgc5j5XG6ITsvVkpNVvthH
TukfMaBYMDOGWwm+CRzyMyLJZKusHDiTcYfV8BVhyXHTNfl3lYPHRDLhzsQddXxpqgsZzNPZsi1v
xPmiPZJyMWDgS7rZy2eYJc95Mefgn+5UdBXqUUDUgTXfxZqftX/AmMei6WyNKtFDGhcNMNMgWJlc
prK02OJAhfsD1XYOXvvHFKk75bpVYpL6/B3SvXh6hYmpFiIUp47PemjsCCu1OAdVz+F/GKv5MqZh
WtMotyKHC2udLuRbVx3iT/B4YIdYO8GwHzyhYp9eovz9Dm19uYfPLBTxnxNtRrkMmrEraqL7tF/C
ROdUWkbafeVsHFub/DNT1R3jGd4sYOA2iPg9q7YqbGwk5v9k9FEiYyLo0JbhKHJqtT1nmxcK+Jh4
xcQ0PdPkjzbfEZWqkZGxta3v8uaCVUO297JGcWG4nRdfNucrGuyVjS9A/U3HbZC0ektB2zZhYfY2
Q8HUu/SYPs6rZzvPX2WDNvRHSiQ1uQ1St5xPjWZvMKmIqD6qGu0gH/40FSej8vpW+x210KTejp9R
GNZuo96tVzNr94P+T8OFWojnYZR9cC2vLOGeqdd+AWR72XrEMFu2pc8LqMpsfYJ7Zk8E7QrTRvuJ
uRRvxfHptVWFPHkxMGIfum/y4tgMSultk8TawtqrZr2UaqmJN1/DDVBBVcrvb0OMXQ07feIx2vJM
82fatg7KKHLHkzmwNKRaWmPt6vajZXaLWqm/c544upP7DPJNIiz7NAyOqsir6biQKr9+BGUC89Dv
b10OF2N68CU8xehM/PzfCX2CYLtFR6DmhoId4TdfrBWSMazV7duBYT+cXlHTuHPtaAUvcJLIUbSP
ToPva8guhF4zI25SzG5bO4Qjpm96y6/60kEJAC5ad9+SyJ0YDmP2ZXD7mI6DoRw4UBwECVKWwjss
A6osgM+gY07cAlX50AWIL9yBmTwFnG6iVqp7Dfa8dOh73EFZdgudZG38w2QH+0Oc1Laoz2vNzdd+
tYkFobK8aenNoOoRL9EgN1GECx4x/Zz8lmYvTBggcwA68afG/oPF/G4kqW3YtRlAtN0TrPXoEUIs
VgGGAsFLUzq5OHQqR+/IipsYcGSA6e0iQj9t+vfdWlV26IoyLeono7YjO6nUh4556Yrr0AE+I/yJ
gyYC+dsU2qEUVoNlks71T5NLQ2kQ1Cu5btFxJiUiceWqZJPJM+mEqdY9AeS1hHnuUwUX3/7hwy8x
fgQE0+ihdYupc9piJcBXoyDqeYQVC40aBCA4OaPTTsuvPNsRe0aJ+/joFjq96lQPYQm44vXqskTn
Yag2Br7qBCROdm3C+FT852U+r4qz03j24ual87WFQgRQwtcBMlvZkS8Jnbd+VDzdOc5UW0yULJ2M
64GVZDC6gOilsmaulhxmBpaLLyyP7sW6PGFYDZuD8JZmcRJlJUeG73AyQbf3XnXxFjeO9j6EpXJH
dXXb8VYOOmAj36cRWeg3ry8DQMWb5wK1gFxrPhcA1vvjtunJQQ6oC3Zm/HeK2666yvrQV2n1cxOE
+HEaLS/NdQs47Rr6jsnprhJWUFcLZB5/xrfrLZJfV7avkLk0NJ8NEDqOQHVaWYDPpR6FTt90YOJX
NkX/7YmmY0CtVXnCF+aeHLQl2cm3McV52i+nfi7zJ+ru5qHjBDdjbkUD9eKp20FCNvXNhO8W7QjZ
kLjhFrbWyYmi7eI0PzDWvvXY77VL+PgGtPZWf9hB2o7dMQRLsEfzE+qIkTDBk/1sSuVrI6uLwntV
CY3eF/QVUkzDHQSefFysUlg/pZzTtyKgpV/rgtGihl1DurBRAoQiB+K0wzoMtNU0R51d2fDZNNvo
ruP6CdS6bF3t7ynnYES7E21eV5h+1dGtzkkCcsuv7O8jB3sYVmEnluYw9I7KBHfycO+WaBRS1MIY
bpd7oBclWGfsa52bFQlWn2Ee14QZ7AGZyFL1B9rgifYD8xjzhjdM9sd/3gFKy/92fsdYmqxVeFId
x4L2/y/+RdYWbobiXKBVjCcgPf+qUZ/tynpbeBOC5T30UdtYAwdfgnSeXREIRVARmCVn7qgFbOJw
bMilUKEW7qMFOcBtnwgd7TSBzV59Crx0YTTZH1st21K7Aloj20lKN0yNreY0VvrYt2v/Lp9qXNcf
DfGsJ/C0e99LnjgyZoZNMLhxkvTABiV3IcQbFrAjQqNLepRw2WYGa22IR0XtnYWwobUlgjOFPD41
BoiKFtd0QZ/dB6SLBV13Cd9K79wA6hmY9MLBJowO3n7MzRFN9iVUI9eA6MQNsPrV42r2C9bwVJhL
PjV4GlrzaBkfmTcm6TzT9+rapIvrpzf7NiBwNqih57pVzJ/jhs2Y9ya8l16f0+dF/BC6xZ50RLiw
7YP+V3gIBhB9HABBb8ivi3u8WLiQXut+Y8GrmD7KnyFe3C6ZtHNBv/UFfFxZHxFla332nSIY2vyA
2OB7Iq0Sa05B3cH1OjatzSzMh0CjUuYi1nRXJpt1Pdjh6jOa7Hm7yghKcENOjrZ7MuLbZ5is/gNl
XleKtGrbYtIBC1hqrdjgFICL0D7ztwev6zHd9avO5kVtQuAbfpPywbbIX2BPdzGcdCEdyWtq/qQz
5RIUTmnWf70OzwO2q6gjQ+pvXaPF9doIuRZKB2RG3FU8H92vu999uXZbta9UfHJuCzizVR5tkcp6
qX+8yBTGCmIzAFnId8psHXaH25wm9ZOIHAFMvGzfkGgXbUH/F8W6kpbQfTihQLE0BFiz4tzUYQ1p
hdbsBfrLyvDoN4xRu0jdYIvo2aJB++QemKB0ezdJ3WSOwHKNJPEfn0q1MQo346vGKi/X8i5ar1Mx
Ng0DS8SvqCwC2OKWYs+yF2ahD27tLBEo3OKgiQV1vW+CsajyKgoRQh063L/4okvlh+VrBcBsXY2g
lEeeik9WRbhicpORPRFa/wrpDsAC3eSi++XZULbSmHswD9rC7rszYPKDIlABD0mWUon9FX0yX6ge
TkzJSyv64/9FWuV/3yIDa1AzQg3BHhzXmOAvQAtDRquyT3rQVuonIso0uPOW5mOR/E5OnQarI1Eh
EkS/PH5dYw852nf4rkEM0tTAvhuEqmmyOtAlNLIB9z7RAVFoxynQ/kruEFmcKU4ZqiQR06ZpXqq/
8m/5kC5MeZSGNVzTqU/u26O/bM/a2W8JCu/VFDyQARIQDmbH9iRf+DYPn9MRIsB07fQft6Db9xlN
X7YBs3zThTsfk+XKcCo1NqGW21Ud23SeLXwHFYoFUg2VPMYgWIw8I2+2fRoecj8Lt+eJBWeWRj+Q
IY+5Vm6BuvodxWx3P/JrODfoih2dXDfuRY5J6y9n3RhXCJvfdtEWgYAa4MK5L0cPbv5ewuEKwuDr
OeaJ2nAbVOY7/XjH2CxzKOKD1EtgpnMS29ihuEK/+wAdvKHvh8wnAPnj7p2XqReFBdGKWiY0cqw/
VkFiJhC/6MCr1VPTneRcIbGQBa1VkWBdhJwcHuu/lpef39qOW+shF84m1wQM2m9a86UEZb3KRVXV
yL8oipPwyF6Cw7hk+XNBClgmRdWBBdH0KpG+/Zrs5VATkVnW4sbfcOP7HNCSrqDNE1xJLkr/j4rU
1x1BnmGsgrKpmKgZF62zL5m6u3s3Qk1RVTxJQP6JcAS350gez0CiEjjjxYzxlQXuZbKP+lUpro7Z
oPZX52IHT3WZYwNGOwUtQdRRSDpPFw00B0DCR6X4isb6/FvY9lTej+Jmh8KhEfF4iDcN7xVOvbcM
WgElvvbZWV5exCq8dcmXb3ojEpPooLThUGMIf452qObpp2K8MQ/KHATxFh0kma2DE1zz4JwVPkRg
WSH2Ty2M5wZB25HsuLDAFBbH5462rQcuOBa0Bh6D/qrFr/mkh1MUvoSwzikA3rdzAF+xST5R73dq
O9GasofiaXQPHWsANUDLXAg31hP7lftvUmrMgmfWZ42teBOy4PGLN2osOTKO0F9nMU0SBHfESwz5
Gm3sugZnZJj6d3mRecT3oxqBY+gxJ8v0hKfymQvXrjJvz0+KZw1pml0M+/X4e2rbwZauvv1Vo3Ch
GYecMMr8nsOAWcdyVpVq254tYCMjJRwWL8+4ulbbg04szxHgdXYkebh0AbYtaGsBdiyb8azdAog2
BssMFfm/YKRRcGGfcwg7n9f17Y4tqv+/Ybm5yH2isEwPbc1/Xea5wutgQHcDB6y2/j5G/ymAsnyW
pjeFcwIzWbiiy3yrHwGD4yE4halx3u+uJV8+PD7liuJDxmfCKpHRWPI7jryfOTLGiKuT4ebXru7z
GkPagNXkvbzuNgH//adlX8FIRZXnFCQMuc5U+hsMkn8I7FuvcRiZH2jE7Z8O0PpUnCcS3ZIoKLwH
CBCouzkq8ObcFQ/b9yiTwWmU+GDMlSLTh1eNNPrMz44Ay6jpWYCYFdNY4XWZM+A4SnoidufJNGyl
7yKEbbp12nc8xG/kcBE+cAwVdxUYYfMVZR7llKzmjbGt55j5lIboNYij9cJ3OIO5gMWgW2gj2VdX
BrCyMwW9TZXyMcgHiEZRKV3O8co+pLXNjT7HYNPMq4Tu/CMQaVmAb/PoGyfiYagKVB0Wlw5UTJhB
d/1pwFEtUvtEuuNmZLnPDRlpstIXuEnVyjLP6bl8D2+ygKTMjPKSKDJ+eylnuI09VYSLaVPbp7UI
dUEiqZDOPYQV17aAatMF0aMEae3sUHVYjAtQY2C2iu95+dYQMe9BED/lYdsEQZ9jGVLx/RTlxriL
FCHRlrcPgNp0JM4u+gljPLA870QWr8uyOC/uX85qyMCdkxIlQ7Tz8wDTQUOv7MCSXryD/E02XUqD
O5JvFlJSFv9mdl04ysKXCgx7ZEOyJL0Ffa/DGUJb3i+WSILs1J1C+aC7TijAUB81wRVGLI6ESkn1
/L1uMjJzRQNAJE88Qpp2CpUBSkpAgccFf+TeOhI8Vnro4JTQWtgcZ2kHClN8QmdvQnBa9InEyBPz
FVdlrcfIVpp+HfTc5MfZA6j8W8Cd7xgl0UA749xzy8Woq6kGCvq6iJWlvzLeKDwnwcuzlSrxMQ0Y
ZDv3T0fBWiTAIlzKeGkTA4EZJ110cP2HWz50IVaswvYkvcIsyKD2bKP4zCb9GPEJTIP9vC/mV491
Is7YxeC3WHW8YytULridhvd8d8oLQ0wSX5+hmLi03gUFg+DDDT/IiKkwz/heWteR/xlXlGhZfgYq
LMm1mB7RZrKoLLSwa4BA3GbwaGCzuuSj1fB9f8GU2M+Vckqyvs3rx1/m7xXJr9A1acUWLSerw2s1
FOeZUm0KHp4WnJN6M5p5zZ/aQ8dTBXGsUkA672/g6KSc+zKpma1XfbCuJKIxvJkrOs0jgzc8cVED
eM0Ky74AKleKwai7gx7Q0k3NCFD1CB9zo/vSyuMJTrssBypABRIUb2LQ4PeoQ7gm0kKs1KzNcqom
cVkVatrOGV8Tx47ebIl0rivZDQiMAUjMdNFTTyY54WrMtqnTolWkbuzO7ECzx6JcuBt6SEwyHb8b
qdKaW/5nvl6rDz42WNiCgvoQjZdrG81bHWHzifKu8OIs0YyJBbeyK1iUQkCDkQEqyI6QmarQVOsP
AXFUfjowza4zv5gwuVLQO/2r0HoO0hJRFFTyYRZ7jf4TrjgJPuJPyshtQTpnQdCQQ8xk3EkcS9zC
OkIFwvg68RZ/ZzVN6ML5CaNAmD3sDJEXeCiFWqgQuxtH6UKoEb7lmeocsH7DHLm66dBDaA/Qdbdy
fP2idy2lK8RSAXo/IxVaHQY9Euq57GgQHHnVAsfI39PvDA1ZNI8Yem9OE/2MynTetoL+0+Wy7Hdv
kVxczez52O+slIHUoS4pDNHgy2Y106XKinEc6KQLn3yBIlv8TUjxaRiwq7HAL48YQwQNf03pNPh6
tXFigL4FTpORdUOUVWoE07GnSJ7qJ9C8bH/JYnU3eqQHgVLBid90ZRM2dOlEcels4cPF4ZznbAq5
lgY13bjyfoUkF2bdRkUT0daHfLxQ/dF8xiPMXDc+ApQZi7kOms7WVz/t3vZoK4mr/2eEEZKJjdTl
IZgg1j+/Z3OCRGuDrAxJCIIUyn+F31IgaZIiMsbxGjKWy5m1Hj81hchXIpieg00+aP2BFC3tO8UT
hVy9JT3ULVub4pRCTMVqVvSUwH+3x9Wt4m9YA0itfU4jq30qDX3Njx3v5x3sDkq4JTIGR+EPNno8
CfuWpgnz9Iz/TcsIfMR4PPrOvZ5PxqOk2Hs7NhytsCoChbxOVRGSOKuHvdF9wqnu34IvNA4Y0ICm
Ir1qsTIOyAQ7I74FwUvVd79AY2jsZFGo3HW7zJRQKdyaM3mlXntqTSgLSzsrKD3iF3EOKzV2nWx9
Ls7BiL+OPQyOnm95+bXTuxak+PyK88BDSg6ioKL8I/31AnCXDfsF8w1RitjQrQL77SGdBgrqJJfR
dHSSv+igg53SFx3rqSpDUc/9wUw6FDfgFf8F9swHKeooJWmAfcz4MK5OPXYzSg3Ij1Fi18nzGFmr
i6aDtInzai0TvaGQJMCPR5FgE9gn3jaIIrCYd6dyHrfFz9XoMinST841keOj+B9NqgVtdU17oc4d
kxBcJK5tYrBpbeRUQpLFBzyOiP/wifS97Gkb16/9fzXWgLvOj76xFreFqCMXo6Ne+GQBFWH5+1AU
SifxdBmHByaf+BTkeHIjgZz1Y4MtojpQrVyhqcJ3RGBXk6XEQLUXe769YGiNyUEKBezoNLM1x2RO
pfEBu4IOWBl42solDmKBDXsDVJnp5cpG9bwmNMoegeN2RMdz1ywOQb1KtMC19tKgGNjViRCdBPoV
aQtHi5uynJa+D4aA79zucvyre5qHjf/PTg2AHfir8Qu4Q04jvkAZ0xbr9r7pAfhIoT+JE3AvqxQL
go4LsmwHRmLnEjKvWQFqgeHykqQuXqwyLl0HyOHh3twLuv454sOO2SVPD9tUoxG9OxauqXQ03Kts
jH3+Uwfc5TKZ+ZOclhHtCfAzdMTVfRGNzbcyP92+p9ODWi9C+gVhFwkH4fexcb4C1P22wGL34mkd
tf3UQenaoK/sd6Jvshzs5fHfLUEHoYNibgendjsVZDrifwhah1J3UGT0vq9LnK5TDQCukyNBGRD/
PKqV/b8l3VnRH9wiIxhnOc+8B8Kl4EJNJp2Voa3jRgLH7Jgf1kbY2Mkzhe2ScRb9jLcRBAzFXMzv
Z6m2pPW7zsgyGosos86bahd/PmkIO/z1SoJdsipRBhC5X5rdXSP0ZGL1JQF2MVqA6AjXXvvYuOzj
TsdJw9JjJTf11s2Us+Z8KZCN7sg+4Y1aUz9nq1lnX6N/c3klbdvpxfUiQGxgUuI1qZvEID8ma5SA
ese9jbI7C4FNhWtaRYFF35L2uU9rpATyEYYpouNUTIeUCcArbGZ5nqm6uTYGE4swMK/a0z57+7/0
9biZMKzaWiKZrCRkAux9Lgb9iG2TEuoMMPp2K+laLDksJuYrPXf68MxzTTy6ULiY3hFWIM/9FBe+
P0hmjkdQv90NFFP0CIPPOUnbQuVajsxcCPhwHMlXGol4vSsZMhhgo0QIRXAD7Mq79NfK/7L5ZqXJ
Wkk3VyoRqugWfvZEmnDpUyDOlGrB0IzFsRAtX6zG7IB8a3jc+kwMAvyvX4z0NxKncmx+RvurhGJ8
ID5b0xIL4SDZlccL1uTUCVN0hEAU0xZiNmqTaubih6g8vMPCrFZmzcLj5/khnEce3nz3fbuWyALW
xSFRMNe4vGJFx/HBx+7d1Lq7r/g/u6MYpA2GPIr2qqu1NXiLp2PJdD/ZBrh+EZu9Ajd78VQSItf+
Ugg2w0TtzE1L+evs7JRs9MKVcpyz69oGYSthm8MBxtVrbe0yCRTpaquUeA+4+p1CmNiiH9jQoxx+
oeN6YhGRKSj3lA/ftXcenVmTsPYDKdjnozNinQeciqM+Y7I/3R8hiN+r3+N8UPZK3Vp/WtfAycIw
u72fXA4953ATgAjrDvSjpe00HvvBDs4KwoJMiCiZnSpXEqTIqURCycb6qQsnU20HU0cfpfMxSFBy
b99tN+xNPU3giiEJwKTO34TQXJH+gPUq4dvKGosZfWjDRvY7u1l7zex3SGKgf4FmrBjAvtPK0hiE
PIMLYKwORcLobNV2wzb8cVMD3UxKGn4n7GhpKalvfb4/5FOONlf0A1aSuppZpTay+zwb1HwDIih/
n5KDVwwcKFXQZnwdAu5ECxd2g6Orxry16OfSN7H22H7FlIlka80c1O9NMTkkg5MNMT0V9HRmkOyo
m3Lb4RBu1UoQNBecjOBhYUrue7bxrWYuCSn8k5MqHX2e1n40/5Mw3dh1i6Az/1q8ZmZ92wvXA327
+zymua8rFEN9QvJQbOjUDS2ZNC7/zV19sV1UcPLgxSB7nqHLMfwBRfC6TNcEu+wgcwhtvqGrQunp
WeS67nhRnYviMkfHOs2fgQcctme5ZQoF77FzkNY4+V9gggIjOfV4wXlxqplkbUimz8FZPcWaA7P/
dBw/ej1KLVMhiKQ/vbxYAHrRoGQNnnLgibusaKLsyFe77sNwq4Nd8/uKluI7aGPI2UIYiknQxJWe
Qd4psrWS4FBvOmdkpPSlEZlJbbGqbJXilouxC8n32jUe6fiPyrYvA71k34mQlra89slzL3q2D18Y
koGhvCeztHStV+5CUdI8fGn7lwCOGCoWAyozP17ja9L0E8j0Qy7QRozFeUNpTUiaf3ytfMLmRV61
0Fz9AnDTignzye+0n9oowD2NhS/lPP/qJ07JdnWBjmCwog2Jpf7Kzi9B2laOC2DvyJHTKFZq8uF8
3dVfen4kkbwd5DqugxyAf2cc/l10Z9JpP8hv7pEVt7MfU+TlQbW+8VlwuLdvII7WgOn/qlOAsqai
+AGaD0DqPtMXSBrjQe9LPNzvVEXJs9BQHV4/eXstNE02WtUNW0Ph86U6zTvU6edFimBJhmo27Ss8
bn+Ds0WBCCSjawQxLhcPGiktbNU0H4VIyGumLyh1GDKexbGnlEamCTf8Uc1i8hUNX9r0sc24FC0a
angpf4xUIdQaSNrGj8E6wCP0mph4R4coKXvogIv2OyPNhUUt7u/0LvemFuHsk/5FO/Ku735rzB5s
jGqixxKIoEBgEzjqQFEaC8KTd8tN7Vdq0qOsn8Hq7TV5goTq9zoAE/GRpBnRRBJKHa14q2drBOGk
WXR+bXOvpRVL0GMVTfQzzSk9UJMObYU1lF4U7DkLP3kUBhg48lNpmHDnS5TVgMGHkXeYpDR5Dt1S
7CPp02xwVfs7Zpgx/Y/a6cBrbplpyv16/EQZaMW2cND8We8N1udddCoFjJ8TF9tIL+xgG7NGEdU+
A13pDNa5pd2TuTGVCbyH2v3yUIa3ZmLhIYepnr3Qa5NuW3y+V4ByM/Q29uiABgc+cweDAqcAeIXq
Pl9X1A7tPmZuvTBWlYO2VXi8S/6zRu3l7577MNBYPoWuh/ntAJ+12lWWUuRKzswYoTU9uo8m/M/8
kzgXpF2+Px3lJZvGV11e9LzepNEpjuk9Y3Y/k3uqdyztt4RCQ4wqxPHVybZz1y0eEn5s/gddLvat
EV0d1X4nAPxzSCGjfkS0IWXY/g/1ItOFWyFBPIKqbh5PpRGlDk8PpL58jXWYcUI0AEGlDH7j8tQh
Cr8Scz/CtboOLg3rJpi4UL/VVog1Bl0KAxxqs889IM/RGgxbOmlu2P/6fufM6vbHiy/rLuUmSA14
4I9iXkD9JfPuWzrplkJbgLExJZs92A8tELRA1brextkV5pA7fhVX2XZ/0q9E6El/ILdIJmYUoAvF
6MHhilWbVl6xh+stkXQ3Eh5fgUnxfRTTpYYu6VfuedneFHeNZZAeHrVn/arexHr1E5TnYC5dkCC7
b4OyQqdwuz7TwyaKX7PnGFu61daERNJ4qSK9K8XGB42FY0HuuZLrtfUXbSSOclCbTqCHyEr4BrT6
2nNWrwqejXN6cXR7O6qhAd+lcbI77zyxOBaubqCy04LVAOpANGW8Lzof7F4jx8EpoHcgkm693qCb
Yg3JPMNys7gHsL18VT1lgm7Hle9xu2ETCrECbsIWIGkYPMXcrKVb83mxER/rDNr0qwbtiJgT7tZd
ldt7Sa2ZNKryHl44WNr+tCRsM8IuCHg7X3ROMYvMXF3rTeaptpDqx8PFOGu4YMtLDLIw7UqPwa2U
D7OHXLK+FE5D2IXzdA7dTPOK61MZtkQl2ArmJN7rCmEVyWWj96DZSveBtEFlYn3FU6oqg8e39TND
eV81q5Bii1S+93vVzlQ63iea63ysAB7b1ZHpadK/6u0uvqQ44M8rKMkQ01Kj/APVHlTv5/ZRu+a7
qOK8Lewu1D2uYztTR0+h7RdbZ0jXh8on7gfyfwl9ZHJGiliIL22E7Q+JIJdmTSjJYoxfiCT73cXP
VVwmUuTpq4zRMhBQRoHtfTMGqpdIUbQZxS2cu1a2/tE4Xe96Q5f4n+N/H6stPppiQwWC5rlYnOTR
5VrscUOAnbjniVQw8JRyIyADAenaiFdlKbwoAx9Smh5m4DVSpXSuawkZpbfzpTXUYNnHppttmVC8
KykIsiKVOaCA/FK6/NMzsNr2z09hvcRXAv8O8EXyNoxuH9NDiP4Y8XfgPHAiMpBvusu4L/fQW8yH
L993bRbFr1Ptr9HT6kUu9cCymY30+tekk1D2LSed2493lubZtrEhy0PAl+BQglRPlmAwX1z4Lk6s
jrvPqj2qqrD2hLQFVut1SZk2fj0qPuevvaZA7Etzk1ViTANgzTVsPGoBiF+vSbjD+o0UsdhFHHo5
0CaZH+lYX2BRqV0prUeaaGci5MGkdlLN+9UV2YpT2v0ecRK5nKvIDiV/35pyYQqybw+Quxcf5nVK
cxcrCanXfwx8SJ3BxwIefkeS6t8/N0q/0kfi13BPvDgTFaju8lfd2JEkoJUaQhq2e5V+vCrlpFWF
+M4h7jAo1V/VyvA3ITF/8+Rud3DElvlKs0xJzbAHmwoySRMfBpoSWDUrK3amprrYBxVQS34LJtUf
70nIwU1nu/3Mmm7Hr9U1RUZ29vPgu8FPzJQWahodmyUKT+QSn6IBZTDMQ8ZIQW6IuRISIF7tSOSn
CJEXVvG7SoKkRPjlpqlIN+7KiIAhLof7/EQOhPDIDMFZKYXDMMx4m4CQeom5WYjXhVNn4OMK0BVw
VuBaYGIu6B66dD6W44fuVuSy+5dBSS4rTZLnIyJghe7MXl60DAVU1kpk4yVr2TZWFe97y4c1TGYu
oH93i/+eG40MiUIqXVHe3cJefzz380PFjDMTklRL5W4+oe3rVW37S5IXa5XuG5PYQWchgyLPDp/G
Qe3H47Q1w//9zNCBcJwsUsriB/fnofaflhtwNvUoO+ecK5/EHTnTV1VEJv4W/VzFZrUT27/jSDzI
phpQ2codd2uxjWEinftvHu7Zu842Q5ft6jTLLQBJh7T7/XHZIXCMLyMkiDdVczb4Nllv6jgXYb7T
4PHMmt+eFcISD0I3WNb2c28pb4y7HXaVdHx6makRUEoJWF6l/j7lndmYO7kbV1KnaZJvukcoeAh0
YAC4HtDbJzY+GiOT/JE/JMpiexhoU2NzWtrpfaReJGqB1JMSL4McMf9zaFc0043x3tq0YPC5aGKw
JIQpBTXg2jMZvnuXDvmwSablCQF9qDdzAwD9RLgM6WMGeJkX54VlSaYamIoOdwqIUaKqwh7QywIM
B2h47jl6MzA1Sldd/QODZcqsvCtymhgkGyciJv1fDD6suqs1/jZg6tNfQ1BrDs7pBZgv9qBpIi8B
oo9/+5Zq41GNgRql0fs/+x4byU3anBCozrbcvt/EgffJuPAKcv1N4TiNTjt0pIf0CGcSuDkjEicR
5ErGXDPUNZuTmlruH6ya1/6sFAerGYfr7rTh6T1bUgRK5lkjDYEn45l3F4Zq5Uq1MM0DC9ltVRz7
YHiiGIzaaO9hx76saO531lXuYqhaH3EJQOV6VaJbidHBThiFeRhT9lgqthq12Rq+XsKiRyjrd7IM
2KmznkYp4hUJtFMYWJp5mGuAkDWUZKNeyMONva86CvBUIjlIUUshMjgWIGJlfNeE2mynybVFul9A
uPOn6QbqoVTToqu4E+Lfmh/aEbNYSI2U2OZF3svs7vO/lLrowgslPlBpiLsKrQSPCT4fco8WBozW
Q0df+xEBsjgLFp4BwckLnzTNI6O63ceZ6Bu93wcXIfkxowo9Z7jfkFz4JgrPtkzWp9Cy6IBDnfIz
BZYX+V0VsOZaBjxil28ihXH+y+074cBavbpD7zcOr81TdXEsxud1SlyrCY9XFXxEYnjq5RgNKItp
NZLU9Lh6ftjz3Yml50nDu7eKjDL4uTERJAClvklS+LmDMBypPpaVBUUF6OnqsyGOxaX44icph9qV
UK5AI0S6j0QfkVmoNwz5OxGohrDtkisPrL7ZZaMEKMkbJYFsFSwcLZQQ9ZazUcOeV2XyJgMjHp6I
vRMX8zDBSWDSwYvtcDvn3AL70FslGX+mPtfz5QTMbAYKAM0pWKWAhz39EUYzlwyVkDZktW67cD3O
gAwdj1RGfswRduxHaWb+MZEvRPIGyrW1c4xW0E6rbreoAU1USFMUmQFWw62a4tHBOJDrAkBZaWtQ
83p+9XZD4/1i7hjVoZbmU6HAjsvzLlYI1/3L3XzWNWzHmSVA7oPo2TrYojGeI9RumjswZ7SW+FNi
lgMPN7CAQq3U+Q1pFT5XkhxwXsx9bR/I4RweIek5NKAeC5FPkvjzKt4KnASUUD9PPmoDRzYp+9is
7V08GaW+0dwR6V6ZdfAfEYxeeoTTiF46RwHVcAljOFVoZ4A3cExpTqM/2bKqtdpEmrV5B0q9OQ9+
JbPpwKFiudcF3V4zgAOkCfWkun66uKcOAxwceqzYakUJg4euEQ7MXgJB5VLJ/br07KVljCctiSZf
92QQpRJ9xnwuGrxNa3IefRpkA+NlunqYNIt0CJk4rZWty5430102Fh2l4H474p6ViL0EbpqIsAZK
8UOMYneDicqPBGw4KQCfev2UNNZvGIx+lauZRXCZCz07pyTJa7f4jkvhfCfEn2v9dhCOOQ7Jcv9n
lVRU9DdyxQsIw0iaiDS8JaTT9R07MYe6t6FqVKu45W3Wgtk0FdasV4pJcROiQBlCbYmZ3zjsUyhM
sdDDRuU+IYT4U9uSCMjBPKBhlzlKckydhubyLgvWwLyObcODc3iVtrWNM4SDkC1Xm2wePzE0DD4O
eW6qJ6ShYPXl/BV/wFLvUrZwYTtb26r8PuSxavrvkLrMbGpPR9ltynQUl4en83nrFqL17JwNeV0e
GzfgVGcK8xogEBaswXYM5VQmXSXC0YNIc+T4JVVcvM/DlXNXnbAU1sO9a/UiC23EZBIKBMmLEaCy
7eTPHmJmtAp2t5agY6l5cCtZ2gv8a6drY1MaPGbjDpZCw0hlNVeTm1SKHTWkXfGxjN4g/0QPrEoH
5q19DWcXmpxaqL9dCgTAkAqFvIhVFjLfrclym3KSTdXdmb/BuWxGNWteQoKcmr6i4jCUSvYMbBX+
N2TP6EZi1C5PF5FtqKlFGmwNh35hi+HaFT8DIB3pRPgF9iDZeo77XtIobaXZcMt6sFDSfsS73Rnn
HwT+TPFxXwzS34VzEwQSOsVYZyX1VgFnxC6Vvzdo3meSnXkuIs7qYgdGuejz9djEEVxi8+vmAT2r
RbVdGvT27mrPfQp7nsne1y19N8uJfXZmxhzCsU1pD8AzaY9SVPx6MDPTeHXR/vT6up5WPRe0CJ9O
/zreWiNgFxvEpfKKKulYIY9aroL0H7BossjOYxWnRQuf1RpcNwqmedIgZ8EZTeVhhIg6j4Baz0SJ
hs7dT23rQU3r7qsqHUFWP1yiG+o8e5V8/kbsYni9Su5FRjOl3Z1JUUkGAIBPXu1sEfQP57ty0RTl
aJH/w112ii1b5k0DnAkm5UZRc8o527kVF6Wwa5umigEghQ3AW23gHMlC6lUfBJLP7T5zk3pNgyLk
jNrmCO2kKhTj/wKt4gWnBS9KwBq+gU2L85NvjqGMeKLvFAdyufIYiqX+TeuJRKNcHWNEm3MaQ/WY
P9hTEMiFUJJMjAeYWcj8JkQ+c49cmuB8/DhtMaOprBe+EnCVVrp6tcGiYN0Vv515Kivf+AdcY9zf
kgBXJayLT2/4IH28qnT/ngRHz5JTqIDKeMB7kVT1XppEAQxaR2k7igdNz+FRU8UBev8r6mNeUzki
HqZY6/4ShIg+PCjd3eeaaAZ1vyAAQ+v6QjXmPwzbJ79KiPc2b5Fsq6drUSz8FqZ6+v9QIj+GRx9Y
Iv5iEfJzLOmCoZbJWHtZsCCLZGa1sImZJBH1CAgkR0v3d6iMoKnXr4okm7omdpWytA3ZbmbpXdWt
YW47Lf/dK3DTEVMMNwE4iXgT3r9xSUDkc/nQVPZreECrEPlBAPs1lbMx5gguI853jA+WZiGBkQAs
KLbyjurQJ/23qhHojJbuzq1SiCNuUpd3Ntu7YyBl9NhwPNcd7v2HCaAKxV7BhklDdsoIs8OSAQHz
cph9/Uc00TD4MFktgzOKrRw68GY1sjWvL7Chr0vGWHZhogSN0kklJn4YbHIg3L0lPB+l82Njvyjh
uzXcIq+EcqNt1RvTbTV+FE/vocj/Inq4RZFQL+Vl00iN4otbU7bW91Dq9qnj8IZ5itFmvk7609hc
AeVdYN5fBI2Xf1mN0Ja8uBPNKb5pYmiCvibSngmhZY5GfyOf0y9JEre9q8xQVwPXvGCTnV7kHfR2
RZSa6qOK/GK+skuTi3MY35HRTr0VaLhd+9d4FEJsIzHkah+D6UCQKUEuJKD7uF3z9wu6IrGhswwq
Ub526EsNbmTMPih72PjLLdgDKja5NnuzD2iaAwZEdrmeg6yKOVHdaJv9/hwvYDL7/O0tGCDw89pO
BxMxQHVY1GK8T4Uw3T6UQeDQ0ZOClDX12S2zp1BhFc9QBbPirAYthgdaGdZOqQmcO+T4RyPkrGEX
AxGpQ0sJyh1lwZFImFhkpHiIBQppORi2G9VtB73ROfqM7vQxnk4M/46lnvud266o9yRrYfnTrpfl
dGxgLkwktttMjqRfg7UlgubYQZ504FQ+6HUN5LOuqECnaonh8DGACzEEdxiSSNg3UCsL+V3iibF+
AwbPTGa/acN8IEH5qg+iwyLnk6x+if82tHcsxWUvz1RXssFmlwA7yq+5wWqFmVdiMuRyBWqJWS4V
wQxoIrU9lkTLAKnSyeVEsKrzHFoY4IJWbQVheOZOAdcnuZHLINuaFNUCHI+xpKiR0kBRB1fhjsLE
e1mu81MvDDhtR+MV0gP3PnkAbafH6xoh2lCKUS4/KrkFgSlVOBX44rcMCbGF10O7lw4IA3vQcDAT
N4SVM9Ix8PurLPPFjb4YvYRwsj3+67ZU74NkkYW+2yXb+8As2WOGZrbeIrlduJZAFVktgb281Q9p
fRSut3qJ5olO1q27aKUolhqDrhNOJ2xfwnCVab4ozD2kVZ8VNyKPuZk7FXLSRnMgY0nGzOU1OGbZ
KAFHsiK/xty+4Un82llYE6sfpDIyeR4NXEr6mGwzvTSR6TVxTI99jLD9ZhQ/FQh79OYEw9sk5tXF
3pDth+xrLAM75DgqAQYwpqkemPQJPym6JSHHXgs5L/qVnBRCbvUpjS5ag9RXyfZLSf+qsHi2BisP
X4hPaBwtC4F4OOX9DPIhMjrR5n7881gA0fWcF4l7vQgSZt+y4X3dFx3VsIp1ETyUk8dMRwRjnq0b
ndyy35L/U5QQjqdDVPTuqC+0GEdym8HVcj3dVdPdxAvuPTHVz5uTNilxB5qHCGovE9iMvoMIpMtd
JoZPKZ5p1vXCJGWi266JqI0CQD8CpXvVgJdBtlyBdOgi87ME0lU/zT5xZ6TeN3bmurj6+ZysFJxk
y9fayOZshZh6ejIBwRUcFYvX4ZygpTSmLuC1eYZc9AtfH8+mPoFS1bwpeIzNJZp84WxsGjTTLscU
Ujy1U0iVXNM6KQsXHtOeYbqZtD04KlNm+VwgK0WbWw6H/QMFZpgimMEd5O5oO5xQCfmLLFZAQpJn
BaN6yeTMiqRsd0GKbSZtB9QsuN5PVbi0U8q+gWdRCzItFgjguWSyDE/poq/LuP3uVEnhj/kKGrcB
JXVZUPPNPo+wF0ixkW82vRPZTngS6FEuAOnu2TuCRpXK/soEIyr8AwEdZ9Bio3nLoNnNVS8a3JB8
0x0sJt9BucsdZDEVrKjRqewC6YNI7hb5Bgc8Tv3chFl1CIwBYYcPcwXu0uSy9jqawKp7fpL5tuSj
aZeh5NRvqR//XTU8DMTSNLyCdMLnz4aqAU+uh2ZsULGwdldM2QHwg2755eaGqPZ9tLdmATHclVQJ
Yun2RvAcjavHHojGGMUApmfRK3sHDJeTUhNI6rEVFT6AtKiToDGy3BXOakooXEcGKVx2O0s71f/r
LCV33z4oaHlmqn7PchumHV3zdEZ2H/tL3YLD6eEo5C+Ga9wpjGM9WMFJO76KwiPcb1KSXnZR9dbU
kPsJ6vDieVdK0H8C2dET3aHJE6k/FvQCDOLl9L4UzocN+XOn8nP14YQUj80QMj727cOsnrvrDr8R
vXSG1sYwyP+wFZWB3K7vDCE/SlowA8goSmioHIX4ZYZX0Dkmp351zHTD9NO4Hvl8TAv5hbCPO1WO
IwfZOLKW+eYrcVJ/L9Kn7HbCU7FxT9CERkn39HTDNrX6kMBdorTGvdz9umBez7Pg+9kI6IeIUW8c
iP7oxaOa3g09Xb2lLx7FkLS9GflX4UUKGVrky9xv+CwmdiYlvyQBVN9YAklLEnsNaE2JEL5JwzyS
1ALCAxAwpZeqmB7V5z00/FzyHTyMkEdqyZ0Xp973wWUoF04yA3Y/OCy/IErdo6zp+ODgj84uQHRv
/EwW5ZVjs9erG0Jc2wxXfdRb8gay93XnQADchIw6Z56oYn87fIOcPSGwHDJcj1uJzvqHH0WKUuKs
lNWXTQCI8Iy99pAm4cf2N+h4Etsj2qciKF8OycYz4tEusWdt4IOxOcx2tTKjPFMwOxIEI92byIKz
NY2X9DevOH1IBvcNHsvQUJG1euVZrEGtyvOmJ8o6Ibqr/ke4qtNwEPIFze9uUQrqXfR3CcGX6alK
jFjgUqTfkG5Khol/zfPA9pJn8uGyZbiYMkWIID32FJPR0687rCqeaE5rkJy/1NR1tr752kZ2Mi0g
SIN0IyZeC74E7wO/9D3oTtEMJ7HQEifOaTxg9Uu7YybaN+DKckYsK3A+FK5NtgtKUDqa6gt3rYui
M022mfuwr/MgUHpN+2kYJYR2vleYmxS00SNrDY9h50/Eqtxwd5fRqikOjAmqg2wO2iOOdiinHko6
R8r0i/Zygp66dCMGqQXSD0vmCJHrFdHLtTfiWTvS9G5/lvbN18HjTmX3/U1fVPi89sg64uTZD7fY
w4AW4UuiXXBVEKhFtd0+9QAB3dVFspeo2iBIlnc9PSp77aciD7IqlM0oITogEzYwAh6qEEsFxkaN
PuPZrNb6uVSIerPZaLR97mxJTq1kNjrIl1/Fa788ztasp3Rfi+EDWYtjhBKiyJHUu6YzgnUCWKZK
Gdt2gYLVZUBZwOA275Q9SKIsSZKLdSY0iu2fgRzN36bs0JoF1y/0tQKdfrPnPK69g++UHuIYHnNH
PDdlZiIUBfpy3JdS4G0xBrsgr8X70mXJBGsZT79vex6ilQ6rHAyeSrZOsM7vAsRdYyN4FA+Cbkd9
C2MdnC1sXiN9MZmRNVhS1ye5XgKQfOdt0SLpgMCbYErM/SMDo15M1LV+uRG/xeXxiamdeWQq2exP
4G8XNuh2j5hDVmh0SRdGsPf/IF+zW11oVTgcKG2njf5S9BQvFOwMbTPkr2sdwVSNShIApQmwVHmN
81v1ryRDjUqM3Qf9A11tH+gK4OaFA2tuzzyOCsWunHgdqpmg3g+Y1dRUWHIvWZTtqoj+H1vi0wOc
+V7PmyyumBrIkhQQN7xt/JtAZ3SipFv9csBsMjPrsqqkFzl06iUN4PIv5zq1UDPFd2qrk2nbj7tY
Z+3OUdzNCGvQpZTUn5d+GS3QbZsUIfz7Q0JxKs5v5JU7ylG6oCBmcXxYt3O3tbKTC6VHmjBH10w6
CesE85mYh+o3Gmw9yNu4y0jaypufGoEHuATj7he2bW5XMj76An//yycap2oUOsIzCX5QltysHz1M
XuGqCkhx4mL482iAOkzffoweADcl0mR32H6XYhNdz4aDgCq23e8IxU5xAw0dV+ur5WrDA3oeuHeu
78i2ajIV8Zulayd0fHNfUrA+Yrjw6bbEJ8/mY5vXZL7w9ycuaJt7TPLpHCVyUQh1nfs5IbYmzru3
/O8L2yUSOYMU2VzCMROloC9bF2qYxLakAZFj1UcYsSlRF9qWQSAoxUIYl4CuPFGG2Xda337XZjtD
ZlWx/q+3/z6DwSOBkoH/dC/XFFS3SZJSPElBI5FE2JZx8bY6GYOLMBRVMmfHjkDYr63Di2k1jz2J
Vp2txm7R3++rlLh1jNJCjSLxXENM83+3m0KxyMSkeoBW+sUlYvP5HswbtkoLK3IK/MGQ9ZBG0zrE
z4jtHU14UV/4NLjH+SvW0gfRl7CWn2RPGIahjKIT8oECCMnwb/BkXk1qkGCzoeSXD8Md7dcmRCC0
agO6NttwYqKlGwWRj/cGizsASdJwtDgMqFq3iEznTXEZfl+15tpLjOj7Ispi8uZdqWuNvlo/Uv1D
MlmL6ic7qWE9MNw1nC10lZl0B/kDZWsyiR9TWOye2hirOvpWSCPEUgWw0AgwsuLB4l+VY3V/nccn
clL/3hXIfHOQEwVVN3cbKZ2+vU39h1mgJGHga93i1pUAdh5FSbWnApQdOzv+VjWYcZ2M6oBofuWB
0DWxSZnj5WLOZUeX9O1IT/btWUzhHko7V81Dc9kSX80SmwFvNfkNQu3I3TgexzMxV6ofyaR3a/hV
uRVzQQ4niaaYKzO8Iet4gUtOLC6wvq6AWKyFAa7TisHQzhB9lsKKxwEgUWx9e7JHjeR3L4gjguW8
cJTS//ZGZyxbhYe1+ux8xdqFfpL8G/nLIkjaHQoAcXZGu4VZbS47488ae6HfSK7gdW7cj/WzZeVr
PhFS8oyB+Xz77XElKPp4aShOfPrADGPz8AZEhBE5dPHwWOHK/iEFld06O158MtbuQb/fkmIhqWFB
0BZktdviS8xyZSlRnV06kyJK01QrVqFZo2oBVdv+518BOajXyXmGXusPYsB/WV5bUSnlKLjlHy6+
XfV2a2F8YiQFmY+LZdzfK/VNtkMKdA0oraruP52xrMbG7oyBzv8ZcoRBz3elK/EPPdbuLWrGLQ0j
9uwdttuwXfgPVivEj50YbcnYbcjfvjFbPgUKSs7TmuOpzsvqBFhWAn/Dxv2y9gVtX9jx/ro4dPW1
SMmzaVkzC/tPVdOn+jUPzLJxm/3R8sbx/vuNruIeVg6MzvuiBAGu2/J3X4p3d7jb38NZMdfbRQzG
QPRsAxmPfVsIGPGXo4tQG4KPCu1Rxgr3WH7R3OcZ2RqLwLIsQGy1PUES5gViQVWAtfpv+dPEPfli
BhaFdC0QT7TwGkadWwPQpF7TyaVLUAP+U0YLZTbYHdUE4+iS5D4BpLvrd/XM1XRsY5MTanmYC5jD
u8vUOUO4X2PyeWDQ2P/6/KvEMtA1JqvEOkXfY1RMSMtdYW/MKx128kdBxac7Bg5eCCrBuqYq6DHw
L3lHaIbomfP93kXIcy5ZsZMI/L7zkMcrjIcoU15fNCODBDRj8C8OcaK1+7ijwas1AcGYTAwSggcU
T93mTijrBZqvAM/8eDZrTL+HIRhYyjOITUgqWpS0RF5FcsnZLYaQWrwhH4TOoAQZF43bWqOulMqL
Cl/EDrkiUlllJbOThgi339MvHs73iUJ+9VzAMH+RHoivJy5cIzIpJyNzQDa7Sm0HF8q7UMAhPIOn
G66a+FPb4/NrgxksdEj2f+txSvYdG9hMIXCcX4wgRvJ5TJYF7Y5ivz/YWV9X1558202o5FgEbMlG
zwVuiuq93TOoctf5NLEZd5cJOqnjAt/RAsS/peWNlkZOpzazuetnbLo/gFIM3WShDkCPi0oFLjNs
bHejQpQeA7xsTJveWVq0ddDXhBRi0GpBkALhh6PW5mtX/G3Hz439ZBzf77W5gi67Ze4NN927RAgX
T3ZOmG3QkS0Pl6FEcXh/KvhjH+K/OtRdDCGlPh54gSeR/eSOx90NUzCr/MxnS7VLv1V4/ehrkias
suI3Dv4+lK71KYWoEEUJ0z4InwgN9WyeZFbEz73BaqnOdp1u7mJYdwZU+yvOMiCFdoHvkQCcXD07
D5Boatr4hQW+4wOqycD4xE2icbWS9rkc+QibFIW6q2o8PuKSFboIANRMYYLf0pORWU/9701yksxz
CtwjzxgevA5ImXTamcnoCIgXBcb/VE2Kls3H0ZcEYR3n6ZSNOVeBfFGJqZ7SkM6cpHtaFvjKPuP2
H/TxgyuCVddEK6Ww694nxm8ChnuT/EUY3LX3ZiW7dZrHdhw3v03unWFWwysOcaNga6dKOe5+0V0P
sfQoc97lzB65tIOmKxhupBhi9J4VFpc3FLVA/+D1YWMAa4zmvY8vbCUl6E9qERjmDLlDbd1lH5TZ
setaekKTBiBm2P1AWKvqiB+z5HuUAwPlYfRNzOb5nM0XCzO1VsoiaO4qYTwZo3va6RMOK5h5Xtag
EN5AvTp7yz5+OyJB8CsmuWI70xBszdZ9/xkVE+Cv50zUwH2VAgy9RrZtbR8usgZcTv7x+iqjiSzv
4XTdQGzxp+8m+E3bykf4QVxWeFAA+hh0Lcmbt8SJMCFFf9gBVMnc4UN+PyrmFxr4hNZwFX/tCUap
szw6j+dv8M1MR7v0Afb1krmJ1XtwxzU5U+oOcZebysj44P5TIZ7QrRej+xWmQjFNxFuBbwRpD1q+
L3IsJwrSwlaKjYFZ/Cpq9M3tq1ytrVdmuuqj4mXXkTCUO9ho5thVU/Pc8KPyNNf658POob6mFctF
QrSL4Vc2YM50zxNPw/qCHv2HV0CXkm8VEH4bjI3ql9ifesKvGmvZfm3y5Q6Ve64qJnfikUMrogsd
wgJJ8MnEoNWX0ANB2TE4z0IgdnxTZt/HrKzSPAppr+ZkrCb4sOuFT307lmie2g/0/jFR/wXNunsV
zR+hf5qF0PxrzsWabiC54bv/RNh+oWgnSGcmSoRUFFo7ibP5M8GRRFABSpJ7COAkTpJBRxzHhqG3
1dwSfH4iZJzP+AYskvejep/AwKmXJk45+o/E8yfXHGgu5xqE+mV4eKzk4ioiFPrxdErpKT58Om80
vDtW2uctgV8hic9un7vUMTe0+L4/fon3RIsmR8W2ESATvZvbw4P67OC4aGG5docihEjtCkEVlbaN
b4cXbw/m9ay82jB+y7nhYfiSoLjKgaZCGCrNVltL9JHnB9JqU+EdMgdSt4L/LrIZbTRpF2Jl6eec
SjcCGSvV+CkexFg7YEHnT0Q3upzJWfoknl7oJwQrmSIvO/vB2cY8ZhSzySy6pLThro0bbb+RpuIx
sczceOChEqX/W/iTv9O4J1yE5urDtde2m2zVxSU3jtJz5gRG+/9n8km0faaXLaxcof4+9hQAgQrB
P0lA1YUi82dX28528rjd9IOg8QU2lk16FOZeH4SsXS72JonAYWu8fho/HfdrU8cbvhdhC44/nqiE
/+fXUc1lsGdJndXWkLFnO8JB8cBz4afHsk/NNK+M8VxylpX39RnYpcT16UH/LO/2xI2BZ49dDyVc
omIOtg5cugtfPdmDUAOZvXjMV6xC5JJKsh3AvIEGMNfR0EKz+ImbCa9ccHA7tSfTMVZ/D15gzn4p
lMEXTKWBBXVCfSr003rCjFVyHWb+AWXhMOPqzRk9Qqc+SAZ3Kg3OzoPRDo0to0ale/M8c6qoYPE1
1M9vaVPLPVUsYzh6WN62nlkV9HMtdhI+0sl7p81Bkw6g9W/eWF1AEigDGnkZIwuN7LtqBDVKDaax
52uFlgBeNpgRDkHnxmT9+HP+Jcn94QFhd9Qpls/wl0D0UtAf3KovmKC06+GLDdy3b4tsKWmwuC6X
Sr/yrxWNBDxD4ptgQM3/G6blJhr9oCw/GJTnJi9do/82uOQON55hY+P6BpmvBqPlhCJyDhJNPump
1xvBAcRwjLcpHtIv+2nH1CX7iLowzA7zEypvZWAkv8jSGNJmPITmYHilH3XQMirYzqVJx8jOFAec
eJrRSElUdbiFhkys1EABIjbppiu0JMNIhePj3xbxJoe7go+1/t5YgiAPbODnM6nfLKPQcwB2WCdQ
xnDjK1ZyctGi6EMqJ+lzkvsZ7+S5mZnHXlL9OxwJc82Pk4BgUH0+jI4BrQh81uFamtkRW2BgDXGV
PQcAMgnBlIA/nTH5+SaImBlj47ULQG83rn8dl3fFC+ismK/9/x6qV56k1JrhciiNT/6+D0e2zo+W
LRQJsBvFAtIyAvWcelArTYqAtoF+Q2mF5SDg8ueu7fVCyglhB/sfXTRg/OVSTzvBwWsEt2zbVRad
PK4jmy5DNFm3gUM/0etHhd1oufvhAoCY7EnWSmvbcvYpeH7ocgx6w3sCh38Of/v9vcn9ejL9AivM
aZLwtP8pmKGhRv84lZ8fdhfc8Ecnv4WdSMbyYdbP88TbUd2v4KwJA9JKQv3EMksXzABX9szvwmfD
fuJ9J4xDNx4Us1e8KAPI3fC7vU4F8IQjK9TkaqNHphyKmxeaF+vtigenbyeMIhOrhcH0abjybTZl
Fr6WYryKn/e3UHgdD1GCCalCVb7N9LGFmibOVJJUJKfFcsKuODfPoYPA9zQB1LAgma8+mVk4BHhc
zpXFT7CjAXJrc4/mmZhH2jfi0RsvecAr7hjr2s93A0MiQSf7CHFVyUzq6K3utUY8VYSvoSqUcLtv
YQu6n/LSX7vGBMs/OCejVXLowcbjbL4Dc1/19y2n86XfUGHd7TZibb4AVsMBgallePoT3fChZDn3
jQ838H02bMrwgFJdEDccdakhRkS+2KYsayO9tip5GEk1qXun455DppRUnhToeDoXs9QT0fqQ1Dlv
n5Vb4A6WVcaMHH+WT3yPxYd2C9kOjGWsn5E/yC9bNwIaIWWgUoj02ozSvxOihOYM4LTvQpwhSeP/
CfdgIAZ1dsXW6t1FnNSLmkYXXNhmu8VerIOKA5rvnh+v3PKOcdsvcBHr9uiTBWlBQlM3Ig+XmP5U
DU//mgMj4CexiLqQ4kRl31uy9WhNg3SLAhF+uCzP+M3fG4K8I5FaWJF127LDxYnPxKGcQxj6t2oe
mHgNtANz6XDxVQPB4wEBksN2+q3NuVojG6tqe6ZR3MS86loJV9Oc5DDux5IMV6XahyqNZrJTMaho
4MjdnauEobx4ukSxUUUnXa6Jmr6lUTaY/KYww3adB+jVkgpFQnqLQwGiSCZGE/8MKvUABkmCwYQ3
2vbM8WNrXo/HftaSCDVPoR13ngbF7E/OpoSmOH0yYPy01Q1uq+JF6VNHMMzNR1tCGMl1UCULbqAI
Cd7EIAONLMDgqbhoTvBFSEbi/qgfIv7MJyGfdO+dCiAMoykOJRsRjX/tifn3SXrnRXr2yj6TS/UX
tm2mRAQ6GcxTNklbE49AY5XDQKDck6UrQC2Jp3gpIj93Wldm7aZKWZS4S4/C/NWED2iEy/Pk4rPv
o4Eem/cqiEZQ/03sYvwWCtHM0GKhk4vWDF87OMfy54nkeDJ8EYAWSG03+M/6h0qR7IXhYZMJMwel
wR3FqhX2fp4PiDKPU4AOdh0KilFHNHNs34eTi5H/BKR3pHb5l+wEzE4dfCAbBUHwsiK1lmHzVblX
ttcj5LczG58bNQr2udO4BUCmFCwvIw/glnf6FO8hQbQ/pmYJKOTUHbzJir9/HFfF7mON7g8hTwLq
S19cACOxs+q0uJDLwSe5n37cKIB/mVEv7dqnH57RTXgS3ebRsp5S1A0O4Jhtjtnk8iy7ZOi7Mtjw
Vo8ixtJ8p0wE9UuLYxmikGMN9uUUDOIXxxH8BGLARFG2bZ3c0PCOWgM3eTVVrOmtABpMEtERT7Ts
tbPVvp2bPfaoYfFF1oNYWduqDPjzXuu+yzCtxcszdNyIV2LT29SYKf5JAQMgyP5pVuJuHKH6lFOB
QrK6/e46uf6WoW8sA64l/0EnrztTL0s59CM0SkpG+U5ZQmbNB8PTK/EFEC5cNj3hpCqPCE2ezvHM
kthFWz+WP6qi0HXq9xNiPNEhGoe1M/z+Lkmmqb83H9NmvZdavyAV5Ylpdt1xaBVN/3zub7rn1Su8
+H7t+71GbZADkMCZavB+ZrNXqC+5bVhuySjIqqOL4+hl7etMAoRIIUcVop61NAGHfhGKu/32Sd5t
sHSIIFLdPfcbOmpm7nUhYR45PEZiiG1qk/uv2UdXNSQJCXGSak5bz0V6lH5rJG+Ib6XZ8Ou88MKq
1X36NFJL0zaxh4r0tdDqQuxzx/Hq8dboDll2YAZqkhKtnMEnP7eFZWotyisWrZmIncnLFNrfs7H0
koW5nIXl3ZoxLj4tJHTdMocXe0kVRgfM6bXxmZfUzf+f7ajC+rqa/fKdF1GDjBAyp9UfeqqW4stF
Jd3dgy8m75NXsN54HmZWByraVg917OUeuGiqyedeEw2bPhuI6sd2yFdgssAoSCK3QRdQHsJgmFaW
cV97KBe80lLRwUCBZk3WZEdOF8aCju15CHQowVe+s9h1y7Qqg5Ys/4oxOmaIMn+JdH1L7MBlTU3x
d56ROq5golAPLKrMWFAHlyR/2lhr2L/EIctgxOZtFDg2CYwu0fWXU3dUzfVzPDiGooCprf9MdWvy
6WK2Xz/UuR03Y1GaPeeaLDQXe6eQCk6Wdj5LciKh3vLs8O7UCFSX0TS5f2zUxj7CglMVypnyEVXR
lsqxu6eO+Tqie4ycq1JV/Bv4V40RHg2Au1O96U1jWYAtK1Gas3KjJXAZ4UgP6/FsoMRmrEKh3GuD
LA1QyNFSHIo4ulret2xD6bOCgFlUvPEgYE6gSy1e1COn5fSKjdm0DdufRXTKjj1QaJJ7L7yekeN6
be7rrmrP6XRsiNikxFctwHOr9eJrorLmdxPMQUEA9UNU0DPnGJPTsqJ/ZRkxeEFLZ2NU1qQOO4uo
PVaqugDdD21Jv1OWo7s2q/6aPSr5xNFNLeXSAX8Cod1LOt6PEhmkn7Cj+mzQ/Y6a+E/z7xVlzooy
j5WHO+ti57+5lmqMiWCpbp3hLQ+zdou5fKG2kAawdz5Pjdy5hGB86EbGQnZl4UtUuWla5wHgRRHH
vL+EjrDbvp3DsA/W7eWMFRaM4K15gX4F5EgFJrozLdhrgR7+DMWtrhb64CkB66iw2zDvUD/lVPey
duj4lFIHjout7RjYf05e6T6pz+UtrzV2R+Vq8svKK6jFaM+z/CmCLhpS9A41LHbrpfWMEMXJ4YeX
rsfJ7ZoFdLsiaXvxC/HltFanoi06QJFHRUNzwAVpP9YdysVxZl6wxNincHqTT13yD3CVezXmVWzv
lXFVBj5NjIX1TW4Mt7+flICTLdRylRurlaKhrUqkh9t5z/k8qaujQcpt3Vy0x1aJF6sEtLbu6Ktq
1S+cXj8GREwc9rOshTSgqu4o9Op7Bg8EiMOlNA3pY+iuQfJt/OurH9PlQH2S0RJKj7bUnKnGO+LY
RlJm+DGU6GOsVOZ59aVSghVg4fmr0x5FI8JmCy5pZKpiTt2t6/3QRMxCnMoiNiGOCdv1M0yyWchr
Pype4E20XyJdIRYiE4BffajnGWVG6DxqTgfs1lMKTXpwLotGKUlawtUtI43Kfxixgfh1MlkYCwbx
gC5jJxZfr3ImZpbkj2wXXNhao9OCo7x1ia8quqZpCsmftqz4hwNxe5/RktegWjGm1mSPm6u6yf8z
v8tBmM5yeKVo3cbAoC95rDSrs4YjRfDplA0fL2CqT+L6G1+SiB5xDVCGir+wfFVlqfx0fLX8a99k
gPByMSSPZMNNBkqZ9WAtDCLO/06z9LzG3gWkj4O3dK6L/SwhhnVws4CfztWl85eH0vtdq+dGS6yE
z6Zdz0GWptCXK4n6IorMW22HH35ZC++YpzP4watrR+VRny1UnNHOAivfr3jlsk9H393SM7osnlPn
tO+GQISapTViDW/ssjP8s4swhTg1bqYn8xAiSxgbCm6kb1qlYkpX3mqwaIiXf/CqSBX2yWdxCf9o
ZVpc8lw+8IHyNpRBCdI43WavvpctZsTy+yHpEV+3B5akRQZThBq3LaqGvFG0iLOoItkZSrVLvfZt
jYYxtF5l9/lAECtNf3JKsHFmgQJx5rPMQVPyhKhm/TklbVjGxMPLB+Zkp5O0neSTVn3Cp4oBglNk
lZCsUpDue4B5UUaOG7/rA2e/83E6IlwZ/ZflM5uRw2rnLRuQlvTvRRfT027bV0kpaHM9KoWtd53o
HWGS2q5I/mxpgM75hETjJY9XyYVh1fYg/Ld/6iYlJcGDAT+J6NGmsMqg72iGqZU8nRDZHa0GJ4Dt
1rjN0s8/yzBBRdEyL0jOxQz353IJ6wsGaaf39noj/7Dbeipb4+Hhns8LQEsbMxIFh8BrRBiG3t0p
rfOObGw3xYjbirfKQ9VTZ78tmoHIARq3LZqri90n7VIu0S5DpvdR1YLnHVC82phF1OKys0Qbudri
dU6NSuh1GORBN4Wesr6+0QPtH3K051HEVTb+BwpumeWx3eO9csmGdXzjxp8H3F0XP/iXrbw16dWI
6K2olhjW4lGE/y0B+Mtt+u0Zn69EdV4+DFgBHRZEQbETOKCLTOeRH4p5j4kn/vt/BFKOo/FKoGFI
jmJEMtbf9oSWbHhQCchOtVySsTLaWF/oJTT55JbcTQdbjWLlgJpcuu/ygay2t3mb9uKyqrhPhidY
fbK0TGroVN7bqGZEQqHIOX4mhAlGb9v0TWOsMt2MuzcUwhrTn9CE82ZZ3sDtq0jYInPmW4q7lo+q
yUMK5ZCBZNUYDVIRbmLyxNTSbIAw2pf3kE2Qe6K6xaPoTL0O1gwzP9DzUhPLoUMqN0n2gH2DbIAV
9Qkq90URrPw5xBtaQ0HpmMY+M4YrFI5b8Ubf7GR1Gi3J0YPJINAoxhdNxCtqngQoFtedwrDGGM80
4os4T9I/gXci4RA0YJxouJnz2HXqM9JdYFi1xkUXL35jcpzqyzpJCNU3m0sksFJe3PatqFrPH4Fn
L7wp6XXffzEUzNC+XM4F3D6I+3rRQ/IfROF2sEEtuM0Ux2hHPnm+3aVh+OnJQIKySlAFt2PlSdX7
/5vvRLe+x4xkr3xwVuocUwHIRs3AMU61Vza/ZgtHbpz0YUqF5EaYaDfJBxqCZoYTptGngxLVNlYe
3U15xfcttqNfYb7krX5e4z5Bw5TMnUiF3eAtzCNaUDtWEi0WBCAbNJ0PwSI3AS/NXYRwbKKGvxCe
2J9b9JKGqwyG65qtzwfiOdMZUO+ijh82eFJJQHPYYfcYg1lZRASTPmx1mJLqYjvELjKpTrp1ZpjJ
XVU/c3xFZWvvzqOkOcmpQ9HwWtx/wr0vUcw9fGdK8zk6u+i/YCLn6yaDvWFUYE7Oc4lhI5QJhoNZ
9i8okDVOc4+1WY+TeClZPxBQp9r6zLM3//glin0YkC8D7qHO1VJjCln1B/GUeHETYWDyt5yefikM
mkANt5SG/UOev7yDsgf9GxeChcYEjNaylysXhnV81qxYM1ghPO4qCRNtsfEjyWOq2z7CgEzvwQSU
UXjNZacjbUMDK6GfcdRMcbvH1Gdy1wnteQCKC2vgxang36yNdnP7FxYpxGFLTvjqiC+h+4pCV2k3
fLyXorjSGuLECjvwGI8u1jEEjV04W/BTIdT0LVNwC2x8oG45ZtsBzrhytnttXRLzFgfvf4HF8f7q
U4MnINm/btgazsYazM3k2ZbCMzTL3jvOsGR7uU/PFYX/aN/mz0rchs7H2xqWYhK9D0w1wODD8Psp
79bOtW6kY0U5wwbNkaX1SHL+PvyEgLvbPPKOIxSRixBrmXDrtO770f6jmtLpnFcHFzBy/i9aTMJm
b0MFJKuaf5ZeD4aRup5LeMAdGPuOQlXmZmzVZsX7ahpQ2vlpZc3U8xYeY3IBkkdtUN2kfb67CWOs
pR+8VdLDM8bkashNe7QZVNiSrliGCVhMDHJFZWNqOb9uWKws/Zw+F+Z+9WLIQUA+fCn5hfLrFIW7
PeGM4bQvrN62tk8Q2o/vlyrzxJNjkfOFBg3dVAqnMhajuMCyls8xeDJgTFTK5Ir6xVtS5kaXWYrh
UyEO1r1nIQ2dU8bwHQlnIdCSgyHClH1W2FSAw6azqjsSJ9/Ud01q0Fy42siaXOXwcs1BLu5ufi9y
l6xXPX3Y/VhgEh8uIWOs3Ia9mGghCNMySvZCSaC3s7OgAbXoJtqU10UuSLMiPm9Fx2a7mwKvIPO0
Tk/yDwFi/GTTzLyBbVgRHEiakKwc4Htwyu6/URKCNQB3qD9inFlSVSOO3eQwefGM9E63GYDGKfSc
FteE0FkKUIi7pVnmc0+AbGIInVSUtRz0+jyhRfcSJzrT3JGMCp4RARPlf9l8qj6KRAflSpDmlc9t
9ZIMWl36cJ7wnsOzTj5rad524w1WkMK8M1NEK64XJ5PMYnGNNpfpxD4G5RQbEhARwJ6bwW+dJLDn
8zdQBoaQXVSWgsAgCIoPM0mXKRcg17XXMHHXmUzP/vEIYpb5rERSQlXJj0OyGJJ6AdpqqMud55pU
t9+98rZnA449sJAL8FrSQCvZAeJeRv4q//qZ5J2Yvr2jTMGNFjfg9dmZvc578voRigmBGtQyUzgJ
DOj6I7eK+V2Bzu2OzmTNHPzLSkQFe7stsNYw7XEvtFHrEHFRveqCpStdqp+4k1JIxIIvJDVlgJK7
Axs4wXvgO6fOBfPtapW9YO9aNFMMTQujaSmqs5rQX6uv5GHVpVC5EP68hV6dkYTWDjDNX84u4vqh
AyeCOWwrjz11tb/YQxC3G86/P6QnQNP1MJepOKepnQ4+pccmi4AzqxSfsrSiZMnH4jGZ7h95/IHS
2jnUquzPlELI/o1wvzna+L1+QeJ4vMapWJn/+Pmej/N8t/7p8cdRxaHcn/wLB+hm50XyAEtws1tY
Sjog8ABSEClzNhx1ArAiZGfzhG2+LN7khB1McIO0ciuQEy6x/cgJyA0JkSdyoFozLJav/9ZkjFXt
IlnAsyigi1ZpHYPNcj2gHhZg1JNaE8ZE9NlQNp+dIqPMUr42jA9uWpwIK8oqxtjG1NNBNYBUZuvM
+NL9jJsCkuUvaVLLK89EsWTszP/Sox3ttMNchStJKY0W2+gOCyNA/EQ+atwSG0wp1j20pWguSCaI
hawjWyh/HktApx3UYQRYq0OfdF8PJrw8PHBnMxnVLVKjlvFTMLkDCxyVoGb4n8J1t7D70MwipKtH
xM/7LFlvbOhUbI+Y8bGEU17H/B5jC9sBSge2ioV8wP1tIBm0NpVhJ0dvIwRPwHHbuosOocXHnTdY
fvK7YtVA3u5n1pWAdY4nWbDRG4y3v/hk5N3dAWSi9MNlPE1VyzTteecn6wxxUiCBuOt7gpnRFKae
jSzoszKfovc4pS98m/Von27cqgM+HbHGXI2EyBiaMf1krSg5adOHyGfQqsHrWVTV8+oyD7Mg/TK7
bW0lM3mowSUkgl2e/KtYG8UDmilerJnA3kJoMfajXbURWbBJMOR9CYnDLpcCWGFC9iJ6bt6vbiCp
e/EiqknIZj5YyarHRflsmgMOqFh/7sMLTwxpCiL53t3gksssi/yT5en00aqtEH4c88n5GNxmDMgm
j7Lbxgu3MHq8dSGxECWNOUPpPxVy4clWSgQcIJ0xzK4s0LVzjtcz38oGeBXoWTDnm1ksZ1epuWG0
RTdjtOXsQ+GmvsruOMjgUCmdG/6M0186T7TTpgI3aFFap365SY7/mVApM5SJerdgchruce9CvMWj
8xDC8cZF9EzXnAQMK3I5haufNIlvNYCHQBnzTzNjn21xISQcXz1SEsNvILnE1CU7/d3E6iOUpDFr
kQKsCrWCw6/gWzPNo+UcKCaUp5ddF/HX6WbY1jM0XtzomWsKRspnYvdYc/2VWM9a3/IagJuyCTkd
ehjN/Sm8gJ3OhL90vxgywRjtvcK5S+Ugwk6THOjQnQ5e1Lbyb+MzkO89m/ACdpLsSwT3/z5vuiWB
yawCynnXxb8djteigqqUm6Lkpqe4T1Z3dktwPmSqb8nHCV3uzZXOp2ASStolceXF5g49aUQwy4dr
2ASundtnSXqa9GCUccXHkZbyrBn6ivqFMo/iBmpE4tUas6x0A0hb/iYmTuLKR/8s5S3U7RBoCPCM
39m/OQkzXTCESqW0EynHN5VNxpFmgk34a5UPXcac82wcaW4a9MNYQz8K2EfYFdHi1NRFginYjXtw
4ZdXhzyzXZOsNWnyAlE1KPjCRocylwvxxlJeKeD9TDlVpS5S6loTZ/wnl68SFEuYoE/094ue3Yp0
WX1iHX/OMl3zVgH2LC3inOU0iNSmOIs5yphjofa30qsk4uXX3AY2wQTRDY1MSCGhqkyKtQVomswr
62cyKUXpuKwWfR3qyyXYmsV7tIhGK7SG8Iejdu+pd/L1JJeCK/9FnxfaBHyqD0fyloYt2ye+q9/R
PLve6/6GGPK5hT1qjABtwok2VtUJ6K9m6Gb4kUMMYYL2HXH+JYTO6Ig2ezDVPqii5RjcNpsbFNzp
0cvpVhu8FKDEh4Zf8PLR3Fe394y7mO5C+USHZ+/34X5Dsg20YYzwBtAWG4MxbFo2fYuDW43hu8BS
bnBF1sDXY4YGvnEBLfVouhylsiA5ClFRd0Y6Ue88nOQmR2JiLQyUvNhp8QRxQl1FZUmhI6maSCay
uy26qD0gIqg5PQmj/latpGJXX2AfCXpoeIBifeBvnNSsh/zpPrKQvbdUxSswjeslpf7H6q9MGXdW
hSMJNxi86F+DJxiO7MIssP2HJkybzuNmtrqwpQLUqLzhj7lr3uVLUDSUB8MxiWIhQKymBDpwLDJn
Rn1Z4pWncLTzhmM+qNhtlRKmQb/hsk0ItcqhhW8Eh8zHyaAYk8+Lw9h4YdBRDKDIxo67nkRVRIs7
LQq4FgUZupK0x+TIrYUtMcQingnVwo7ILTDlRJA4bGBxDULHHJxO5I88zMeeMzu3FI/lP0jMJdfW
ToBJE63bmkWM/sF+Zbpf/jPAmHuc2vLXD6KpMK6pjA8Iy+rAERJUz1H1c6gr26Y4FLqquk4GMEcs
RDbJ0VllkPscKnSI9PFeynQr6NT/zCSn7aASbkF6DpOYvgplThkDqvk0DVOlTmJkJUA2mbmyj1sk
QzvPi3Mss3E8ca1j4zhvSHQAGtp6Ukxg5cOpVKRsEY3V+un/TqchIvSKtdebJS7JEOlxn6JuHoSq
g68UlA8xu8s5Xfg9N7k9i+d74R/BNBU1OgKViMbveY3jGF0Yt86pq84jaHJEDfJVt6t9rdOoLXQ7
0si7+GJr5TDtAm9VCzELeaC6Mn5g1Cyj8Cj9lDtj4wvAReKIu84Jit8igQK1T6InQTZXE+lqMH5A
Bfa75rEzzJXMha55hm9wOocOCPHnIMi5iuC2fVcSiQs8glGeKhwxrAMwxS0l6bqCjuIZv6SEAs7h
Od3QyE/NAITNGREI1wndQczcdeuD8PJbFHthLIChPeOySdy54FyZH088mjQwBnWhliFQuyIX9Qqf
FjhWXDLSJVDK/TKABDsEZbZlh4gabUL0wIkKBmk6FvlM86K5TNSVEtgwLIwGwclJfVrDzF69jZJf
el3l98JwBHrLG8KCFKqnDCXmhq06i3jx8oO9CUD+VX70Lza3Vz0C/x+RxzGEZ5Ao0K9W5JpGMBHC
utqqTvaiEitAGvyWy+zKC73MwxFrZZw3tM+dGpQtKt1IYebD5tpyoF96GjzkDj4HajBVYh8mknvC
kfbpFjuMKljg8xaO/h/YA6O5iDMSgLP2WK25YvCGK+/DjGYLaI6t9DG+8nDq1x8HW+75amp0uRjB
TNlCGdrMOvUdCPqSSq6BOmrk6lBblE80p2QukFoRZePlhiU38zskET5HsrR0agLeUgnsQK821TyP
+1Vxv9OIQpbYzgenPE2ZRSKsPziPpgobJHO33VaHqEZhDtIgYt4FTO+fEy2wDtUuvyG4EA2AB1q9
EpkewIKC0pbgRqKOvewBBBNfFevqcV9A4+DKEom+EeoHhH/citC705r0oPzO8EeMsX+w23OZzeCz
NUuiYJW+K+emELB7Eehm/LukgHJaNb2MXD/YSyY2MU34sOm6dVfOCClmpBUgecRHiGLhEycsiuPJ
hFMWJy0FiSBqInnLUd/iNFJQuTV6xQSAWC2AMRsdNg/Kz5JnvZ6FAnVWIzEeAuWv7d6JkwnluHAS
2JjH52F/v5XL9Hi85jhWzZYTjB9b+D3MBJz5cHElsOF8j9GIEug5p+09VISFkeVistfhNrGfaU78
Bd8oftLBveDTFhgtcEperPJM94c6kUtX/rNDypQHX7krwiM4Ljv3VDL8kyYY8cF3FXrAK2sSJozl
WX5CLyZg5SJuYGSH0E556dMMVZpAn9U0RbZnBL90u8uLHhXRnIb+jBadN+svxw+RVZTIvAJ2w/d0
8lMMVyV3QRnHpsVyVc3PMoWuZjOg/qDarzK4bHLmqLYPf1EkOVP7YgaqbA+ImIb9HKlcuEeuFqrR
OzHcB2YPuwYXP31dr7CdjlWPnaHqjdRj5KTaHCn8S4CxDRXDOaDuhd0wvX7yOMyQNw9ygBU8/ZUz
bHzFhChyhJg+tsozrrU/QiLJmdbqR064u6M+MGPQ4a7EERlNln1t45LtMS60eudvSESTnuAYg0sC
iIsz9FrZxLtvwk24hScUY7ys4m75VwWA0Rwu52I7S36pEBf90FrK85Ob7drHzpBK1HhlHFMRLxc1
xM4fxbZHOBra7WDdxOQnKS608+bLliD5bYv3wCc4BAwXIEEMZbF+/uHf1l9I+wssMQKvCw9jK8o3
76lWGcOe+OcnYdMpJNnX5QkrCh+TNMSYIrY4OGmD4+bBae+DftYnpGZsvej7/l0t60dOiclTulc4
+DeenQMV8YctH5E2Zv9aI6hj4vfaTzxfF0QPhAbzCsUpUMpB2m4RFzo1xIBFiPAqG7ByXqaE4fRg
mnNPm+DaYzixW57KwlFKD+7dEquLz4YiIN8mKvhNbed+zalLYAy1hCmpf0t8RhY++wteJa7ixmQQ
Sj3dnWZo7eiNan/Ns33nJyrH7M/yy1LvFsetAgZDXylJMCSOh6wxJY9IYPdnBQf9+FoooXT/7VgS
QLb21HLtXjqz3Q7ozWilKnBjsJXcC/gZf+Rdsf5liZpjxDHHvbFRCPIgSoekgiyrWGr40okw0T3Q
/Fr4Mww/TWtFlJ6QuYWrMPi3D97Ju/asY0SSa4bjzpBAOv2IJPHPGM37C1ZZRkDlbITQASR0FRlM
wT5irEDMJfq1Y8Sc9Dr0tsbA+v+R/tsTnk1zbphPzfRYjKSBWgdJYhoLxs3jL1hRBAm8fcSo5aKy
pWSFao0U+4JL30ueVnk6kYHUS/Gjoxt4zuVo+tI4iKNjksY/w6RSqg9k8sj9pq2Mv/WZng0NEDtL
raFcnpsytjFkAdBFRncKZIkYecJZfbP86w4ILbeZI6MDO+O9ylmGuSbjRCZUCPgn7p5nS7evmkj5
yFLK8lnhSHbAR4Tq4Jwu6tzogVR28p+cePZYPECLneE9WG8lw8reW3E7xzX/Znmczn/lZ2QlJsoa
NjB9quGqbTA19iKgVR+JJhVOJjL0oeiMCnLBAKYoKB/LcuhjOec6NJrxpLbjNSNZxtLtiN7AWxxF
TDNQeaGhahO4D10oWVOrlp1wwKrCFNDBBCBlPAk/tm77MWOQRYfdB7I2E+IL92FajyrSa8WpfejH
0GlFBsN2E/50PZkH6+aFFeGpFop4+zpulavs8J4ENFPfkvG87lMaczJinEA3bRSKvNU3aqvQcJDx
HsFWOyv4dsKOY44ALyFcBCk7mM05b4NNFH3vuFHsChjPZv1ireJ8umZlM8x2jmpEbTeDX3e50xby
0JE/YlM24A3KuObFKtBM5hbvicjAvRX9rkkgZ6+k0SdG7UPS68hmMgogkA8pbJzV9TagsmArntEs
3WlwjDazRiFEe4UFvmHFoH36bjoUL5DGkdgpX4auyW8mz03BXGs1/hNcLL6wJFnI6JraK0eR5U07
q4IyeNrunG2xeEVzAuHYUYEdIMtaJ8UrJH6rpfofG6LuuWBnTGRMEskjjQFyF90OBb4ibK/4K68t
cAxXP9q3Pb/LBZlG/krHB54CxOfYyyaEjBsOjjEoX9KqVNtLI2oEN0dSeK/SaXTsIDv9nIygaSky
YuQAPk5olzG2O5nqmf9IR0HrZyD4IK+s49QjmeCKCksaf954RWjoz3/spuzJ3x7o/5DLqYLWH02t
BWgZN7oULFYNVISjR1gRoZIVfzaWhMaLNfOg8p6FPn1dV4l22Kf9sb74Asw41+m0gwvRrw0YJRk3
QulatFMHxGuORWCm5SxPwgbYYb7Inicda79ZdKDdBl2Ma1IOUeX/45IhSiwwZFuhdn2OlknuJUpZ
y6Q/ROAwLcIMjBEV8LWBCaJDKzcDP5UdbORuy9LPEga6haQ6dyucb2cgJBgnb1omgZEB107ypuZo
dqMGteOiDJyFFsBvFQV1ytZXSVokA5Exz2wFxC317u4sWQAtrMrZqcSA+swQv7JXQo+4wL7bd3ZX
EhwEJMRJC8D4u29ZBn31DlGxR+SHVbA7ZLzHVtyUuDFCbx5JodEBaunxeEAsTj/f/qwiayrDUHTq
gbTgQQgX+SnaT1FQntMU+BxYaU5frdevJBoBY77QhZDwt9LWv8S+V473sbD7dWUi0hw+aIBF8/kM
sO2t2DCQ+2nMMRiAtYgqufoXtUvRTbqP5nsh+fjOmLB9eXWrqVdoPBNxXsUgW8i4bMV+ncRF7CUM
N3RB/8LWuHy4F0EwbXaN/pFIpHtRdU7c4gb9P4g+ksQ89Hx8KdLDu1rc9btFZ16zoWx5c0cQIqNU
Yi/gerxdi6mP+/+PG81nBJeADyJwXmBgO095L4a610C7g+HqE6Si7DplEa09w5jHDYvyNEwqEBD4
39EeJjUWj1uI6WITB3T2L35aXvP1NwD0GCZ+VwFg5b1LkpnbSjP/oOIyFpYdpy9S5wSnWBdBfYP3
FPsIeRMyIid8nRC3ocdbKNKT9lVDaWiy2/Gxpturg7h1ZDh0B+hrVTmuRYDdtUmWGhf0Tnc/BGVl
YyZl4AzLXKFRJrjji+w5YzQglkU4mRIq2TcQ2xAvCFG1nyJL56vSE3FAmJGeYhfzzmnS1OrS5bIR
BrWuXU+ztCY3HVS2z0TTnlS0smJZ7KacEbz2vNnv6gYrGroWN34fVBXmnNVjq5TqU7/sLJfrrQpl
/lBUuJpUhlzFyF6Bt+jBdrOmb5zgB2mm4ydwOx/DEwWnPmSoPJCFo86q8YTCWYNo0vt9ipJjmufd
GUtWztnm67we5INCCJ2nUqUPrnVQ4Zxw0VWXLHHwE2RxmSdwCJzIyDwfExhSSIhkx1UTS9p1MN/S
69FPP5QA2irGTiFwNazbfa97nqfaj8OuHqiYvHEbPcO7rkwAFf1VLa18Ej+EzHeOx5rJfwpT3jm+
8vicES1KsFm8hLvkBjatreV1irCmmOa/SwN6PS41LciGGNss5h7Oky01IZfg1gjHCQaMHVKurPqI
aM+XXPytxCoXGK+WbrrsQDLZOb4zY/AuMGMlNUoyNNqh1s9IoiK9bCzaOMGWKTKjT7M41xqXw3M5
f50Gk2vSwzzlJiDaS95uHYlgo0Zjq/Tn735dHO8Z+hGRV711vEr96Pewpqed+XM723n5HtjJMZJK
qB756YbkzXxxMehVgQeQhWaUR8uT4Nd5cjeQpQGshiodItBFYGpsKzmiBpp/4Zsv6IPweQeE/cE9
nmpkkCafLaOoMkNhzQyCEKp03lR6+COeXeXlBqAQPTEu27sgBn+QtYTDN0BTmFaApV08kDHbCMWQ
+QhxeEJ39lxCAUNAuVTsQn8BE6J8pQT2dK8ZOxIkZAA0ieNAfvj6YE3ukOdODZKe81dic+XW7h+e
YccJlzCWLBcAjI4mFzINNWeiiH4o1CJR46SRkEHilcCIHQkPgFFILmlqjQtZFX6URYEveybLAhs4
DNouKU4I3tPzhSmY4jnvIF8kLlbBKThcMhWUC3MSlbnhsghx0RV1RDiefu0ICD+k4Kl5PtCqnZFB
/E6BUww/oi/PZsA0kZI5O1VuKJHayOQrec7ECQ1rTYO/p68V37Qz39ZiRSYhFnHMKdHQ2Cxu5iG3
xQR4pGnI8tYrMvtPfaMkaELYKBsPF8U8yBnJBVoERDSFeDa2nqxk1aq1LoD6GvkasikzeeCynWx0
R37e69z+Gck8WmRAnPPEV5gdqfns7Yo2k4HUBgumiW3rYy9y4XsS/z/GM8S04+uEtbuyq0UnfSZK
zgGWoUIP9ogFNq0DhQVjnM7G7Ity9wioj/QKz+qFK5OsKNxzr43GRqsnel0S8MF7EHi4j2mkn8zk
aZNyGQOseDguj3RmOI5WknBtGL6T7/8YTLMGIVHl4VCarxrf+nVguo8jJJHz9EE7vSWLsXLZwoj4
aS28A07vuWsouTS8VZbNlcEk7Vsd5UrH8WOzJ//34ETf4aOVr7OkYBzym4X0JMuAPy90cc61fxxo
dyjCO9ibhGKsB7ROyScBJi+jhH16BPjmSlcXIv/MMSP8XFctr/ld1H06R25slx+thrpcSIBc1f21
0Y5apZ4XZUTllpyziKBtY+3dIt12iJbKcHhSpLh7UtF1Dh2R2yGo2ouAjUtvclPkH1mRjA1zU/7i
1LuyWBNUP+Y/0S22VgbcQlk68pb+IpJSPPUeohFPrTVMu4DCPX8RjbPC6CkVR1rccCiwXL+K0HIm
JBrW28cq4CVSFL7ME3D9cZ6MqZ4s8pTxm2+Asr/up8MlRdp6LFdyjhFlNXq3CZtM/XgqoR0hRV5Q
h3aezNDjU/w7FEXlNxJPeUc/CZru1TJBW3KX9zX0CTcqeeGQrjPlmcY4ycSEI6mG4lVSXvm441Wn
//Ptkmx4xiFTt1ZiSI62NzAcYwuThqWGREqzPaMga8pFL/U9e8I8qAnHuV3QnYFqiCObbX9LcmVy
ENwKVJVqZpR0UV6PeUXQzCRc7MRJcTBGejH5FEkhdfXbc2NjmXqV0nPeKWbQ16hKtW4eMV8t2jq8
PSBNlODKUxE68sQdOPSX1eN7vmwbJoXiZFTnwl89ilYbUVS75sAu81lxMhcxgAqCF1807ZnEG7xy
zmWKNJ6Od22Mn3h3RKa7JOXlBbCosoAsJQlSLrP6GkDL6CgcArgspMXBsCcAxbWsNX052Lpp30ve
C1ls5STuCjugdLRXAs8gz3fWYqUaplck8RhnhpSJNIp+7lb3BYEx12xxg+BujEBZ5t9BmDVEvXTv
MHfeG9lJa3FcwUys6m97EO4TjsSZd8veCaUB78AXoykIk1ZBUIDHOIshAPN+f6nOrzyf4TqT4wPN
49fgjr+v/ZYVO36AYtWRQnQlNVeReW21MDapWXibt+YAuTAIHEclxzdWyJ02lmbxeMNMnWRCe6pm
Fhu1yfulK3dOCC9RnXpLU2HsxX34pNZy0b941K9UdmEhm9HvNz8hHPAchKjoNgDZhvRUzoAKpz3l
EhI18UPrkoXedTCynZFCMZ2eGIITDBacbP3pTWoBBLJy0LNJ5T2li0BSLF49eqlofAOvjLfezlbH
xwgSvlwZWdZPF9yd8LVRjj7R9P12uwnN0uy4AyiqSwO1PkTBGvd0k7k6o0rk8nK9cgijJrz8zgy2
bny43euzIw0eHA0Wz5LQytwPRqwcdG30KQ7bobT1xr7W+h0Wf+kE54MRB4vwMn5yVJLjn3krjDTk
KYnkrbSVvN5QNWu/R3/I3x/fzeJXhoDq3i3QrqwDUE52voBDk9lV+Yn6CTQqJEKW5n2dknNHehaX
+VRb3mnUiBV7CXDrhg/xOsPx8AJLF+uiJEZo+7ep03L1AVUw7JXHOa3khTaFVC4N5Iq4VbIP1xj5
APSvNICJIC1OH1jD/8tnAQOpw7Cs/Pb3wA90300xCw7aT0trq1QPrkETG8fsERBfJyxip4vB5GRP
iX281IB9J/E0fnRPeF3YqjtjuenhHkW13REgj/inFwhiXjiNoCnSxaUAwcfQ2PNUrXk5QwRFFQMC
frg+XZqQFtsmGuz/SpRY6gx50fh6lnvXhgSiwsTeyFGztDeSkq83wK5OmFIZ0dE3MnxzGMi5oUnZ
H9lnMWyYsLAvTgRLCBJiMtICpHKTzfe0FDkUbQCMRPDch7z1nDKi5ZqzNBgGD8TWpuE3hZNmz3fO
FV9d8xTsoUbGdREPU1vdrzl7mY6lE3Efg3WcIVAkiAHi3yRQEl0xFBHBizHi470HCbD4PgP4tB5i
+miJlMQQPLsmxqc+sR8EeJFPTgPIiLLeXC1KlY1Y+8az1m+/oAoshXxH97H+WPPZn7B3M5nVtIeU
VqBsH6wEjJwObU2K1igZSDiNLOfbHMwgvZPNuplIo5NKb1wE6WmLTxAy47ag+FoPDar99UnnYAJB
K8KQHaLyF7tDp85nzcCnI9jAsLccg2fR4ZFcD1t/xgCLbpjOUt358dBk+LmGf17iAlPoYMPJ+9ml
L/aYZYpFNmCyTgpjf07OWGHhCGfI6VxCbnbsYOfRXXh0fkaSLuBlIpv46fN+NnQCbJ20liXqr+Ti
o9wSrJbECw0SBr+0AZVf9s88QXqdhlCrt0jc8s9xTCDvQUa43k2ObZw2fKVpBiboPVjMq9tGRo/X
aLtGMeIU8rfdjIHIszK0ormJdg3PFXacsNGWTLdJc24qE/yvguqrrkvpHbasBIrRtTdsGPlWyU7Y
Um7JlDqLfkiLhzg3WdSa6lVwp9G3XI0bzWkNhFPI6rglhZGdsOMGkWWL4V3yXNNYCx7yBNAjW3TZ
tsUgRbRvpIXan04sm9PVENaeqLMqROdse19tKn8paNOYB0zTFVyLz4HtPxStFyHuENCEAur0LGCb
24PzH4SyvAIqKhQOJHNG0TOpjOrkTTsN0pSL/qx4dsFBxCg6QYfB0IItPdLI3jK6jfpp7HVORFj+
U+yZGYOLeRdWXzWx6LvIelT2pvwUCDhoZIabOo2FQt2SvTNIc1+9M+i05gqatly5sgGGs7hiVKnN
DAAac44W2iJW1FS8q52whkfmEuxCG9n322ASYlqhwcuvVctTV2g25ht2ZGeD58gynMqiIe5CHajX
gPkBkHozf61ou7wwfAcXWNwe3mfyXcxrrj6bYRcid09a66K/c+TQNlpYZGAmBzpzU+mtZcFeEc2C
V+gayQGPqKzXk8WwagE9gefzREaxlzpko3UsuJCt6VXUdBaq7CvfoCv6CrPx/xXXTLBwgKE6JKRk
x1Sv7gaBYNEQbV7e/m8HNOoEcae+d8wE74GJMdPa2UlMUrXlOsmJtYOVOfrZyja4+NgjJIlg2zhu
SpHvMTGkVFpzZK5Wu6I08nXlzF9jKNoNeoXCH5ZXkB4n1EDjIjqm6SZ+gcsAlp8wS6i5bBZiXOQ9
IGDmmkRXJ1p3by4oVbF2z8E0w9IAyM4sc/azDz8EbEBKni7UDaG5Tn8gJ5dbG6vjiVNjZIEno/Ak
zG8DxlI9OqYPfziVTChDKxAeWVE9dWc3l/0h5SIbYcVRAg9bBev0XtF3BGhs3fsMFm6UziSDygre
FoPX8vy0TA61LTMXHHVTTbjeB67mhIsNvdxna7a3uGySGcRASqu72RX7D+/mktXuZf9h6V2uRSOH
yvpMQgH57Xpn6nQiN0e4S7cli1yfWF3O2i3z7TCf4kG85VvgIGoXl8BdPSeD4uQ9ubORTK8jYCx/
QYp7vtAmbKv3VlgNHxJOCX0cP7ryMpYOcyt/+DKOfamRNW+zVcU0LYGhRYYgDrGutK2vKevEGmN6
u8ITEQbuyMbh7+VYMD5Keyf9lZNoD+Trh+LkoKBlKDt7gQjL/eBRitmZ+iwBAlU1k1kTC2qeXoj0
TUOSacIoZJgkD9+3h3J17+5fNLSAgLMnRcq24TOrBvzRsILEwr5wtHev8RAvMEvVaMQoBaGUWS9I
6GYCQ6kDfxaRbBJQUbsOEMKis2G2kTXn8bdI8P9vi/6efU7FafzsjeQi8tTPkN8J8Abnk0d1VP1S
zG9c0hlShEbfQLw/p4ULamddBYf6BmGgXFv6DISc7H/kZWUECL+/ZrK5aJlPU1MF3q4DRYEeG/yL
KWoO8pAOfcW073GwaOGetRKOSiXt7ROFZrD1ncPf8B906uQzkKFWuPg5BKuhkIjQdpnOLX+zUWz0
Nrl2GJsZ3OQRj+kHWvqjrmHY2Yky61Ehe5jyAwMCRS945o3PnBzrVwHMl7Paov/hcZOakIZQ13Em
Xg1LG3UaePMi4Jl/InOJfH3v+CvxfEp8rI0zxQ8FbqtawU0vxRj3kpV6tJVNygL900uriT1FtMmg
iJGiZ+CrFKD445jILfWIeb68eJiaU524TLfc/Txs2AUiEsSsuSV1pY67y8hwY7nloabBs4U40oIS
dqhXiBHrrfkoOLcuB6Lt0M3PayOc8xXB4Oi5SRnUQW4FOuZutpsJHx0k3mxjg0lbMnwIB/HcFbpy
2ejvYuiTy717m/2Ga+iSFU29CtDR2w+WTcMffbzh4CART8Fjenzmh6+p5mM39xqa95A3UMROcMSI
hy3r9iCeONBFvsYLPwuh7mZ/i6UvBAQK1W2PLbNBdqJsKg+klEyeYYQvL2VimxrJlw5IX2UNn7YU
Gb6QKgtl72+9qQpa5sBWDpCGXx9SYA9eLNfV6oreQ8tej+xr8Bc+7V2G/xwssoQiY75aDnMJCT69
iQBrWRou1OVooKEReIJX0tO6avkhFRKN74d2Q9fPQLtNKd5SLJMlZcqydAzad3IlA1B7npmLS/KI
4L3kBm1SO/PB26RgwBlKiER8Wb2pgHwa141d4ap0m6eCFiEKlG6WK6DGn2WF0i0GjSYAstrzDeXi
/+TKgdYaaWirAS+3onfIsMUl6FceoLOFmOroyVa4fex+/HTtM/JumPBVhPxpzy01Oeuv9DpAF9Je
9g2L51NBv6P1TFpSv0dE0QyQSqn0eYQru05zo//xaNh07f36kB7o+71qioT66vteB4zLUtRzOXuQ
slv0vXnX7i6Ou9fyqpll+l7rO222SxRdV5v+9DoXqchMaXMCKG3zQ++QhxJavm7uLHrlIlnHeYfl
BK/fJbJgGnn81rsbY5vWWjPegW94Du8L369zHnrIrzm54mzC2EQ16/z5LSVHZgQFrgP1zlrApK6s
92ysw+1bSBHgrSkxwANdT1iY9JlToytiZBwXgcfiOIJjlFx/RSv9on0XhQTyzjJf7nxhKdL57b5x
5shS1TGkiguw3NPE4n0+wQVJgO3WdVregBLVMeU0iK+IInopjJ5nYWXw1T+fM7wDnu8joFNNGI0u
6RPLTdo2tLihZAaSUq4iroArplT0ikX2J8eFdMTRnsVZLhSsGNBkNq95erdGDaAtXoD1dXD3RYZj
9mmKabkU3/5CyBr7T9Vk2TpzJIWKvoAlJf8AieHSq/g3SFyOqLftbdwy5Kwep6Qkb4bh3ZiuDot+
lB18lBIb8KHZnIKaw8m7Idhu2C/n9PCLn7w2XUuM09xfmQj3L07d+8Qgka8tQB+QxoXf7JhlmSpw
nH07mLzyDC2h1bnMaEMOKYpeyIyGmN51R7iJsneNFbCMoih+eimiL8enwoTJBqKzAXJ0sypxGYLp
QBqeC1+o0C6C+NLvQOhY7KKU6kbDf7KDM5a/WG5efwlk021bGpI5xxnGB2hi1DY9x2BdQI38zHZu
xUOlVyxArv0Rn6JW/ZlDjj99e40+6vCfKn5NFMbRzUqqO5nXRSsxkmv4azncY/AI1DOipEy+jSRx
djb2Bx11FpYW7I6UADDh03A88+kbcKuNj9W7uzMQvZU13KcYlgPOOTFqTc7mvQ+GYRKO4FAKOqIl
rJSl97kEfUKUCg7qjozCWIu7OUZHcukr0w9AuETRiIUqkgaOXWSe2mKnlyKJD3QXFvK28gom1hzB
Um9sjQ04BkfKE69YliRuifkc19Dxa9tpzyo/MM+ONQPVVoe9jankADJLaviA6IuxCU+W/rwJe5qA
E3zm2iR9a/1zKNavFuGoZRHuQqsebexLqHID3mUOZsCwJI8zOIjxTNj6Havj/l4p+uykndo4/82U
SOs52c9gh5UhSHjvpuFSgaN7ndZkxFYq3iK/QqiTr+ec0jjVR7/AIpVchkJpmOThDV7wB910Sg96
FMcWXzq2W87au2fo+1dTMw11zI/2Q6zQXtOKk6jSPGB+OCE1uIDY0IMlJW7vu9vtdWygzpoL4h3o
E2+JCQG6fYRyOqgoKDq2jFuub/vTRJSpZor8Pl1G938OVmWBAapYa8DfMKHKE5jFTT93zB/wOKIH
OWW1fhm/ievG4mTBjrYp9CzTfuLTyzgWocYfZmWY6t/kdZcuKhHxcXg24iktPteZf0jtF3juHTv1
R0AqR4s3hNswoS1xm0+cztjQ7/kcBEwAyPdt5vIiDueswx0NaNBGpnH355do6V4mgK6NEq8HVXBt
HK7/WhNx8EDcIU6YgFERZs0IJJlcx400WV68PfUxYtptGMLc34v9ujIhZ0X9AfWFEbb1khdNWeeK
wjLYIAuLRVgS0svhQEJFp08Zdu+Rgf9m3lbiM7wF0PP1+RGnwavhtqhoiAUjwdvN+xqbXYVIZzQG
m3t/FEJdjytk5+b4hoVafxdYMNviaY556vWO3Ktlg7wY5O8wz6t4Tf1nvD2PVA38KMDlpMeXu8lf
fBHRDsSdaA8bfisaR1KLzGrag0jr752Tin2W5JfxGRwcYJvcdkS6ZkKRnGjaxrn6j8oAwHovoJd6
Ktxb9HnjAtv/0hdFMsglkweGMX5NkkgMLHV9GmmUrYt5KAxno222OQ+3rUrmMzq+m44MdVScLikD
Jw05xL3gqzNmZ9KBA3C7htXaGXtdAAGMIOd24mPZaDbBR+4KCi/4ArBBOFHUIVFZSkHK5wav2vD6
JiZ0rbrl57GK2z2DspEAfOrH3ezObDgp0rIag7a28Rrl79hEBpqQAt7uAAdzi76+0vSrG4ySt6qE
vbN+gaJnBg0iiDFDPwGi3a7rcFRwTlV22ADvH51CqpoDX0uWi/7rm/wBVX8R6dfg+nT4m+c+gjLZ
cPuCe6WDSvnDn6bAi6i0fawpRz9zljHM8rRlfApxmMv1OUvrC9EmFznD8nHpqjaaJM44wkABcWZC
7PW7URDpMr1fcsC5yHJfrtm4jNVNeSf2wldKUSeF11glsV3yBIHotyXUCl6ZpaeqMjuKF5b4hIlV
0KbMK7ocgs3U2Br5aBFVj1sNpdhTYWLx9BmoNnmUw4PM8iWAvtu/Mic8ZoOUpL+4YAa5gfKMoSGH
G63eJnMmnQYitwGgCnZVhjl6HPrAOy0vh0Cgz3CB3rmwsSwcV/jYANd1e7VbUP+tqBdUkJefR2L5
SGyLgtKqCD+V4QUoT339hoZorP/xyXs5umJo5VpVLyw41Zg1czIYqlw5tkyjGQ0ySwqM6TqrzwsU
FAQYCQpKgSknVWfl6cXnRLbHyfYOdaXvPcb7YIv74At3sOs8z4NO5mNhxqorF5uZYWEsU5Seswe8
IqInzDZoz5km54rtFZv3X4Bxlpihhpwu7R98xz+IP6kEL5w11RHPXOI9NetlXbu3z8tyJ/I4aDu6
UT+SFKRgweKHhQVx3tJyGXN3WIQf5Q8fXbfR0nbsNBcVv/Ku9qJRXzVhjB09/W3+zqXzb3jJKeV9
rtFKGJXs7rvnhyz7yCVFdpkrrgW3P+A49XJo0x7foIh/lsKXzOjFjwzoVW8N4ESz96yAc7lY+zXl
Z/T12bXyDrehb6igfhHeqeOX8hs+ThPo2Sj7jMxrulUJwOzsyYNtG+Roat31KOnvM8LSinXMZ7kN
eE81CjdxRSk/p/vNDK+hKTeg15EANVI+oJ+PA3wFs50h25Nps7lI6IL14oPUH4K9xFzuMEWnQIkq
kTl0zasr0jIdX3UYb2PxLok7WbEcpcDqRlcUx90Srt0B8WLe0Wz18QrzwkEdqyCMaoC++U7WsRNB
ENgKeJIXP/onU6iybz8oiy0rWHw7ZwNUP9lu0b/kdzdpsZG2R7SCPFMm0q924Rzyc1IDpRAMUEVM
CB2n/RLVKwfLLvbj8Bs71lhvA9Ff48wAJG+yFBlmQ9uTMU7HP7tQxTyVKQODv3eFjdPIkQqwe84Q
1qFRpu+qRXCmqU4CVx3QiDZOZAWqvznP6ra1FRI+h+xcqNRh77RkLBq18IW4IyaXmN3eofP3+dwg
m0LI2w7yNp5rvfJn2v2ZA8wiQjYc3pcqqt0agNqvbddkT1kNZ8w3JjcopxGACtuC/v+F8BnqlJgY
LZyeRH2q5Wv5iCiPjvVTL6Yndybl7TlGxlLXFh1G9bXnHI8JWOvgyKPpZ4Q8tkZcBRtbYyFve7yf
W3lLmZYo5zOxUptci9Ah/JS2IMchxu4AJJnGcNWrB1M2u4phPiqgbqvsOOL57OvMUW7QUJGu13cH
/eXKnAJXdOjVZ7uuwh0TJfTeCb6MLaI8zQgXC52tbhnS8zSrzlVnLfboP4W+xoRVRovAVu83xdQw
7+A8fLBgOHrlulOl9aa15Ms68jt6h1BQ2aDf/tVoanX4YRpWbxgqEldkeHL4DoKNEaPGQz8p+6SU
Jvzc4GRIBH98sak9yy4HkLIO2pGbw6mhKYeCQUlCSMgIvgJBa3s1SWGxIURyZDG7KqKlInuSBZTv
p/s2meReuk1EbnblBZ5rVntvmIWE7JViZUmwcEEZIBrvJ87b1n+HcZfV4/ipDtesiDrA/OURyv4+
uP7dZbbz27SAUmROmjzv8efgyCqx3bU5OQx0e2iBhFOIEUWCbmTLyYD9bFDUMi41LaCnpsxsY7hf
yt0IAJDTsSz+Vg9jU0ds20NpXKm3hzidxyO44vzhMVKtPn1FEG623eqgp6kPrfmIBIXjSxNZ937K
0pmY+tvNR+KlmEJeUy84AjA7UX/BPMHKOOfzVKE6pdZuTpGgSfCtxQFSXqYcq3td4Tpw2VYilEUR
JSWqfEqUbG1hOCPo4oUvM23SAl2oO1NABbnHgFXdXO7tiVz2CifQwTgQnaa4p1OtSzd9sYIg+XyS
lVRuYt/yc4X8CI1ztJVXFPeueaDD3Z7Eht9i06MVUjLfGHrfp+91juAHr/2D6BChQQpcQcWPJ6ZM
3AV0gGVEQqQs/16VG+W3x+U+GZ7GMJq6/1JwUyQwNq73m18cPEpce+4Xvd0s9nhCK0A452tfSF8b
3FLDX1KhCiWTbtHX9k0PjcDA1hg61yzVzRDYs5Z3dHwvBtwc9eI5sHvszR0w2SkErVXmW465ZELA
4FkvPxXz/hM2tNfvdl29yUTXzxT0tNqvt4FtV2KlHodz0PsJ2JVz559SngtW66loEPtLxRb42D42
mjiJ5PVPJMH/iuJZQxq6GoEK+VfEyPXI6bZfDnWWKuekdekp7g6ahIYYuPCwoTC81pU8Sd4jg4FY
/huX+6sEQ9B5xiZj47hGWz+qCqkxl19DNNQ12TnUYJlyseBciADnoMYpClmfPTe0DdVJb5H3mpCN
VRKo/aizVnecNY9zX8nuKsUlS9bBK0Dgg9QLi9CJNoKACL5F3Uw6p+YaxypkGZsUUUNw3gWGlaAE
Ft5u0wsvK5EUi2dfmVndUs7nAZZ3ExTBwSduBAUT5btTdaLYQclYBpbrO9CAGzEDJKG5JNIWactJ
GNsyzr2dY7vo60P469BPeQj9eEQI3jCw69WvwIQ2cZr2WlzCcbN464ttnWBhch/DYi4FH14neBzg
EkpX7k84m+e5Wa9Y9iHQJ1UtE6xjomF7gZ9t725JkPFUOOecWxo98ntL3EHV7aM6Th6AuolitCUB
+2f27G0rdwlPzNkhMyswMk/Ot0pPphi9HF2GeWs9X5XmxOeDN6pw4CUvHpdQlUCYVWbo3S0dwkhz
eX+NMxhf2acKWMOlal0RrLqiJUm8CaIFMTlnvLOQorAWNYm2fD7P4upa0sjNSFqFW4nSXKFfNFD+
ULg5fqfLY7tdmGTo50x4hBDZkzCw2K+YpeMAcr1B9CgALeRYkqcA6sQzBfKkaelKlaeBEi/4kGo1
efm3ZkZGaTl6wfVfHiz15tlQIDrHxi0QjhKlcdLj3krctOAnIHc8llj1oQ591Tj/a/BThLm74kuv
oZv9/4gvqhCGs/uNLhcRVCqovUBwOZJDN9OAQU/5njzf7ITy6HTSXTqsPvRNfu5xD5wClykvDVVe
t20/ZNBfxLf9B/NOU8HchvsgyqbMlrLsILX7UDRBL4m4Oo/ig8oE99WydswdzQT1nBkAYmqlkqgm
x8a6GeuBqeEDrmG1VGNxwc7wwm32c6aw7Mqa2wr1kzcQDvSSTsiHCM0TPnZks8IazgAKoheOTYJ/
gzAqQY6B9V4gBxUdaKBAkTLPDKrNupQdKagBEZxRFz8cx/fcxbXR7gf5LP49shRMiYQQSdJJ65FI
yfqfwg5fSt0+oNhPzkwI2MRjsJBuDA5/9oxR1bqUd3c1MZDfpLOGiufh4D+kI0Tgliah2KC4HFv+
Y9ZyPpRJ9FyGv+m8hsa0LUyECKY9LA3EyRmhoG6UxTxmb6LMm9ucP/l1zvfH7W9vPIPXu3pi/wak
3qexz/TISR4LhLBL3kKahHYbplpIglk1OJiSaNV4jgvjMbpPOHfkW2lLW6sgfBJ1YolmV72oBQ3G
D3zIMhO+A0LytULuL5YLNo2JblR6DwnPM9EV0Bt3HVutkokvAUsUXjURQfZ9xKWluX3rTh+yBL7f
M1hJMEEinGDw+3gyu90gnf2nfsCCtW/NI1Cd3zzSB/E6f4OTwjNUIBGrYiDV+uADaZ2cOmFaGUEu
FmV1hkQA5k1ji+wMyWu0nVHCM/AoWGf6OydM8Tqf1hsjyLMJfpC5JO4XJH7TP3H5DxBYZhRTvYAC
N1L7TnCdTpUC1CU+fyb17dDg/OQi1Gou8BJlqum8Wy6mDx9lzG/GJWfrv6xtVPjF4GTJZITFCOCt
04qvf7WdFwfUyWjCCkd9d3GYKqubZlzgaQqfXc6XxU9lCTeDLJWkTDKxt2GdKOJiHYQx+YGuB3Id
ozxOJW1kv9pYutthY35U8CAEo8mIaeWa54lnyoigAg/WWvD++4k0mFXlAov9+aM/+ETsHpa46436
+zfDhkvAWX5BAmk+CFJKgmoqmV8EjeBvEwCkld7Ke9gNdPy9KUTEny4Vi9kJfGIxNQwe357uzL6r
dXy4FvkdfOU19dDNkraFecP3IbRnT7mWMwdT984LcN1S619wzKqF1zNMInn6xvA+asHgIYL4NlW6
S5sDnii2aJix1GPsxQdQJ1+uCoTlomHMsiyO+H4E2gHRnc5I694njaP3uRIzwvcXCxFa4tDIfdwM
ueWpjJ1upekZpyvxcne3XjryHYivhRHmTzdahk4qHjYQEs/MUzVltrBtYKcMO66sLRYCwzOfvMOE
KtHfeb8tbyZpBiUBvTOVzYbIWYxO0uzGTNjUwGZ4413OWAodz5TxYn89kuebvHwrdH41ZNuStGSh
hnsPxNVq8ede4Y8FVWzBrG2w6oAIaNF1X1fMpPKw8JCp2v5TzuF4jUzLYb/ovZURuEVwSyCAAFhs
q5XI2xGlidTsRRScBF7t0mr7+dVkD635TM92XRFlO8e3dVAi6sqGgd3j5RtZG5m6ElqUCH40+Nq2
erOvI4JSOxXEt13AFReEVKfoc408MTkd2lQqt/uBLtUeID1UuFS4hQY4cjY2jYPUmN5md3QKIFzI
upf8KT7JDvPerbEbNSy3Zw8lYMDgO5eRWYgFdZ0Swrt9R/BkednT8KSgI/ndNB4ywb/UVEBbHFhZ
MJFFUOAI+vj/UjtF7YqvYWPPDX5DLF+lT7crQqlY8XFjeuEF0RuVixEsmVV5rBbqw8OtszLyCPT6
xYVO6eSVR7rdKmVhhGL7YkIoR7ZoWiTFpVZi0W8GUT2CySvB41AXQk9dIj07ypAkNh9Ya/lGWAHv
i5fwy+lws28+fw9JePY6JXnymmHodgqNXop18iMGisTdmvgbRrhanKga7ItCcWnlkNed4V3hNDcW
8Mt4hNMF4VCNWkyys6Zuq1zjNnb1hsS9/8fYc5x9OqJVoOBlNvOvIc8WlYTNNUkVjCfU5wnvZLpo
/xYu6AQ/D1b8VEUh4itXT2LVQ/Nxvh11Se+9EVEsxFCQz2gjHdCRp//fcc5OROsZSYl1EgU9cFqM
7Jxa7Zibg6KASL5YSIeQCvGcRI5Opa3/EtCdwmTuGyGZnTOjjsgWJNvr3H8EI5rrPf08BPX7QRdN
O6X5PDPNd66Xhy6xC80gMg80fC5BoqDEpxQeyfSdQN6+qsmLYO8S9DhqlsfgN3iNIHRy2Fnsl9QY
1d+ko855CYCopj70R0BPfO9n0wb/ASOVaLKhRcSELd/Aes2vP/7N1RfB77ugmK31TYSEqozg6xrG
80ERvctLBxMqwBGwWEIoR/HeOwF9g5Pog4kZXcYu+i6kEMeIuYSAoGlfsehBTCbwsE/AOBpkx+1Z
NiALh8zOa2sZJhhkDXqoz0ziQB5lRrLXBSZRITjxc4MO/XbZlpuQz7KNIXI2Oj3hLaZ9Tc8GzmSj
1ctLbUzji9csfU9m0oi7HSsLwl13GDy1O2YRJZ9AyOThTXTEQbHOV3NReqT5JZdj8VtANLN0iFlb
01RIh9+xVfzauTcHFbTseu430M15OE0KDgshDKMRs5BlOlXIJrvQqiCX0apOcTQGcbjCUx7vsyt0
yf9BSdK3IfzZiZFqvtFfqPF5AYAUce7+i/1GLXbAhUCcXK5iHumeKqeQl2EgjQ6jjfz09LeNU/cD
f8gibB6CBMyc6N+1em/AXAw2Kq5b3dn9fDzAmYOn09iGCB9PJD1sH+NHqwMz//5OPCFdYw4DZ0Nu
5kYcFqzbR1amn7OP2Rd5KE50NJe4thUV8n1+gUAS9b20uXsITKH171/7H640S6+gTvtykn/MRaP1
Rkd0kkpcq1OPm7ioQQXMFpMN2007BsT0n4H8amo4OjhWY0AvqIWEKPTLw4vTbfMCWzw2Yh413YE8
XTY9+lDtP2N+LBvo9qEfOJx9i2566j6qDpI55IewXT9y6j7XFnTaXBBduscDbU8YQKevg2plNIZq
SHvD+SoqD0/8Q5cQ0AS12pZ/KiuOOyef51t0awduyZ6UPQ8ITx9HP1NtdNQvvwUuJ08WgEdo+MA5
Xn1DfyfT+2J+dByHizB3w3EtIFYtGRQUIEx7HK56IY3wE1u87oUtYQIDOd6Nn76C3fRJt+mIhKHD
4i6nprCCO1zNTZ5/5hmBVxmiMUmS6in1DdYIx6gX0hKX9xk2RYy7HTrfm3btZTXuAoFC2mRxIu6e
AsaZpXkXUtnVOABZCoByCBG6TbmzGDwnQYcxZjM0xmJVY45DsaratKWXbtYKCENCIA30mykcv2NP
bll+p7e1dfLSKYJqW5Tq5EqbjnzkNpV5ne4C6ybsJcDbzt3CwGGh25muyJCyeqYIejZiwIyxlNx+
IGOmEvBI7PLpyQzWDN8BipkcuXXWRCzs+3znA/huy862e2bXbgnn2MJEOk7qvGv4nLc+NEDC5yL8
q01cVyFqSs7dzD7oj1/ZtoyD7/HgW7Ne92sCvNoA1dWfSbpJxTZl8oqlTs48vV3T+kRhabGr3k2c
/oEoH6G2EOEjjqldFCfjXoSWhjR2tC97FGp/sx6AE6EsRXOw8UFmBJ/+NqH+M4hInEEhAMUTmFnt
vo7xCNV8DaLgC/VxR7Jxp6kW3PCNINg6FAdfcJRlC0CT+aQQP/0+sAUk7MtJYx4/Qq+TYWjeR5EP
MGw5GYWVJYHHseO3IKhKNxrYYqC+tVlEuDh4Ci0tpFw/XWFlHxor5eVIg5epu/HT0DYcKJEmuFg/
DrmLCQRLavJ2Eet/ZN3GxDHjtyFdKAJzMbMv9QG6lA+dj3VrTgYefqudJFdy5U01oWxE3ETpF91r
YSd9RzFHN7REF+jgqTJU5gFq7DL7qPnjULXByV84Dw+cHG7Lml1wfwMaWA0giESeGDmOMi5pcDsy
F+s0ECdPX9L5AbTYXVF4NfQSrK661BcZHz6PscMN5P+ILeDXa53SmC7OuV2UlhNA1NpyD6NB4E3P
2I+XxpaYHaQ1rnwutd1N88LVIzNAWKrcBzdW5MYTkJED7fWaKvHOxw9h+0thwbC85Ge49Iwh9yJT
zXP/l9hn89mIB8xpQdixnRzvVF9zxt4nl99ZtX7e55Zmy47Vj+Cb6MVlHHZDunBeIBoORmZmyC5n
wCJxDfnAxbIT+zQqSUIfx5zBMO5oNMVeIQ6Uy5qKr2cSx4yx3O3fEQ6KiT/9ZNgKReS5TUFuqJyh
E6vWKFc+lUM336n8kZUHaScFUokP6ovSgUF6bPa6R8cNSL2sMNXpG1QKuKYioDdCwL4IkxnZmusE
YLOxXU+GxsadIqyWMkzmKgw8Ai0um4szm1QAipqR0j4NmMZRyOtqdlWlcd5qQY7Z9e0Itr2oO9xP
SKMfl81+3TUTkCdNy7QrD3bqMJonezfeQseQGsns7mklHRKRs4YT/1dAMYyyg9vqZM7uguoqzSp8
rzfqVqXZn0zcN73cBcxATvWd+iuikrrluMqET8T6P5Scm62Y4HmXlimllvIw8g3VpUn4tBFkPB4O
isOHfzfY4hTgHFdOUYtaK9hI/cpzNdeIA7mmSLGT88HRvDt+Zq3NQyBKhiBsPYjwPclQ8/Ox4BjC
1Vx9dhJCTS/W3WH1Vv+zpb1D07PsMvFQitKxGmmGPTfHKUZJuiKmVVN9m0kOOcet2Rc8r8+XNynH
d6hVCNBqVEHebTKZZva+8oXj9QJo6rnGrn4g7FafNGg49bK1CD0OhNfYJPrg4JN3sNm0HVAu4uBV
5Kq8rGwlwMUr4bAP2ohlEmb/u6orYNimu+ULcmeiTvELWDyW4MA2K059r/Fwa0i0Kk5Rsqw65GTg
lc3G6UQB5lZxtR5xWDJj0qYeZGDLOkkzOjgUufhoEerqIspQC4QnNsqYNRgaN3tJWOIT5b1RC+7B
YCiMMJY0KB5QIL0X1punIepbFsCNKI74JD2qAvQLeFRclCJMoGFxaXDrWarYiLT1KYbDtPbLObdG
TcGf4Rxeby9lNDJQcTA01RIOeEfLib6XZR8bAfpyYEqYZdne1c+cysYEt2X9w8znjjk+HdRMXjc5
+n+WAvQHx1Lstv6f3w9aUASVXg7lkGWeb1Yl5VXvsCyn2bo6ENjOottj3sx1u0PbAzlSNAvlOQFZ
2qrg4BwtaX6irmBNDlYbR6Y6YJAN61LTjrOIsq2JhcpJBUiHZUyf+OQ78WmTapXss2QC4iKVfd6V
PXHuBgez+AvXvPTAnAJIT0xWRWWf9nlDTa7eh9a3Bp+Z9Mv6Z5glG3J6j3kKNMVZEZDMdkqPqRx8
FrhijIxYoOYyVyOC20gn0wCiE1h1soqHPIy8sEv2+filPEFfLOZaw2Z4X9jl3e5zHi3UzozWAwF5
fA+VN43cGvsk2+JWI9GX2qzgOKduRuUN+imJZGOZqyPtVaDQY2Pt+4fhFcX919Df5uaMhY2c02pj
GRzgHB7E50iEBWHHt9lQnhXT2QX0Ew+vs+EUlWeenVXx0naClLzvHJFsIxpg1h28FTJLbN3wcNyk
GEfiiavuek+mS2KDhd+2K8/R7+T7Y62rIRwCxFSVZ5+sXLZaVo0jfFYqij/cGbhuHAkqmXzjxgBO
vDflRm6VsCicGtyT4sUiuaiAPQwaEXwU0+9z6yr9iNpGTszyeS61nhurUVjs/PCtGhtuvJSngaVo
DYuGegy+KdwPd98GYI/E1DQUSrpnPWkTr1iaA+0giQTZPtO2aHpD5ii+W3x6csQ8KLOD10YjvX7J
JAxMHgmNknKDMyyUWCqaMfdWyZdJ2u2Q3pFAHmw8YRDNxYZWSCNFSyK07M7RXGO1ZJFXz0JZ65WH
PaC6fjVuMltJgJ2j+1nsrq0SOIWBvG+H5skZQfoES+JNK+siom4a/JHWNoxG7V5RJfVVUXAfxZrk
6zauuQCAFAoqF+MarSRc4nUgQEqWHEJxjbp13nnf3ek8yT7WsIXjqjb0ZNBBd77wmd78Z8ePWU/M
pOyaSIug5tpmG8vvWesjk/KsyUiNb/RMr3YhIii3cLtogBngh0tHZRR09wWISvjk2ZN/0Gdi+DnD
8rer372KrdKcc0PacsWIu5ZGePo6Wq7UU9yXQPbe46E1Q3B5LbTTUOSZXWsOf5Y+qQcHnWYuYOsv
pWwp0Rv715kWkFL/2gNQWI/RtG9X061AUP+lCfeAakLYb2OFup0m9oOdvnYLXEFpQCJb5sC6fU4O
LCCwz4flTX8PFr2sbfeTFJqTSXjTfVR1GQnvi+e7pRKTYJpnuIsdTkXR7/sLgb6cGWiUTzTcVGG+
JSpSkVRKurieMe6NF6wAB4zlOzq1AY14L6MNl0Pqkcz/udViO/hLMtoWFU6Ks2UeWCAUjLDakgb0
NeLQPdoyTgpevUhkzA2m4DB5nS6HXKdtc6z2BSYBHtTZ6BAJyaKsywKKib0hdLpkQuA2t6WG4Ei5
CpVv8m98Q9gXpBl5zJ2Q07rH8GY0hQSjw+lOIDXG6F8dHpDxgZfmOT9j0B0eyggRi4w9zyLoNiDY
IglhXnQcv/+TJjcibu4kb2U802QVe2KU6l8SwHlEcl9ZRBJWhiiMKlwShkZx8P3XgZXjWunZO7E1
oXKQIbI2J6D8uE0RAkA5irOvd2x2GJI1UT1G87ukibo+W5Xd8WayYNp4cmHQy3t0xqLt7QnnTHah
pAAdH1l0YRp+y4BWW4uQTQ1aKRgs+Afhhafaj8/brHOwzXPBhJXeLRmOnWFxC3GG6PhSoZiLn2hl
MLwZ2r6j3A/lZMKI7TFDb1K+Mp3aYXxeKmecoEcn8QcQEy0tthK4+FULRg+St6rFzA6GCggOURYT
ftRzak1G3HFT63+UhD9wURJNg/ZnhdJQh4VJqnYSXHw2DjEAOPHC2MpdJDBDUr4+QUxUnQNEa6iN
n+dmqjlnd57mOSXwxbH/u81T1btJzFJp96qbClWUSBiZvhBR7cwE6OFGdKLEmmoNXXUL5HF881Me
nz0NFCpKCZfv5paPW9jIKM6nKyFyNVLMFO7LCPhh1RCGOAjjUUIuIXblONe4/p7jWZHslxQ+0IuP
vNfSmgSgMbkGOCuC1juQ+6GcTySbg1Zs+CeMoNSSlx17lxfHGrv/UdmX6SdPZ4pcBViMBF+Evr79
rtYasJR4I0dWLV/T0xyACgB1hFEuh6QLWrJVQM0pFQjXpyjKEc3h9DGXAMYxzC2Rzc9/l/+t3lg8
XK6h3kVGxlyeMU3lMZIPVwO50hYkFCxASImVy1OMnH9XTFZgm+U4YufT+EHhf6yDXlW7ACMh6OWQ
O2gYgSdQyTjKxvR1mhyxeyocGEY94IPXUXxwtcXjQRY2cdg/BNWIs5oAi6BvHJSu6nSeorcVrLBc
TYkogHDxj00mbiWed1Hy/m+6Zk6VZbnhm7QIPofasqY4WmaDIlufbHmE4P0p+9+co89NGBpNFQ/p
fxpLgZTyyJD5rS9tu844pmURbZXNIIkjyAQ1XmJ6xSJZMVaJKeiI+E2tQKgyvGTc1QKfglUhhbjT
oJDybVHGER9ge3c/hQO/X17CY2B45/qbNm8mMIHG5kSuD4qa+fRBxgZPMjAuu7U1BIK4bn7HgvuS
SEbAINhdxQ2X4fpDHgUgUv3gD1jQO9qvUu6byZmXG1UXhh3URXl3deF0TNj1sCddN2TpgTWhYjBO
Bg3h1a/fhDtK0zLiief50ahFQ6Nd/qvuqEBSdv8KfLHofXJjOp0hpfM2xpMaH02ckCIgcyKVlc3N
r6PAtpyCBkq+vDU5FfLJQ565LNL5wQ/KHiAnm7g4eOD1ygJoVO5GSayGXTNCbAKK3HF1KmGfKUgy
IQWDno38Euzks87omr6ChMK4HVSpQDay9BMi2O9E22y6D3QKidB5IKtCqrxLkj8Xre8kTC1PTdIr
judQvmLvyXFzoopdYdnO+pehG2iSlv9snlSfuGBPwL7jYblPe/JCDQltnarMr5Q1xVLx4yH5IQ+8
YDpjYb3IDIvlZhzmq+UO5u3E2kQzbJSE6XnrTj+bATyP3X5eT6WgI+mNssg0LLTZBk7MO+KhrWjX
Jcxa05BlaQvBPaw3ae98A5SEz0nktKXrLJ8ci7EzAZQJuC5QTM2g33nx3GxispRuqTeGMJJKI58L
uZ78N63e/1nL6soYsr8YERRICbC7e5fQt5nvGXgCZU5zk0FhSqwQ5DQpTf0iV+P/hKks8222c+ts
b1naCKuOM2k4tnCNu0FNws0sPcSD8RMFRUawPsRv+rPrfqqYvqbRj8hqVKpTpm6M7Y6Vmr8pXuWm
FhYTFLPF9hJOvRy0TKwwo2CZFz6aVIPM3ijUHgWGQQXiWNEjNoRWtG8bKZn2PX+Fs7tTjrWc4P9G
e1oC0IM1pmilj1m4G4qqGiO2x6NDcSJ+6n4acCSjfnUespohe7drAQHuXAC3DDfnrQnRfBRvn6WR
kKbfDpeCe1LMKMLJw+yudBbTksh9hD/Tp6PdrzVPPNyIv5ULqmQJlqXdONsedJYQIYOSmXte4+un
UQqT0fkj826O8Hk4NoaLoBBgiSj+tHJRY4ZinaVUI4FFLSowpyMKm8XB3+viO5194fGD8RQ88lHH
xiLov8vaZ2XliGG0IlklkUYQTL89VUFwHc0UvfSi/0DzZ0+zKMETsXHb3bOhB5Acid07O1xjN0mP
EOBn3BH5zloYTFQvPBsXn6uqxuBosjFpObDzHGRI70YTWbcVcV8Gu+YiLrT7L9CaioE8tlwxXZJy
uiyfhe+/WigJohTFZMDAc/gBuUszSor9b2gTw5Xhugj9KCsJ+MLYMwMoagcW6RSOArLF9czU69Sa
2Sg96frOEOnq3BVzpjOGDsbpyUswbLPXfINev2LupzUYkH0wfcT6sC2WyuKVIA1Aw4SrE+AiU84I
HuXT4JQmHcMU41m3YykqHmWX34ZZrttrRJfzsMPvmnbXbRSZBzLQIbLlC/lB7VOQ6fmuxfeYGCJO
2YZIoep8FerCu8HGKeD2usik+ZvfEEb56K1OIXFA6GBtlS0Qypv2KLB6pKKQwfLi84S9a4CU3HU7
HaDSD4xp07SV3ONCI0Xz9G1xvcEz1udUYkA2qtd5n+j2gHfeqCXx0eKVC1bhLx6ZA3iGD4wEDYXi
B3NFoZH+ZaxH4Kqs5IZbxlPjgdfVic3Ve7Fmh9wPr2RSrhMctdQySgfVdgvEpYwrZ4fTC1M4+XVR
dxA7Fpeppv8nKhnbqlxZw1c56HduMfkFjK4eMKrfTZl7NFD8CXwUfj2Z/8FoGJG0stONv/e67W+s
bhrx/sKks+j6Mo6NFjoyfEJEzt6x84IruzvvyGUT6wNy4wjrI7BYJDzt6d+OA0fhDacZZoOkswf4
iC11hiAuxA1+wBNWr0S00Ui4ecYA/uH+n/aOcUGhObjHXTv4dhEcgK9z6bRjdqK6ITBw06fx84ZY
I8qCxWDOLSupP10fTAK9CXvoAKdpB7JBxOMkNpPuAq1+vQQLL+pMJKRrcip8JxFnHpwd17nFLxey
AiGVFkVfGRcBjaCurVSWTIZYFh5g9MxUBIGfNNcJrE3MfrpHIsmvtf+mDR9CCjT+2jCl2Zw7sNy4
/izi3C47yq2huu+xyWjM5iyCDgXfSE/ULote3UKfYXqnTcMnNglUhnLQ8LvGdF6D7T4JoTTTbRjq
RKFRrtsTSh4p83Hc70CSAcP9xkz99R0MddS8Bi+fSgs50WiRzs3nhJKyyK96gQOZ1GI65K9XF4Kk
U8a+o6lMFjv32UJrSJ3MtPammcFxQW674K+nFYW3N94Uh1AlvTa6YZENebdgMu3j82pMkf4vsH4r
4jDyoD8fKdfqx2Vj6gpABq1dum7ST+TBixl7FOQGWSVTeevluycQutvXm+a9iQrNslO2uJDj+ScL
joNg0w+ULjxQKY9GwubZtnZVxMF2sh9JgSRvFM14WMxFz+mqjIXVIAwshWh1zt86BhApwCuSIdUc
l67TlC/u/qoVwxWhPONFvEXdnMQushRx9Ibm6R39GVPMIihydO9coS8TBxNkDJ1oXAxrl8slWGxg
7Ae1tgxHsRj6nbS3VwmbXJUIxTNw19mViTzldyQsKqAABWAx8VVd+A+oHq1mgdvlInHHgjaHesO/
cTVxcPQJrFkJpXEBZkJVpupwI/E5Nd2Tf7V4DKZH1hBEVzpUlffv8n3maj7cVkfafXklk/X5gH9p
csx479YyaT+7KQz8f+1HHKt1Ps3vbAa+hNcQPAoCaSUTIgp+//a4KRA6zBtJZtzfsBM0L88HTfOh
Cmd+GeLPNXovbvl4QbHsC/F2nuPzZp9c2mCeK9icp0oXfF2uagohNKshFhF1VTAXQb0+tHm49tgc
C6SiTWhufxhAdYkEPFUFgzUeFkHNNZlXcccPJByrY269KaLjlfRW9pYmVaUGAIH8BjdFattnl44A
LV9LiRKwdh12B1hBk9fQG9MIQCuzLUzIaRk/kY9flD6eu+j4+ob/sReKK5iDqNMPoTHkqLr3IBBg
jIIgf8cSK9FaCshIHNYUN+pBZsBMeqoEEdu715fl7mHHGZ+b9FtMcu7bRZSW7ah36Y+OcTWpnkmz
tAjwfIZ0Tw9r7qwj7iQeZWXOHX+7XVclF9vsE3rlx0MZ5TVY2ynuTxS1l8jsfK5Mta88JnKjCzbx
Mar+/c19hWQZdcMs8aEHi0UYMzPfmLGH7bJhyKeNqArUpJ3ADaU46HWleppADd8qpPkOItYVHmzN
QtNz/DwCUvf8MAj/wcU/f1Pjz8AKboza7Z1Mpe+X84nB7pm1/a2qfs9/7frO0xofOdVkQZmDOTRN
J0693wDYfAd1dF1eJr2EFxA6jTaaHCHvc8aw8lVc4sy8sVoX/kEMTJ6TTOVR/mt54531jjIZwjpa
7fIW/s7bXdQ9WTgtAQAKKvzvSOoKGxYTkYJcwBvkW/cYz/+4lqB3LU9FYsoSdS8VuuYtMVuBfyJR
X0+BIB7Zb+ASogleaGqpkWqjcgfcaMgwBfQdbyCUzv9sXWDjM+jyFBEof7Z9TLW5cFc/oMqPVXP7
LON5bNyNJBwVvBwC4wPsFnY6uDn+bDndnwnm7SD7vRphRFhOkAp4yNsyFsnJlFoZw2NazKL1LoEY
DFMn4yr07xnwrFITdopXO7UbeIA6sDMfgO2fMx2S2e7DyvoDds4xqjsqnuIVtqtYCKHwql9RycGl
+EBEl3sZQI0rn4cP1puCFQuSyUYppghFngDm+Wu7H2h+0MAWkhIaGchaSTM6mpKjaOT0LszM2VNn
HyfBuB0Fsugz0vTDwtrL5VMIaJUKj14Nq90WQiwPJObEB0nH4Zf2nc0woQdvjRGcnIETtBK0wI61
nv6qc3NalfM5oKZrq6gYP7SP0tABY5TYCFw+4O6/lFJgp+Nqx4KGD9sMFmNymce/RU7ESjdeIOpr
t2kWJHLCW9F6C+Gsg2sRi2QU58WE/v73/gIWR4K9h8xc1kqeiG7Y3lTCH5aJaU9xpThbVZqg9y48
6t3pD+u+BTdoE8kZK8pzdhNdjpU7aFXOK6ulDYHWNnneZj0hpX3RUkBWVEW1L5nAzUvns8l9Af1z
Ktj0R4v92IZQI14XGh1KkEsjIk36AwwRDz4+rrJ/6kg54VC/p3DfI669jwsUJMTf+o7tRdlU7sxS
9FAh/Qu/CJgyeIZMJ4tQHcJNCI8Qi3yQYXHHJ3Rr1tFlZgrEA9j0qJZD7mVpfDjJXB/sBf087w+I
9Ruh65sOLHCXlRswpj1PVgLsXTr51YEz0p3vuhzFhs4U1OhqPz+v91igJrvE8OJ61O1RfIOaGd4H
HzRC2rf5siJCknSs6hHOSg3P2u6wpSjfAQsSBqYX9Fm1dFrxB/9GH61K+ESpk6G3WcAIPN75ngXv
K2ddOFjOHBuPusF/O57Egdxvb3JkhtRmeXLmIwBRTjnqUZXRPv5kArwmfe7CyOTmxRN0lFlUBNw8
DN8qwkB6vjvOfwq3fNzeCN1VZFL8UqtQiVyQXbLl/8GzVL66xIG/ip96Gov1xnNj2OUFRpJIlfpv
+vVkWEnyFVS9Yew3D0W8aK00GKu3iTHyEJrrlSxjyJXMCqXnlCf0KfzsX4kW9nvnjRTHJ3uxu5JT
HXl3JsCD/pl/EZc6jj0ze7vfDh73lH/WrNcZYdn2pHPNlviwG+bHqlTJ5m/1OaR5Bzf0yjJFRPAb
QVvlo2rF6G5N7oCwz5hdQEmSvz7GBgjWy6y9NB+Qyn2BibpnvdvE6KcSah5JovtKZneKbdD91yAZ
mQRkya5yh85r/LPDHZPqYv8VDMcTMsTy3DyKBmI1qpJ0faS13s3cww6R35uB1c4gGvWuvEVbiv5d
/uOvPhOuQNp0yrZSifKX46QuXNnxr3UT99l0cPpeG6WrFHmQ3WvSpEAC0bvY+VD+d2y0u/zBhFc4
vfjaoROCISfGexjYOGG0PdO/c2sAHMEv2XBhZpiBND7/hvJ4n9bFBxqfXSbGnkWEUklDGZPaH420
8J25cmzeYB3oTw1J+eAYmGidEcRWwLltuA0PyaTmg+oCO0mVZPT6cUinMzzCGIyXq2K5G80UNJkt
ySjCZ/7vw47ODd4bCdiPaeAdJr/CNKzDwAxLqDi/cmP0KHE9bcfkmiaLH8OLGMeyQ2/iwmnZSRGL
Xv6Uw8LlXAZSudRPU7gBrjUvLbVQETYBa9HFHxxekdCKsd/SeJ++Z6wYYv7I7Xbk88rJYJ3olfOL
pT6BqwVqGdML4ZQy2h6+UUlIOl0UtOHI/ZzY4fABpg/WPFFQ039v7cxv5JodL8e0WS8swxke4+nX
VaF+whUY7JWfqHfDD3sdTTciQT4B2bLWaOyhrvtOiYa9G/0/60i5qMfiFK16r02dA/sCGfytvRkD
8cFjQENOnZusacVDNFygDpV7MMOzFLLsGZvbva1N0b+RxLml8HgauaoyKs8/GsdloB+ydkqpSRl+
jDgDgE1QYLhpeATIZ018Bc03aJ91vMz7z7ITy+4T1lHj3YK+3eKmtHKNjvJQaMcBIFBasJCsntRb
iMcpOSsydb/b2w4nQQctj2BcabD+kJNGRqt8eR/BU3Z3zFTJq24uZ22qGVDFORFFG6TWesPYlS9U
I7/5qlbNqyyfwkt0hWqTufMHM8S77RxMyekYEM/rPsitLEzps/WPlYSpuNa+oJHqTPR7lqgcBzJs
K/PIcks7OEHrD9aztL4x8QH5JkKhhuPzZiGdbT3czBgcJ7u+CXlWoQrqdnclgIqjqBsRHBgvy0Zy
CBOwW31XnH59oI1FYGi741E9NmCWD6oqc1kT6tXu+zQY2H91gXlLUKXd0Yds4w9g/LggCQJqM0hy
9tV+qTi9c3zCcBKCw+pHp5CqpvmCkErYig4iwI7fWPaqpWEVmJEmHna4MdL+uhJyw2IdYAFx16dp
haT9/PwgOiv8t9SqPTQrxG2SUeE5s7BLjd8yuFmJ7RNyWRFz808pl5e07QSSzM3ORj71juCfxAN7
xA84T0JwBj/+XcRDewgpPnF8ProePpg3hpD0FVzArbsu2A9SRGB0Q/0wkglAlgzql3JPycHzFRBk
O0C9RiRTbtWNtCSh84VjY/x5wXbv47dAr63vvadci3rb8tSRneIUPvjjQmEvuVzHIQE2J4nGpavV
LLbqi1mQzHSlnMwKz9KlkbPDSOhYBW/qyO7+eO6Ii4jhK2bc3+FA2d9Bngjv9dcIhKQmO9QklyGa
QhfoIzGQ8AoQQdsqcDGkdjRRIucSBYkTusbEgqnGQx9S0YhxbMRG7QLM1acJCi1/hVUiLYL4g8/P
zuuQr8mcvAo9AbA61uDQY7Le5WYdsZKu6cQ5QOtgL5OuXH/wnKvpdBwQTldZI4KSAUm8PfipB5yP
ZKXZs1MeC6LTWE5JCDLekhUXeDyhXt9HKwQMPxKVAnaKlC/JJrdMJ1wHiTx/jIm7Hfw5/dB/8dSW
FIbl6k4GnyGXOHF2qGAuVWL82i292eIx80zW0WDq8ZQNOMZh2gWpZqONPkdIguzNwjG/KwjUUJ6w
UYy/k0KVTWQg1JmR3hqVtFQdy1SO2UcC3TjYhwndVVnRr/VmRGDx1taNRbt7dAQLAY2queuCTbzz
rQBE7f/9UUiFXhc0V/+BAS8axXqQrAcbgeU3HyOE7hPsm6aZsaoptz/conLuW6ANkuP1hCQEIyV3
+DK4HylfKIZPYLDCbmTWDVJ0MrRoyMHUn3fuq0MBXkkelWDjvmX1xNBAox3sgOkg27px57x2Fdnw
ojfHdXnehvARYI+sCvmEpGY9d37RQPBWB6ZBme1V2b9jw4d/6ACipK4Vmky8+D7O8iM4Szfk4OiX
4ITlHLBUt7sDXvikVjhOXY+IbVyBWQBwWkavpaT6tvL//eeNvf9SF9UxxqISQ6q5jSFKNJOkNwGR
Wed6+wtS1R+tYO5ybSuz3gef7PnEMWzx30F3O9RXsn/y181vgmXGxKhoUY2zp47O0aUPLJF9+MhK
NprP2ffXPXuBPwHpIhLYFhAHT2h0WdMB60wrjMuZ6QiwCQwmvNHhDfISW3pGva3NWVHd9BAQgBSb
NrRjUnUwUH7hBjkoCjihIn+HDzGtqJ5geuQZMjJkn52skZWaF2RB4Key/tvhedixioZTof1mOGbA
/bpB6QobSpjPc8q/pv+0yB0eJ/oC7Z+u2pB3J9134r/4JrQ+rvh1vaQeQFrQP6JsZngfMQtNCoie
k8iqihibxfkDvWtrjFkTOmPUJ5jTKEk1gVyAD/A64qwFSOfWcA4STmF89sMYc+PjIzlBWR2VG16M
9xC/l8RZlrDCqmhaIpXGhxjlmwftIjtHpUER5VPhohCPmx8F/FCyM4d2YSyZKUDYjeFn11sST2ky
O3xagPaFYvmyNrKHSXaP4+YJ633L4IDvXgsVWwOA0pjTbpX0NhLEBncfBm5GF87ZoB7liSzNHb90
Mg/MAfGKC1q353q0MrSy5L4NY8OoDdakiCHbyJjnL9pLDgvAkNfuvI2UfG9GkUXK+pGozIaKjIrg
pxtN1ythvRggtApwc18Wb83ZIR1OhP+6RyvtdS83PTk51BQws0zOMHlSMRbPlMhOCEQSWd5qQfLk
6WR8cuRHhsr1p2lI3Mnkb7xiICLZ/T8xKgN0/NPbpy19DApSacB7O2pcb0bVYx8GTn3ldG47bnbJ
P66TcL3oaygwT5FeJeD0t89dV1oClb1zw/xp2eORTNyi3jyISc/tUK+sSXmYb7lSfvrjZOpx27VN
pacC4riQ1zgIV4es65brNUqJfyKAVgP3f1S7gJkOAk1oOCu9Qu2bnICmANtIUrJ3/XurfKCYYaps
uswB5+fI+kwmbFpSjY2sKQ6UmFSWUYwasR0YCspL63sov/K/KRslPyVEltX+tfTNpmfes6LTgLOl
Trn48F9+sTUD4+cWlLaxMQGZ+F9RL5UFjm/OaX8Xm3fUfnqdqtYSiUqWIAF1Ue111Maui2H4sxp1
rzN75/GVSzoZZ8DtIB/fDFTu/ZNGQWCO6XPffkDGJIrZLImwa2WKAgTeZvwoDAgsUViNt6bYQmIu
L9QhFXxegCNwPLGhEWsFk0f4GEEi69D4hVWUox3HAHhRBCuz3wUQ1aiQKhvp48Qqi4CPxfE1VBSo
pTgoTeDdSilDpBOD6+VFpYkad61c+GvEGtjOh5c3QIME8aiZObJddII482y1nzbfgJO/UBlbcyrz
8rp9jQCA7dHqGKk6+TRKM0DMiJsa7WwouvaHr+/1X8tPE5bjNSrlQYlNL70yrtkPwFxuhiU98ewi
pxcwVQmcjKF6hdrProudMTiYn0Jx8LJqEQbPlhtWIdWj04DFdOSmm4fRCRjUiOWv93w+ajX/W3mj
3CCiBnecuYhOp4vT22xvc8FTVnDXhiVzCVkq3LkyVxNSlTtsLr9jEforE32gLTTMhGyyPYqOMc2H
wwVx972ZkiMWXX6sJqq8yvefBgnGHplSBxQMcA/6lCGkTDdMptS01Pjg/PlQwcaf2751mqHL8sT0
RYcioZW0qWko82M0ZTnqy2uFu7fWzVC4JcKch6WbiwQMNZdMLBFbhmqVcN4MEVuJ1b56Swn0CHhe
StHzi+15AXKAegDP4U5/7bPs9BHTSRe+EgGgI3gKmEFCLUsNwRUK/Sjk4bdSRNhUob3Z9S8y/BRH
GuNCAqGcYmBCj/HVkgw3Smh4GjclP4ENsAMrVHnd71ft9mSumay0D9hTFoBmsgIEuAmkVt3BxuMv
5IlZiul2m34Key+M5RPVVDzOa9NUnZI/642mQGhLbAU0d74cwMVAy1C2qlcyn1pbKsds4ufWVpMh
jyE+vy12t+1wwg13UmDo7W/GhHvLrmAx5lCgBSZ6+LhJFF81MCYthYSYy4wsv2aQ3XUoTIErzUzt
wBeMLm4MATBM5A02UqWBAVoTnP+BVWKaOdgEJvIqRp0VVILfKXWQOv/WVaZ8uuK+yK8vTwn2RP+M
eJi4w3B3IKtptvX1ilJOQgdSb60Ok3qxfeEjHB1noQzYB7t+MvESqGmzXwOCPMnH6Ik1tH7wDgnf
aB+1jP/HSY2Lv1pRbCZNc6zHl/QV69cIjvumsxRHH3uHsxbPsRvc8RMH1pE25rjYAjvljTWJhPv4
yYd0AlBESvuasuD1D+ilZiTGvoho65vneJ84TWD28qFYd5vXuT14SD8xcxCJ4JpOz+Vb7HWdYHCn
T7syx1B6hzN1sj3Z6kdjt/Yv5wT+yoUC8BDcw+Nut/PWgcWuJ4mooUDaT0oM1Xw+v7Uo67A0bAoy
Y9sWvQbMNaFCb8j4zN9Zg0QMCOPMbhV4gzj/DK4WpH8sv9zoVwRhsX2M51UlCHMAg5sCAXw0bMiT
r1b21Fr/Rc0G1OvolBtx3B8IfpwWvOjzLSrRS+7tDxxBlc/TDayWluD72v0I3GTrrNC0N6tL5Vg0
z1XE0Pa7TDJjZlkIUe0W1U//MnCs4nG4uGoV3fJXTO9VEfeSyKkCOFYdFkrVol4VK5F5Rmunf4n+
LVzrmlykziaGSRgpHil4/8ugK22gP0o01pW4OlzRa6v4zHrvc3tn+afRsDdsIGlKaR+rThbGMBvG
57KBFGjl4Sw0FwXAH3XyYrACiAYd3W/ScjUbSf69wjJ39BBYUimsBYUxwOAxcBelmBs4iAgK1PlK
RrzcezF8zx8je8LGiBlDk4ZNjsDkpBK0nIwt0mFTQIjfT9r7S3f9iZqrnSxAD1Vvb4SXreHX3SLs
qPRMaGBGSE6ztCZy8B/DjX84cghHkAnk84MuVfVPhAHKRY5Mszu/cXdSKc2b/JF/ZaS+IL67M1mj
jcc3WoAEpanaa/v96qn/OU838t9Igxa1Xj7fBOaphz+0mV/G+Sk9IINxja8oDKcb1CcBIRSlEdVH
3COrn7Ejoa3D5W3UzqYsp8gumL7YL3GwJhmo21pMSEldAQdz7KgXLIb0/wL9dpcfpK1znPXzpRL9
nrCjWdQDUZ9B5B0ZqJTGEMmCzF6MexRoLtSIu2wqWOZXd1f7S9eW8hV7AXJHsxT+Z+FIFCS00IUi
pd0ZUzFGX2x+2Gm7OVQIbJQu0Nh07tYRvusqS/iARPmhMBUER2vbU2wYblEeNrpGSx2DJbs8IZh/
GkzcUzSAcdKnSX13yJKMvaKDT5XOQcN6Sld4s+ihK1hvtskMQMmDImoc2iZZfAJ+me/SZtNZW4a3
8mbJ7UIDd78ZCmLc94a9uiy8TJBwm8j72b1UCAvT9bz81BmizNkN8el2bz6TT3zziq5LxhR9xTcW
zT1eQoiIni4NTP4uMihPn4NM1V0BYkDJJHwjGIDo1a6JdSs5K82jMMm9S/vAJX7wkZmDha4zzX3g
flyoLn7GX5u1aJxiXslsK893/zkhvMUatvcFMc9g96QmaJl8TINYJhfqGLjLKufEN61kE72WK76G
1mqJnu2W7XIgQ2P4Kk38bxy3Lhslj7/mJt1ABIfZqmBRxRp6FJdDMDkExAfv4UqywJ2TXia4kpog
FZhouVMYS7uzjUzmrAoUW3FAXy7BhZNyQTibxdqL0mdAtIgWvKcVt0LwWrH4tB4GDiI82mQZcimF
7IDKmuu3iYx2EevIqy4J8WviPcaJaMzWUvs+cZdmUuGHNTfbGZR5jxndWdxOfGrp0EYGPaKuUH8V
mJiQ803CbOzdI3/FeC3bW/CDh7sck/3Lr6uWq66asTxqzZFZvpw9PtWSbvmSAWj/L0EMFH3zUIh0
Y/OXcqBphrCBY192oqoEtNJk4c8jGo5XY5Hqb6xSrY7jpGi9R4kNyQjQWuQ/QTkwMseTaxKRdNY6
kDJHdoDYr7xQLlnkdZCJhIewv+9/2JMPLK0E1YKJa5MsR4uP6Uh+oT8cV6ArJJooILM0uyHIsQS0
/XFitzin7Bu+JE08Fann4gxeTQ3dkeJJveNTySDjbjXs0Y67ulYRKQncrEUYR+ZU9lwAaiB56Ljd
+qUajkgh9TssaJptCABUDwhUqKCPZcK8X6R/v8uN9cr/RZLcQr4ty7yz5lJUJACWXXext4KiYZ90
lExMGyQYVfsSACveYPtu1qYVpGge57nbZVBbzSeY9oT3hkRbfWCis/XVmd7xVbTUW9yUXSAu+hG2
jWPB6F1lp1OHtVn6JecipEenm6hB0IkCbMQ2Tpxt6dymHcEwF3XVymGL7+hEj+YkhmGzMcyqexFm
tT2ShTElRX5biFi69WlJObih8w8l25JUdgXNo0Kos9r09LrHIhFnqLhF6UvJTEiE6jJ/vJI0T4k6
vi2cIT8vu2yACUbOtb0JLOM7UBLBnW6NZw1HNAAx0zsVgCI9du3aAKde449nPlbUu3eR2tA4fkQh
FnIduZKL6e3Nz406lYb6f8O8VHljSsMCQhlKItz59pWe0iyhWRAvHmctvOVunHZav6+3Ex0E/MC6
mKLfEebS3maMFFfOjyUGsRLMeTdv6YjXM/RjBL1Ud9wa9xNx/kEJIv/9px9YNz/OpzYcJKm+W9dj
qbeBNo6IAnIftRcD5wcuddHAgRuM0uwd0KSd+6SUtJ0pTvObl6/xTkkAYQv0S9Yikb0xzEAKMl7d
DigDVMEqs0iIWvjqkpQyKg2/hUr2bzTvYFbv0ypUq8c7DEkj4Sl+5DgMvnwKwGHOFoEo72mLpyhc
eTWHTtaASbUBWnczA89btE4cldodWkx/aU7FsTHmXnTUJbShGVQMYqJAtWJnUCVyIw38M4Wt7mMV
RNklRNBPhORWdNjU6zNBCOaMKy00RRmmJ3T0rjxaux8WepIwqdt7a0vX6AgN4F3NbENRZK+fjcl6
2j4e0Aml3FUr9mpcPxXF/ku+U7v6ZpBs3E+H+omvoMqd898rYqsymJnYYTLerbqMpIyFBjBzgwq6
c2Dr2OUchefyrnc878R32Hnkq6cQpDtcAUUrn6720u704EFAYkNPdq1Ou4PJR7FdakPZ2VrIDnFh
9/blvXhfZhCYrXf3E83WGoV8BT+mmnqkH3Se7zKOT8wgZnYVdyWaxyVHL3e+oLVE/BuTltLy/Tz5
2qWLaqyVkYXAjSYbG5qlbE3ecNlPnMe8GrrsFP3ya1D9cTkcGj+NXr+gD88PcBXrFMmJY9rfDdCO
NvSTUPiBgip/vnpUdlA/7+DfuNlGUyGrDtN08H4Es/JLQ92rYyqdXYNr6vGvDv4maKkJBzaWCilr
ABUQ2LIkoYcLkO9D7JMpQsOcKmae1XeP0krkLR/8A7Xjv+V8+ttR6zrqvsshSQjOnHWezI6VEver
18log/QdNyWYORLo2NMW3wU+CgeOeCtB2IpOPodhmMONsH3wXQF3yhoCLZ4yUf6b0agB+lmOIlNn
spfmw8x6I2WnbRlfZRJrChTyPvGqs+xz+b9D1FN/pe0crAb9Eyb1nNtjmDQrHsRpbijo8i28PrbO
51W9Z0mDJnFBSvZwidY5Dccc3ZdnrVWCOgZ/vsqB1VwD8TYkCi83w+titIE0Sq/YwXCoikdYEZij
CI92tC4mg4iGuTw/PkKYToMoYLFTXQovdjZthNl0lt1yrAmR1Hpdo5IrLurKeTBDstJOWMjTIIjB
bMxl0gRWiSzocIxWq4gZmBOh03JWxFAN+YsrfvY0aWkh0/9Vhugl4bxQmeRwofegvluLvSKDlZUx
mNHyak55Fy9c5CzRXfDcTj9tBzskc+OVH0cdRfVXPSH5lhThl7s6wHJ7CqGJiRnvORLp23eU84IO
cG9uI2FXZ8OTpb1TTCBJmCBGECg2+HHtdwUjddXXr4HU4nINgs1w6nU5wXVLQGj8yo1mNTFMdgGn
oDnkmzTSav5xCCrVuC8ovQpk72HbNdQoGlvMOHuL0EIcpsJlzoIoU+MRs+dgOrspTpV7TgILmwom
Z6ukVr4KRNg4thSYCeGXgqwv4FPgE5H9OkIScspoCbo8Tn947prDCJs0agJfN7/50AJbQkq6qOgU
57ADRKbuhyLNbKQGP9xRh9C7IXrD5LZxnFZwTxBbymmpgcfHNWIv4NNcRkvGwslAnG3kbJjHdnQI
gGf6OOTAAHKNvnksv/vygJKL50ZLQoaA5/U6Fx3rdl96mVN4fKQa+IzpKbUDNBcOZ6f44wQ4SqGE
ytnerBBwSfK/OtBd6j7tzo3znTYuclqHB5HS2wgXmG2y7SUBp6Q79uLfKlZV9ubYurRYeUbPhBkD
/y1lnroXIZAN7AqFqvYuKYDCO3wZi7Rhto+rSQ9pAN4Vb+DjKPz6T8qpjWuaB87Hdgm75fDxibEA
sTMj5gMOtrbLRjtyWtqYGIghyjh2N4gHWMficUhE54vE7MeYCoryGGRHNtCMjOQ5/C1PT4B1YRXw
qLbno1zUuPJhdniGbBXGs5nfS91N3EknqzLmWURH4T42Vb7tcI1ZcKFRI/wfDMFQJWdC8cOIapK5
l+el6UXMdyCA5PcKgVHRUljXuJDgfb7sPw5Wyfi7uJzc2+XrGyxj8Sw4lI0ZgB3jF7z6U7NEUuOi
SECyh+Fc2lbFy+AlDC3Ojc7ZuhyplzCgljV20D5Ns5t3xJ0k9QENVCOW7Yz0pV38EJ9xLwt88u6b
YPujQynp7MvqP6K1juZqIZ0Y/dhHQQEktyYjTGLHULfvFbk2s6Cwlp6l0l/VpDWFfhIXsLoNprmU
F1v3A5WaltmCEwvAHpDIYANLPXLL7ZoDkD9IWLveA4IUi14s+Akyr0o+ovOH0NArg7VXuVErFa+1
f1K+T1O28/ssA5/XdFcEFpnRJAtibbhzaES5f3M/OQNaK6b/mQtunwHYY04qFDMn1oRgQ6ThUx9F
ehdnVCZiRPAssd2rPNlhNiPM+vjAgav5lWnqyIyhUlIHslf1RVIl/U5TBZiIRa0o294N8Vo9FaXQ
kle25SADWloDPfNMi6vPcOIvo6H6vK98sq4FRXzxVzlJWl+lj8h1jVJlO722qkLParJOV+uSSp3X
cvpTBvfZ0ktur9RtsV4msk74y8l1F5rUmdUFxKSmpmNwGwcCAkREVJefzHjyd6ZNsA9cFLsipuBR
Fc804va05JbLjXQVBcipIrBoGuyjPL6ce5yHA3Q89YHlmXw1a+3GWOMeaSCK6ngu0N/PmiU97TX/
EZDQ5lC+5iBf/iJ2pQgGF9easruC3rTWrKH0aHK7lzZVhwSF2+KxxgSiDta8P+appM8b4kmttAaX
47hA/TMi+S0LhNUollEd+m5R9sPJQ4s9fo/mHN6NGUjtabM1Vx6QbJVetPfP5BJdefVc9VwjKGL6
0X8hBmQS3EtYOXCBLisrLlSB7ICFzLGcORhkD/vjka9GnQSz0hsP3hdq89cScpn8LclxtlHlovM2
W/ft6crrernuzTP55Uc6vd6rjaC64z3WThsXERq2Xk1NUse2jfgil3SxuJGUdoxOTuJ+fOxUSTod
K3ImDxv7XMLTnseHcHJeIz6I87aqvshbWug9fj7ppikWfb0MNvS+ksUuSD5gInJvGaXml4BQHrID
EXZ1kdP7Dz9qiFoph/IktH3gtUIyKaEwwASQUP3JfYCOQQlLrWJ0GwGI5gm6hCSAH6gwuJQS/+CL
4u0RE/oddOJ/uyJSIwVgAw0tQmVNENXgQyJj+XFFDH/iYL33fP9L3T15JyHS0827w6Ut5TGdJ2o4
6G3X91nMi4+34m3f91n11Wjs1sKw/UJCjwu/chNZB5iAxyj0sfF7NCJW3/gkJKH7kxqKF5cyy1xG
WdTgmxJbfz/35//OMjIDanmu/wF1ZHPDvV0KLjuU9ObNA43y0Vnq/7biqA8JbJh/4DoiH8RBmlCN
jEimVBeWvyKl52JgH0Z8yO10mxNSx7IatdWoPP31Vj2UHhOm8ITiRToZeQAvrpCqLPXO2H8yDMnt
Atuur9N0VbOP1Fwfgfrna6NfUmG0yqfitQrH3S+2Ipc1/MbVj6BNzBumgERZmNX2L7Fj7Xqhg85P
yJeu5GM2pKh6/32R3YDKStP7+mFgHWJL4axJg5S3eBj/vnwgyVJv97PMUlcIRjgVO8qc+fITUUrm
/kJqiryBbP7pY4ENenLC1CxBmcW3VRKaQ7Sb5j/CmuiMLJkBb/Vrln6CYPinyZxJZOwangguCAQo
8zDpubQV2bvo7LQth9SOq1pWPmH8sH1NhZXj8U/CQWpppY4trYZx/nVFbtljETact0U3wK9MldPP
KI/0pH/lUxTYmkhJCe2ShOSZw5qi1EGVBOf8PN2Naicu8rFqVmA9G+5aTSm0nQbJTBPJ2qOLS34H
aIZs6SmrbcTC72eKt6mJDjVWrqROJyX9FI3aweSUjWbRvB4Yt7T1716lQVVp2aPB6tlkLvS6NljJ
wxKwsGMlkdJ3yklpeYSakNBXW7NhAnLH22+yWdemekJzaSQbxMriZEeFTd+i7nMLydn+mEs0bCQ6
rxA24L1R7AYzhSyDiSMkDUEZQXD9cB5W9dQwOUwnxWUoF38Svk0Png/5QikGPOfOXUN3C91HNb1W
kBH122ccudOdK4cMOsGXBjti5zvgX7uHWzwVo28IgpsN7VfXaO398p4l4RjOCf8g90/1PW8aLIba
TKDTxPy0OUPgmg3M+mvQwnx7T5D+7exwqKpewhfFvPlkWU+WsiftoECWZ0UtKZPsddzvRbzI/3h7
poHCN7Qg+b1P01ssAS4zCygQAlCiQfTWNqsUeWvvb6wVHlF+BD5TL7POhail7dG4DJu0JQj47mM/
i2TuxMf0OzYPbqmWxvUoWz7Yl93U9K8gkVp068LvN9KNCmZbXimRp+14A5kcmX4CCTYnVaaiauPq
FXBI8gMOFs08vLDv4wtVcduTEYvEDkb6b20wfp+H+8V6+7F6pJnsbviTXCnB9VeSGO+5DEhSLnVa
mnmcwCSGYZfXYWSD/uGgkN0yInUmmOrx3kH2cnkGCcfqUyNpgsNKzb8YOUr1OvnUCD28WYY/zbj+
NsCmnmRfY4CBRPO8P/nJ4v67pAJLRuqk9r3TjypRABnBhFkPuFrKNF/6pCSDd/466+JaNP7gHNB0
3ApSWiMr7ii8qnDLRgAfE9arV+XnJk6PO6SPHJB0kGmwafLb+znQqc0qJmgADGKufsyNWPkpwXkS
ATTbxdtwa15wXfUOBxXm/CFRJnF6Rly7FWWPSmTwnd7C8gIfjSnNNi34lYL5F5ouLPJ+IZoHAWMk
aS2HCp7ulInwelYOgyhbfdjsSZBRyRY4rIMKJOeEsRzYRln95jADj0I2y1aVGCylPjHx5ZsxI1Ej
E30LbB9hWrkT99mAmkdlSN4ZS2NJe/yvzR/1fojKHuTU7jhPpECZgv8VgkQwyjXEa00W3Gyu2nM9
bGDCKMGocToVkj/azWVJ2r2aGzpZa2gnD4tWTXtRc6QKqzEYnoFSTrLMf426pMHU1fppFSqoitme
olYUdeRH544fqP7oV5DRhmoCHg0UIXXqhcvpWEMNJ1V/11m0+fDrNs1E+LW/AlGl3l4+UQnX/n0O
VVO82q2QIPDiKSceAiOwDxI7BWgRACELSqrbf+CGeyPT9awOn61b5W1G3TaFtU9W2xxXPRNOBY3R
WrzRJ6MhHJtjSTOPNBmcHiSVcmM0SB4VYGiBOIIGhN5Rbp9Fxlj6FnMtkL6gnocq9Uke+YOwrdxz
SwFxl9UMXqC1uvnv+gRRZQB7OVCkSTcZFY7xVzqBXAeA3+OXX+KcvpU5l9MuulS23w8CYdj92VI6
w44p/yKXCfit5bca5JiOkEaSaWqNSOt889eMY6id/Snh824Ig0LFDjeirMEFTcaw1an+U+U1D2ah
fjwga4jcwi9Vk0LyboUuxRD+VwjSEqlDOYdWQVns/XCbe66SpSNecl9QI4jL+/bRSNG8T61i76UF
pPulGuqnhVJBflBvg5+/YVy60Tqvn4UFK1Qj9jdfJh/XZUhQi3SmfTyk5AChYKyQ8dlEl+TYSO8g
RpfoHUQYHmH0hHnWcqSAUhLsoxWZ5sVt9nZdMh2h+sGqgVv/qyA1CMyYnaXuFcb1YDQM595D8qHd
IybbHyO4Adwo2Le1aYUUUoil9vk8KCikEMTPjAWgaIOaAlkRMBKx8Y9JXcu1TUJA1SoP31vlPj85
QYYSwXS0P2sPXTCXoDiiyCErnBhT7QF3MG7ipIj/h7m48QAa5JdKjISaa8RB7rEO3smz2seIVvwI
KN0DqXX9JWQuRcre7xBRX2coyFeYaa2ZXWrGh/6b0SBGsjHGGitFLZAas8qhRDkt0QOyfdZxs6b1
DIiyup96zki/HLVgTZdvFQkxhGHnX/wvx0o4ACbYIE597EyeHuizNyyrk5MJVWPMa3S/mI2qOlGo
XROpI3fg2SIzg8pxaRJ0IDzxC0FJMqoGS4wsA45NaYPwVrSzOErj9NFGaSjUmSsuF5m7SyRIsNZr
zr7Hd7nHsr7kG3VKWy+SjVIZwZt9IPJjiLIcv4qW5suo2/oTpDbQdfduFP0/hC96gJLgpqGZ5MFN
cbeW9su+OEhTsMqobj18O4WfRe5S+9JW9t3esNlRKoFrxwQjngcLccFRY4QNvfhj3gRU3sJatAsZ
ZhlOaXL8D/ki8oCnnycWnmsgXOlcDrO2BIWVrwsilmqxPk8hdbMzIJUwxy8SR44PuKDPuZs/jhmx
QJnDY7gT/zyCv0s/EKic1lwRt445BYCtN2Wlyp8yS8uNkmGVKzhT2/8LNNKeDZhs1WrpI/qX6kht
PgddqfpomZerKWzOukrqeMScfYtFEMeWRCjI4Wmx8ws4AXp/IPLFNF9KmFYZeQiMqaKL4uuDusLw
BU22IknyxehMomD80pVXEtUGZV18zyykfSCGCTXGK/gqgIZ7mnitsHiVp14xXC2aHxAhNYGFyAzJ
hOtWRl/POq759Sx1fds5TcGhtJMs31oQa/CwcuY+n1NSlwXkHVjWW0f6cPuEI4nScVfOzWPws8qd
ed39mc0EMJablpGz/EqvHhbh8juRH5u2QMa3WmjPueT4zdNT7c1xo4d0z73s4QJrpzmOrSs34wpr
ZlcV+RhkHHZeHe6FWy39ckrQgSwWt87ykAEY9MQWm1Yq4lWexzesN0tn9Onsn528YEmE7AhqUF9g
4SkQ00tRRQF/kbIZihxcbJpS+35VUUX5qCNnSkvGgL7G3zSW+zeK12A2Pstcyxs1mSfB4/bpJp52
x8oof8PD3fTLLyLVSqyhEn6MQABvsvevKqYnAd7QrRuqCicAS5tx/hpWHVa2vskiFADQ0YAGLysD
yiOwFftuiC3A1rs9wgPNixs4WqPbIjq10b/o4pwJjRGdI6ELOi49CY3Srve67uTp0juDZ3Ovp3g/
yoyzU+fUZnV6+0XM3iQwyGeeuTvOWeIA0/fs0KPMk2fCHBtpH1AfjrdrmCmp9yQ0vWn9FhCuZ8W/
JSJcmWmGCanqrLVUYSOETHwmovinipZNI5HtIKjW+orNHCLIQH3d9BuM3CP03+V5ExDPZ39KZgie
hwF9rnqzHzWw5ik99U27KQTVaLMDc3cmYHOJsDkmapgs9m2LshH+2foxidL1kPxky4QCv1Lc57ne
Pri/SVi2JaUyohaucMnERsXi7AktYHMX1bn+WglEaHEYYfw+9/HqcuwReNEvjrE0/m5fVAmK1VGa
BEbyZl8wrDcANydqNHSBB8orCPt3mJaMJ7cS77sRUf0elfmJQyJbcydGeyyOFiDCoOC9VQGiRe35
wCk4K7s7UePJdx4ul4e8Vpv1l5/11jet28cJeq4VoGwp+LN4yZQQN8GV/R79zjM+iK+16WM9ThVG
UikZamGaKhP88MI2+eKSFOkcf37o6HIOe/5LzHruzKMaR5yWbY0CcOCKaW2QMK8XCy3wwM9F2NbY
AMopYN4nAlH/eeSwdfIc2j/cZMpxbAC/MWP9llGjGZCi8CdEepj9xOuu2lXSCzbuMFc/AjEAyoyO
oizyclsy7F1PoBNtrd/u5b0Hkrya0XOWGfKtxx3bcU2FIo/dfZpliyn165fpe1FgMmyAExjL2Hi2
HFuoT34x3jm9CTBnKGub42whw8zkmIYfLWMRnAO4Z2hO7124EtwY9LQNFTTobyLz5OsZHx4ccSq6
5B9oR0x9+YXoVa2qFlUVDALuqIPTgoLOaYrIyclTH8ZP6qK3Zez1k/vqtYZP5vSf6TgThoEKggOz
Ag7dqd+4OqUnQ1zdyuK0llgVX7voZWELA85pfD9KIC6Bp3R/I41jZruqrZFP99o5T4fztjH1jR/6
pFp+/fe4AeqACCdyZ1ctV6YX/g4a0S0BxyE93RQX1MUWRAFHkr2erndOQGWy4SQ1Kbepu6QDP8pm
MxIl0AAyxZ4kkalHdc2ZNLffJHurg+xUpFD4gm1AfY4RtqUzIrWpf8u7jeQEVsMe/t7z+yAS6Huf
H1MlPt6FkAiKkvqzBNzn5DpxYpZO+0sqJlcDGi7rKkSo0apS4secvCXjNzCoocErUT3ioq03fh27
fQn/gRlA+hzH77+goq8WENGPdMCn3SKHJl3tfu5Izf8ZSuhWCYXv237Cv/7BRpBM9ld/L33SfiGX
clc9OlqR2xPu+Kpu5YvC1pTSUVD0cDla+z6NGiCuuQnchsCJaY2WpfjKXCPReoWzehsiyZN4K8qZ
t/Y9F4aN9DBDoqetLTxaVaHO5+VT0LPi52xBkcDORv7TB7eYT9G2pXL3EC7qW9tLTCD+sOi+yp9P
nuLzb6Z5s+UD/oGOkGg/Kkkg99ThhYeV/iiU7CHwNx8tb1b6kZoTJtNtcLb5nP+yBvNtWi8Zdi6q
vg41W2NHNOlEwIII0TEZyLf0u6fciBUgFOxyAN55uim4i2Jy2fBIj4ZdjIVLOdzwv0Pvsu4CYR76
adFnbiHEqQ4r9OQxWPgjO3V/6zalkAzgr6N39r3A3L0GCWk51y61UMBN0PDLY6p4CCbWHzw8/RVl
U3G7QPYWdGbBydOPO1PglPBYPRGAnYBt1/3xetD2GvIzdBrqgtDaF4B65cnQTOeOhX+Vo8b4cgrM
miUPHIkSjutdySkUxB2ZjgC3/bOMSoJyMpRXchXberdH1EjYYvULuvObqUiyxiu6AHj/cPCH4ay7
ux7atQHig1Kk2te97Ck57VIjHqVlg+K130jKB0TsUD0u+HpPu3q6EAYHYgsELYg0tTRMHThEYeo2
iCPrKEdPEbuZK/CzZ3fIHPjVhvrRPG4k8dysCNd3YldpGKyCxWlFxmx8zydg/kd9mNnPhsAlFf0p
ZdtESTAxlMAELBcuKDCNpuNccZc4BbipBFUNtS8nb2TQg1Dqj+ymLNeogFNEVSY9/OvPPZc7SAC6
1Un6aUBmSyQY+YapdBPqElY2buehY/KlwnR3galPKAjUuHsVTl3CGJgBxkfF9O8TkydE03y3bTWg
ZVuaw2nNjQgRcqmVJrODdtmA7yFK0rLz2+laIXmnB7Pzr62lQH0FxWh1GC6jbL1pPmRDqmzoFUtx
1c12tFXWIpIL5irEr1Lt43tRWLCC9xkEBVj5eRU23Ua8BY1hbighnBLBauQgpTMSAM5MP4E0eg/P
Hkq80UoPRZ/ZOuEv8EJRO592OSa8PpZUB6cNeYJze8QhJrFZUVVJcN+0+q4N35UcIrUbGIhzJl/r
dOvuis66YEV+70vxoEGN0rbRsmBK5948XIcmdMzXL/LKX1Yfc1GbFKktVFc5mW4icCKqzHzfn7Ww
MbPcj5lQQIDpMd4SDwsy6z6+KGlSwTse7m2QHisK0uItI6Fb2tyfCKv5KrLa1ojE8u40K6yfJWWS
SgQmtFcaKY9mGHZh+UHogrDAVEip0OAYAdRNp0p5LUar2Q+gNLZmfAM/2LLyvMvosue9H6mWdULJ
RoWTil+51FGnj+1h3gQYu3spNDVoNtsmxDb72IKta5heRK27b4PWOftnRf1dCdHtnjudOT7/iFuM
nKQ4SX4/ekAOzTR/OZdVGbTspoi6+vOoA2uMY+YJJ8KWDIamvXGPA37xDAyyYtBCd9hRHTrXrVFO
upIeIQ6GhrBSvFj2TBiHgvDsr/IyFtOEpJZA8eXZrinrKcLWtqTdP2DECOB5rIoa5Eyv4/DSkdW2
anRERxTGb3tH7Es4BhHXN1QKOYnjxAvEgr5rkJNWQfEEz5+e5LHZpxC0lV/oH3e90ymlDPJK7VmS
nec/OzoLEP62i7Q7VPKln9KGkohAwStS9jlBG1Dgs2ePUjlM1VkLsjhvb51HTKJnezNV8eQII63x
KJ+10RAJDxiDHYdUgxxOnPLxPzUXPuT0MyUSbA1ZfrnKDAvGbtZfb16nGcOhElXQfd7ExI2350ta
lhAw568plKFmWRkkKvB+3izZ2XZOIU/LZrJmhc+jx32MRIINVPo9kpzJMIjMxBpDJNznl3q7ZZ8w
ULzjCfuzfdTM3bC4YUPxB9JG1sm2O8NVaSaJdOWF0PHBRgojWuGrFCoTiqfGcukGthGa6paVtUl0
Pn2BnMnwpUsTZ47bUsDAcIXXXQixzElO4ilikEeZHngPJP9ZiOCGOiU27oeohuVZwN8io5ZYhKNV
hzRjAlzAfJg7NqXSsH5M2WfclyjA9FNKysocUcMoEu+PSSEgM51v+70w0FXYKn75wGX8Ft5OyaAu
0iJF+Wbfth2A1qURBKnFDgUPQhQgi0YjyVukzLPOpQQoXNIuowVouQl8er3csaST4mNzdzCw1CjI
v8dge8E5hm1L0II/RBko5R3ykZmiRff6pMOvet+Aq1tV3E5TUTHzuyg1ROU0J50bamITlk8THfBq
sB/fv/2s+8YVNGq0CVlwzseHViSYUpiQyrrOu+jUGW2DbHVsxlq31bfq0T4wMb1nd5N4OvwxCZxF
lsMdM9KkEMy/A4cDE2u+e2ALIV7Wc97yPqw0/q0LUy+38jYsRXxjaL3f+yfcBAsKg7yqP9JT0lIx
5RRppT1KuveVU7VrICuwAAWcXGyxISrpVLpi8pHoOwohXXgdpW3pyAsXmAm1DIWwAGS2K3sDiSxu
FopaPjJQy5oPN4vK6tuJFqvzBb5SzQEWUOOnpq8EbvpRf78ARE/UI44DV5u1EGoEjZaMYqzPeRzH
W08oVWzmwrs+84YizjhyfmwMRYzDazOO1oG26xFQeuSb1BOKk1Cm/aGu+Knz339JzpIJ0alohd1D
UZ3x9g5UC3nIVlc+IO8f3u+9VXmAaY/WDIhxMx0Q33XGioLtCepv6KwVVHZLgsbHsrkH1niTuCpK
98lcYmYrovnLHinkWTMzOWK6YTiDoqGtCpJzWVIZhPjg/v/2y4GpbnUKprpaXhIaSOTakf2veJYH
CeLX7fFTvhoMzG68GJIB1BSVEccIcxgWYksTnwL8spETWe7/IAyX7Llh6Oj7ort42uXTxhWE3dvM
m6iezG0KtnECpE59jbwniMeAUyQ5f0lRSjKB+GUtO7X3Azra2wovcUJB75uGW0wdCG7YmfLDcvEF
AVAxSRuEOkvx9PXYOcMSQyc/iZxzhkO/RoSm0gu4jTN0NO8C7IqSfrU+Hk+632OLCdkdtR7a35F6
y8uhisenInFbVygampBK7wk08RKEib/lvjLW6ckLNFel4a+ZKTEB1uFuH+uZhirIOP1nONKys9Bo
mQN6ZirBUq0+4WKig/WO3vVLoV/r7H0ftLP1er2CSeDfHvy6PXf8i+6TP/duAOFO6F956TrvqVvM
eCbGKH3VqNVFfUBPlRXR1VWJve8NTBloKSE4txUnr+TqcYnNnt381TA08MuYcC2KfbpLx6jj8aBA
r62HOjYCFrQy33jZrEGjlerO7XKOcmylIbKrXwmDmVe16Yh8hDBopW3QWjNnXY3lg9b6F3uCEhpZ
JO0lFiQq0doq1PFF6LZCqa9mA+QaNCrTdwPOhpsDLXIRIa4nQOXsL5LlXsiv7hRJguYFrHjnw7j6
kPe1GwsRsITm0q4LHO/tTW73DZVqJBnWzFq7gdzO/2DtYqFD/O7dUBrYnExqyUzTdoXF4a7D7Mz+
U0rxvcWxenyIVsRBBMzVtXa7cKrQ52Z4BZrShIH8IRX+u1MULop1lBV3z342oAsbVc4067I349nA
zEQjsiincnpCJtQt36B5LJxK+GNVuBPqPP9UBg8thK2SVu3LVdupLPSTrgmPsm2TdCJJ5fgVBVBO
i6UJiXf5z9O2fdI7RDHeWsYMC8Eu+TNIwBavGLYz/TX/fQ/8sMcvFBzpApZLVKn/yuguX17FU4fE
jHS82em9sT94uZpXD7XAf9heHgAtu4eCcKBmJljlOudUoDPaHkFcRnWjjrN/adreCBYZq4oDJcaA
tk0AzlAxcPTUjCVxfm7vo7XrO44W6x1WURaQCc7GFZS/zlojOxhEInTj6ofTWOL7oMU1iAz13yki
LuSb8EPsIxwxDU1M9ael+eLK2pBUZD2um7ka2OpQk2NkDIa5F5KJ0vN7Qe1REnw9sZdIQHub1Hcp
xHZtsRJnHOFBf0Cp8FuLTiXc+XQDS1F+Ov0Ypw8ens7te/58OYOmD+dPLuW0deAITeyJPPeiM9le
l5h/G2Pv7ZuK7TQdSP3ohx6Kqzko682cWv9qCKFr3j7NTfbZWupjS2raONyBiQuiI3zq/ihKWM9k
T5tz0kXw16dBlTnSjbqBZiFGsMrNojufurcFsrlvEkV29/ox3jE/wAKOEjHos9W8dDd6OnFChadX
E8LBNqZGao+tMQDCcGM6SWwrSPRltGWiZiQZqSgTARXrjSaP539TYM4p4IBBkcb5+r4OQlLThIYs
pLh8/x5LtC74rk2N7cr/i6YE15GHy8w7CH9a9v1gIwYVNOhFp+J6cQYdyMqjfY4nIXkD3tKZi+JL
413XlFVKL4fr1LmyRTTMPKdtofibEzVAf+0TVDM8Ex7n14/22iEG4U+KB0HgmrA85bnd5agqVxI6
jYxCL9ULd/zKO9npRpInSEZG48Zx7nkHrmitveym+bbTcucbfvGB32im1++lz8igN8tiLApuvqDY
fGaT0RCdKbwI9u/CTOa62Iwr1U+Jl4MeBOXzP7IPcNsorsDnAODop9yB+ja34jIUAFhYqP+WAck+
/nYk/HZEo4DTXiSeOpaIJzLxMyJzYVSimBi9E4zkqw6grQZGbWleRgth4YmXwnBXR5unk7fz5Uo2
u3JQt/VH53MqO3e77Z5CKsMV5zF7eRl6bxNwyqsLROugOcM/9B1QtQ8dgIqJz/qv5+Xw+SGJxBBe
mX2EldM2M3lhDiQ/RFBFVP5DRiZmybTLZxmxpgzfjmEN09+KHz84CA8f1iHO1PANBQnnbEGoZiQD
fLBBQRxTrf1OZ/JpSrQhSibt2WMyU2s6mCmoi8buSwHQLlerYGWTRDwIc/7OCIPxnQjo2AqIehtC
awYDg4+WjHdl/E9j+paxTzJ6kGkxXZmKL0zlljK1fy4xnleB/ggxwRveGrXSGHugKnDmns9HP5Zx
67OKEECiHv10hK+WTs4W6HJTtyma4/njq9cEUNniGW9NvCwkyG/3LvuzO5GROO/RIRAaZaiSsQF/
BNIrhsF9CPA99AYH9qIvYEY6SB7tDr8JUukBK93eEOpHq3TxyMqyihbqhwUHVcpOcHuSXSEpMjCu
qNLnmrhaET7/w34hdWFRXybMV4Q3ucZMm5XqR+lgVPde/zkFL9q+DN2KYc4G+70KI6rMClPeQ+Xb
jlNfNMjJ5jqAio+TuPcGaMUzAt03pmBZJz4GPGo8aVTEkEMY7lgmdbLoO5xgPoHW9BhpRtXhTfOO
htxVX944JuCrnrknfMb7Kiikt6UEEmahjnNzl4Zm5uvL+txBeJNv7aKzVRVeJzL+cJmXuW5J/5Me
komiHGNsHNK0NMpjiPf7l2BDgp1Euvv0WD5WV4oesNOAzzXTt/mma2uqSyK8YWCKdxj+69rwfrwY
cXyJMGqMG/16VXMik3CTZ4lGi4gECazsnwekmPylSEM3IiMAtjOxuJaYwrdJz43ObOTKjtD/ignN
ENZ8bBabxF7CkM0gG2wWdMl16a5J/QMZFIBz4iwEtn9YiBy1XQldPfm017PFvJo0EhcilDbVsRfv
9PHr/DlmTJFyTV75Y+5qAOosUyiz/dYM97Kx4HDnRqwbXisG7LVLrDmxgbZSci0bn85/uhBZialz
gy79GuO1AhfdQYV6xgEwfzl/J1bG30szjWk0GQMSQkloaWsPo8qg15Y2OetrTNWOUj72QZSVTOGu
J/WE0tCqbQYW3fWXOVU58DFGn+wtN9tc4kF/94v3Q24vkVbREBCGPFI3AMLrObONQudzA2qvKzeS
WOLsd2cknwl1Kr3OkxxGmvqhTdoyqc3TuTIS+ZQFzO3OcccqL8sFKUGpAYNhremJuIdX9mWIc17F
sPyM2y0FNEIlEsNI/hsPpH73ACPJAK83GtfqBV5T1d33h1wwhJ02gyH3rVIZS1XWKqBQqAlLMSTS
dY5mDuyi2HJgDOjOfxB6UWOmrrrHHpCxvBFNiUTj5NUpDcIuylTMZwyvQ3UF1pqBz37FoEkwemzT
75dTSJO4N0pqAzY0PS/+y4r/Difttp0HD9I3EKuO0KC0Pn9s4Af0mHpncOPL9sNaav+2AJVEW1/U
fu0utrZMogreuCc6fVUoKEyuj1kAxLwkjGm/Ya4ZnXezBMX73iXhNnv29Q2T5iHOhY9uLgoeE0fr
ZIivJ1wV53kJU3RHUpDTLk9tHj9uh4Ksifbs1+n64EVL7ZvlgqRr6wE5OS2M743ulv+fVcCIFKxp
1qHr3usLbB1K26I01UQ3fAHNhc8dkH9UsgZr79s8j7tMU6wyk7PQK/sTNtwS1rbkP/IY+3YVKZXE
fNInZXP3n7UnOqBpA5xRUfLlddYP03ivqKD8+SH3e785uQpicM04LW78KjtafwRx/vmOj8gsEgA1
bosiKWRae7OxQfLILp0e8xqbjzQa5U+N9JKdf8JxH5JCW3nYIGxV+crG6JbV39GUGpYOS6DBQRz6
UiM9KJ6axhaj/L04PqPHwPnT7I3VVWEQH34pII6yDaNCyRBR+Oeme66V9JBNiU6JTMPPOOOC/Bm1
hVKt50nERGw4pk+GwETLHaEPkUg/BlFxQRLtmizVHKll4pUbQpKw1ecl87jwEZyYMEIdmHV7PRG3
XLcRBMQF2APBlfHjYEnysUfpf7KaqpQq4+Q3wRhg2SbzFgAzCo62E9/Gpuod/PCmD7qY8tTY9Wkc
jmQwmfp3ynji6nHCVmbPEi8DzZy1SkaGTTmN/6C+T7ZbXUsjZqWrn9gvpKkOYoXQCBk4J70Pax0v
jmcqWG84SCsMDsYm7IlRyP6RdR78pXox1qczDKBh334ydJtOm7KiPj77frQ99aWx/GVe5nL5EsyS
lGpqadVY9Jk3PvNFJZeN+UVZtVkF5Pm7gjg6adjpwHN3Ul80QX4vTUmoG72DMONCt09z7q1NUSgA
5GDlHlfkD8SDT9wbhLrJPXHpgYxwvtIU8NksjntpdaH3801WZ/jhzMq9fEbbThLBbn5ZrKneq9sr
TxK1MEx2crbcoSbt2OszG8rcxccxH+2awzymFWQtsLiA9bD3WHsI1hKo/AHHjty6IIML0XpTEr9g
tj3JPn1Im7et610LfIX/Ee+T7xJ8XwnNEV1TAYn5Bl+zutcEJFnzMqKOC3+xTY4Ar8M9rrD6y98W
ecBa6xxPzuHcYmd6puEeKvRGJ8IxRNah6lUdkrqydPNIzODK/ssQk4bVnWMagKUvP8Mn5JzU2JJT
ezIdWWf5l5TMgimoQaihD+RVG16Vu8QRLAQ2Kc9UoJrOhSYHEfd/YVH6TrIXXtzIzC9vRh3mVLYO
9imCK01xMlEmp0651gaCa8TTEDfgQsQ0W/WPvH3GuB9IewoHWLZAo+1b2JDABz2vB6fmSgPohKjc
b1JYpm4OOnSZwTleYJkfRyJZRRAMv54U71toPkJtPQlWIPam68Dd+qr5vcumUui+2tlzw0cZcfgw
SZH+I/gVAo7ic59nUKOUzUi03V9suy/0x31xR1XIDRffvdylmvfk5l2ZmvZu+J5yECV2K7M/De7b
TniBL8eLmNtmIX1yLY1IMXb8U1sUif06GCEx8ULPC2K3NgGprphunGjEM1xDTgz9NKn+UYj49Z3D
3nS+7YuivKJ9TqV6e5K0NgBcd24KOhdoHFc3CzJgfZTSUjJzZbWv1Pv+ZfIsx+yRSdh+Q1Qf7Skf
capoezafjX0/00ZBD6HL7Ul+xDLdRh08oCzVrupQsDRCOlT3pxpi3w71fT9KBFg5dhkUSICab53j
m3MalKF+BsANwwTDgIa6/zn7JM+pEHiGQbKk7CbjeW/nBNfmtC9L5ONehtkJu0VsEuekmqHcV6Ql
sBV5cMMqyUBEkZr8QtdTvByv9CPjEdhYq7i2mHkDdLzF+8vgmk5NAqnDAN9Zujk+iBcLN82EBbUU
T8YjDH3RK92q+5y0tyMgqZkf51aRuEDZDxknIdJUfODznolRIbMD1VCIAWZ+NE6mvyqhlyFJBpoN
tuhcVpCf+AG4Z02AlxTUMsaXQ/pF2rmK5v+/ElTh4m1tonbaCoBA3DtKjJy7zfO7QCPY+QAcCCo3
U25Me1fXJ7xhKC5yXfum7qFDMg70gCeiNM4CKSxe9ZEMGvvBvndknqH+Zrz5SU6j9sYXJvpTm4B4
tkyyYgaz5BC4U5ZMnI22Cr/EBVos+WBsvMGBGaCU7McJGdKC+HPDPijAyxKyy9WF/5ThV2ZW44ly
8hJrlkceo+MuAZy0HftxQU1uh9vf98/VV3HKJnfuec1v89IZcAzogHMhhwmBkseJEemkJFfsws8g
ssngeernGhKNR6HlR2Y3O6iurbB2NzSgaUI32eygc9TXz0F1j1ZZezT7EhZ4VkCYHpAaI29K6OLO
Tf9PsIrfqCJVFwuyi04b+iyyJqmyDau5sAEh+WQmysW3JFbRZphmMXf6pznNMcylwXTVPIn3952A
2KwNswPcNY9EbNb2NmoNIFLerwldObkQLNsrcFB2eoNexLt/2KpliTlv3g1bg6DVxpNUJcwavH9z
4Pd8++Inx5oLviYBxlepAgvvvcLird0z5VpvNfR+u70cpZNqWh7G53VckJ6JkEId0YKfY07LDcDe
D9ofCblXwatK0hMkNza3/7PE9s9FpGFZIM6WZY6w48uf2BsFaXmCgapcJOIhM8+ksSIFXoNcSs/J
O5LrCFZn+UBQwLvzRdmcvk9Z8F+dN1TnnOnZXhWCJzdhLM/RQJyYbJzhn09WEou+Eta+Ne5fu8FU
C3i8oYDFydRRNsakEB2XZXgd1qv1alwWpZhY+vaEiZwzdiA+jD6oAYo2iKAKkNtm+3arhVIz9Ao7
hBch9eFyrPSpnoKxEV5f5zcmwDajBd3gddaX3NXqKlXYAuZ663cbX4K0g9uK+N/9IUXe7f+6477g
vXLTxGnTmGTYepCAk4SCuxM9+81P3Z1+jPjoLtBM887dwFUtRzkxfDtykFsOKpbupLQ7Ajltfu3s
XIIEznJvERHoLlXnTefh0x32g2Nsz0oB74h0k4VEuKE4HcX9aJ/e9LirS5h7xF1F4Y2eWsyuHiL3
KCdCvw8kcKbsroEXmFIqxprGJ89ERoGATD7ic+3gawm8miHdpZu5W5lTWvwFfLgNrrhHvYbo+6iq
+BFdcqqyrQhPK5bWLghuIZXVMfh8Y9zIQFxuUwcXeob+2ewApymKLd6U+E0fmJvHNMIdn8PoDAif
kOY3IkUrR/q/L8uHuFiLRRM3M4ih1KFH1hSO4/2l/Te7DzRjV9bG/s07E+ycsKtyfTLRMkJpJUPS
s7nEcrZ+WBHT64fROy17iaHeSOdzLcu/1+IWZhTHh8+KzD50Vp84Dcgtf/D/m5AwJLzCMTDw2PUP
by+/Vh12editEGLo48nPPfetUdoy9FRiU3N+RXvcmYhkvUvvB1mGHGcqzmkk1xTVOuvb6YqDifcw
6xD2j9CcAwRBxWdvYys6m/+VEY7f0c9khCq3SYFjd+IxEBmK3ah9N5KOtucsL2/zGgkm6rU+Fc0j
RQMMeVW1VbYj6o1Sk/lQ1cMv9SeMny+wW0b+Zm+1HQtxRkCoZKk/He8218BeRqfO3kdlWTLfwqkU
nfW2E30x5OR6rnW3ALQq9OxnB/yirZbo/sc6W+8pl0YMWYDaDBr7V9+Edja1SZT3xCcShNxLtV9Z
dxyKd1vgm8/oKjylBgi50Cqn10dUi4jGoEwH4iLz9Fxnaq1Nh3oE29FUO0FTtyCo2KAo40TGxmFP
jDgYoflQsWHh/DpP69zxr+g1+ITBMpoVCJj5zh5Gb+bnsEt/Fi1NqEj/X53oU9D8O+z+QgSfvNWY
N3yuvj/e2iuhlMH0qVPHj23qgTE4b0vfrxU8VHyFH+ljq/4SQs7OQ2Gnye2NjOPTUxfBILQSUQl+
WhwsA2z5TTlVltRs4/w74KZ/L/xwHIQWu7YYA+8thYEziNOjX2/2bvnV6xbN15yrkhFWZwkwYfOC
E25XioGdorYI3EdBybwUzGYH8tLQXuFsEYI/tkzu/8PeFPsXPVIAz1QKrC8kpUEMCKSmy9SOomQx
3vLKSn5k9y2QHor4+GrcH5k2C1KaB4cnDN8liA5jtrMFbPXpGFyUU6w5ZLKmkBCKcl5uxjK5MCYd
qWVtvqqF8olGP9gybGdP3izbp/3aVynvVnMfETQvSracygUacIAI5BUIwgdrjqXpfyOdLaHW1R3Q
ZNVawrfMZRckQpxkawZuMJyg+0t1Szif0UxlWRzWl2A/jUvDp6GqqNjdGGjB9ccCzQLbNxJf0Wcj
Ap5wC1ArYRBwrwTS7XPTwiIp8GmmA9OF69euAtcVd1puGyNEXoikP7GtngNKbtfGcRPTSCJNrjsR
5q8zvwfR8AT/2G9NM6j5a50nlDyG4Sx74wsFJ1HEvQ41dRkq3oRCL1F2YjFDX5rd7Fo+sEToRrpi
Eg/QeJUuR36AINb03Ie4k5FGHNyfnM9kJBqFMpQSHizLMC8qcLJO9ErLVQZ6IT6bxDaXV9pRRG7E
AX54y3TZ6/7lmQeGN5EDRzF+V3XkS7PVx5HDlMb4Ep+24FpMoq95kEELj0zPZ11Lqok9NMLIPFTc
pFkgrxdEvKRs16lcdeyMT/tX9STZjFuVF/1g5ULhrmOC8ZPhS/qL8z3J/g6RFfaErSNg8t3lMDUw
BpddNz+DsD6X/mQCykGJuFCVVPbewCxscKBKG0uA7lcEtcTX1YD3sn2TC1E+DM8lALIzdTOqy1Hr
JOKCyMwmRgi0c1aQraNUcnHj9XX1QZO40hB5EitQeiSATBjRBVYr7+koYWAceOHq2UlIffqyO7gk
KXLfE2b6bICb6MHzL95uyT9MzA/cwZAcYGeh4taCviM1vI8NyJ6p7eSRF9BFQCzfCok5gfyaa5dy
gZL2dSr8FLAjrD+VgquZJYykLIk0ad1B/SVkfnn6zTOY4cjeTc5Ge4a/Ehlrph70R9jzi2O45g8V
1c5gEKYOV56QA2Jz+wrW8yWcW0CL1UoJc/z9gSPlC90eNkEg5OIToGEcgzvIxjvkHLHHZDPKhEhE
YywuZ7KEzyKFYTkIpjxSCzhFYZa+aBTkjlrXijaCiDcP+p/Vfc0onCo0H64nT/XE38y/P0GEzrnB
5/1XD8XCBfDgitmMKRqwmHSgKLeRVReptNm1mvbofxvD128pmsNHrl0InGGIkXszVXRGn/uUKx3n
RG4Q52bukwxLjhQgSbuigfTS+rhUR6ND7px3Nm9sl3Y2lNZ6QymMjLEz9XoPIj4B7OVZQAm1nQ1K
qgdeVBctoFVtCg56B5l5vFs+nc07lMMP5pbsujpcIBoAsgGk4gNK9yVzE9QE+dm6x54veCquNQ/n
0npqUIn7ipi9rJdXJmhU/fAmatyNdkpSLRqGtkMpM+RzlzCl1xCMYqcalVJqvD9Q1Ys2Ggn7iESu
FJruMHDnzEbrlLK5j5Z4zaRSvXe+TyWH4ejD9x/5Ixna0aNuqZnk+o4Deok7YIBICuj8OvHtdx1B
aEJfSM7T0b2chTPyP0xu+loiZsYg8Ip5p0CfXviarNpQc50nFFP+MDAV/svjV3xfm5mFz9AXRuPs
YSs6EHy+41yQWrWVK/s7SaJogaAk4EdW3IJ/wS+ssCapwy/AeOhblbuoovl1bkWza5C3WY8/6b6l
PVt7vPcxUXJzJ2/HWQc2rhDQdOEg65sbdhATGc95JATA40RNdjearhR5Wcx8SD8oQr/k7nMMNCm6
QGIs8tTC3cmQ9IrkSQuer0vo27uUkNgzi9gtJKZpjUbWru3yoQ+ws0BCLFV6vsEiMJP4DC2CP3Bd
8c7w2+73GRJIFXE4v4p71ouqmN2yRgic5eHyCaPC3+ClXwDU2Qtg+/vGxeiTwnmWyc5xK5otSPyZ
WIdagFg5dbQQ5ceYBz2X0tCOixbbGqS9Q2eOPFci9hu7NkpAgxKC4s1DplhYxh5KFj06cwxoX8c7
IXOakRP/DpExTpqsFy36QnMUBbH8xg9qx3y8pezGemYJskgI6DozpCbzNx/2ETSGWiOaBBiN6Yhg
HY4D85TCLCzN/FZJBialR7ka2cr5Hi47MQPn62QBBLEWDmF5+HdW3N0LZk5ctgsRHpV89121992B
PAdn/hM02fUWrzs5hnNHak8WT2oF51fsy+8DFp84ACSu249Lexx61LxkxcZIDCHsewZ7W0oMvTyp
KUzbdRCy9D87TZoRi7xynvlf29MmgzT0NOMVxusFwkzPPwC9Sa3vwsTH4OKR5ilRIq6XkR4pqnI4
1XoTwYEN7jtzCT2JvIbTdQrGxmD5bq4beCsy0WchZ7nMP8Bs2AHjvKjgGS2uiDgKpIJzUODbbTg1
nyHadmVmPprepAbI9Y25ykbbM/qUIr11f6vJBIKuyCrtYJYeylRH5sRdsm4XWlFpXkGNpqG8pb69
lpNTzdTRKgcfeTRgpjZfvA7mOU817owoXmxGGkTmcdp8QH+SpWoy6hoHyqxJMjbx8JYj/euWtQgR
ZCz9lK/aGsSdRWLeONPfakgvz1PmxoxX44UD5CFy8w5CDsv4dRpgbdwc6tXJMX8bSy7HgV8GvsDo
ebM35zPbhi2+bZ7ZuhK4kbnhW+t1pwVSTRLUEKKrEdFo6pHB8kf+NuIZoc5B1IKI6hffOjEpeBUR
vYua/8pjLVLf+nAjFF2Cl9uzNTheRQa0BT/GRf4/XwFfT4klQckRnH/F1NrYtgGkBSSt5jsrhO1b
9r4L0xJwmYrJ6OAB+uE1ATilYHyUvoF8d9JJuweRGtSpY8HpsfGW/iXUO9D2wwOGeYWhyDArHN5k
bNoJ2V30ZDwfjutZKyqGxm2sLLne3Lo8Dz5RnY6wB+i3O5c+Ne0yfvp3lf9uBfAukzBwz4X5ZOSp
atJ4+0g0IPZoXrNhQPE0u+JljZ3nDPS9UAACWZqjvk8GJZ0KnhATSCYJ1h0BDPKEUwYG7XlVI3kd
6352Uj9j1WWaRtRn9zdMFuCe7oSqTmo42mpsHdT2YsviOZVFi5MheGr1Vn+6jL8iqYUWj6ArLGxg
dM1KuLWi+EeQYsTdpHuty42jGrJH7sYYLsHRsr2iasOtsmhLf6qcKtPVXApwvuNbdQz0Yn4RCyWh
PLFyqT34kDZhqWhgWK5qkw6wzmRrkkKR9JrWahWCQthakNzcM5P3L2qpk7IlpXEHs+QruMSXkfmY
VhREZCgRY4IWbQuCkdCJDzjXSmLRdDd5pSFijg+nH14N0b3ouSrfdc/vawyWJHNxYgz5+xphWBjd
zT18r1s40yQWKBFGpCADg0WHuBSpwGdbhhdeUR2kgm9UFeY/yfihvB563WXBI8TGvzIUVfvp3Ln+
Iq1vAGpHJyvM1yAKf0pZaNpSXqt1SEomXNGYRqgtOw6umSF5chECqn665Y1di7vGDp+3omRFpUVB
CvaUlkocAjf9Y1iocH7smOxNt6ilTZY8+8jSmWigng7MhJSQY//r8iRDHuJWI0JuZDjsq61zGnlc
PKg8NtE4gvESwWSmIJhBRIhkca5dDYNgiP9b+PekjrNB/tyJSTVHaNqG2NElt4/oMxSjFmJ/IlkT
bylyPB8J2+5/qs7rLVhOoMWo/ZAnHELBN+ewl5V9Ht55ttiPMijns7lGHp+E6YjCQLjkbdvXW4wj
Ys8TMdmqPhnYAr+B42v8UD/THyKRWunJxAcF0bt80QE57ABJqapPJdlI0iprYwRvncu7wEwKWAGn
Al6MAB8dJ8id7wZgRObYuhmB4GGd0MvCbt0gaQpMddPYxSXKzeQkWyoJNF3QQ6TCFrzn/QUXYvUZ
7C7LG0pRHVSXUIETuS7+f6IVMw8aGKBS2hVNwvSaITCAyojmYjsLoTmQdWBR7rpkscX8q7LGGO8z
lsDClzL6xLEjgHT6bCSRUw9RtRVh9FL7hLFmj4NvkDQpH5loo55e8xSrY4vv5+pkv22OC4vHjvfv
ybqjHkhqmq3VwnPXPMS05V1k2uFrnp3782zrQoejWTEYkXWwYf31abraqF0A/SluYrzVCwRxcTTy
wUQPWnMSiKQPGvvS8aEFzZHimlUIBZW2fdO2DRKEz4VgbyNyTbMyy0iA0aIK6VRwiQ/WlJi/RraI
FA7D4iBcSZCuKzFVFNYgcfjjTcydPTAK4WHW4/dBQ95TN/Bk4uHKnaNq96NtZqni2bWsh1ki2Bu/
nd5LHAmcZsEzlmxnjxexO/WuQse1JetQpoSsken4mRr1jCUTlouJhMfA1xinMFGaOMb6acrlmrFF
juScOdWyTUAjVYNox/QL0RONH2gUxAEvNJu3PB3N+KD84nRAmYnDxXj2L5Gp8C6YuUuk32shx7vI
xrmYIcV5iRGBDOQiNUBEdNNtW3u9rQ2VjRBi9WKrqGjq6bQ4eDP6MT1919bGptbSfD49Uzq1zWB5
UDXrjFxE9umg3NfrDIJvSkrp+35MXHd2A6C/N5DgD7Jl70uZNcrBYevTxD/il43C8xHu19Kk+VqK
6UT279ELCHi746SXLf7ausqJb6iKPdudrIpbHhghV8VT0ARmdPWCemuenGbTKDEp2ANxIdC1YAyp
pcI/0cpeXLAoNQQuQ0tewRp/J9tgKGBRKq/3bkcGhXTsIYIFFjWVoLaNSe/Ntx4VXK3ysEr0zu5Y
LN7XgZDbT8jaKOG2TJfXSwel/eARbrq1P2ORubUI9pgoujT3Mp7XKI22/xhATBQYu6/Jsc66VTLk
UD2fsGiWeDI4VNbI11Y+O85tW49TTp2j43JmoRsis3jiTd7KNGLSyFAuoxYSHnC25luADTuqlu2O
QbgAtkEKFt5vcDy54mrMDJ0Oqw/cCpYVyNebk08tDgXTvkkme46cZLT0Q9FE+VPpJlRkA7BvzNOS
+7kHY3q0/m/CkYyIXSGeg/sHSiM8SBLjVH5vwVUi/5f+Snw45z0JQ61jzeAWTFGHVgWwyBX8re3V
mInImJvpEQK9fXsRwgfcwUENYsZ9sWciNRrbAFefAsxwf7sOuiPgQM3FYebpPFpwfkqjBgYC57jt
5IWorZpfnHJ3we6ee/FAQtloxub38eEG1tV1XCcPhvmCMMAHceT18oG3PdM2iGPcqGQPKfEA3Ro/
bxyjx5BLshebJFNeCAImZ+wnbSBqajfjQRcLPvYfrffMna+o4TV/A2X/uzD+m3on5gOqsuaiNIMp
09lgE9QV0OOGHxkyjeyyKqICQ1wNpP/Dx1ScK7RXane1HZPpzUuTrOb+EcqysI9UI2rxoDBDHiMP
FzyyXF4xUlsNKXOPrZAKGJIq6n1omSgdx7xhsRKHM/SCL0WFpovIHxi0BeDr2YzozzTksR1N0BLM
soOD6wM1ucJnxrHkP1wM2DfB/KR7QiSvZFcQep7Vk3WrLZaWkf/VHFCaZ8UfHEBYGuWhzCRaoDlo
JgNeIJLaJvi6dZqNlNp3dj24bLCRjQT9tLa53z6xSTTryLOaTWVorxoN6Z+bPZCAGE5zRhdaK7ge
WMAAx55vT7Nn5z6tYC2wK65RihNeg6D/OIusKyvyyLZIhsA36KvokIZakFxQ25GGj1rbQtY/Gqxg
P3Dyjw7eaHjM1/JaqNiriY44GsHjXxx4di35xSg24USYMtJeaEIJLSflIiNcSC8mL5t1nbJ8ywdY
VLdrGgrO1ljWxWtOjPtJY2ef92U/E/XCzWns/lIzb12qr5guhV6kzWZLqEXzKd2ARs691LprKcQH
H8FvlyJvjRUbVrkNKcLoccFgVHs9nUBdzjvkpOdp3T1aQ6yQ4I9Kh5HLfpxpJr48NAKhezI2IiPi
FPl/HSPMAVGDWuo55pAhAJhnhJ7a6hpVe3wvLsPZVSvyjZF7wP10v/3LcEhZHbAKV2/3GPMfe1kQ
Qsufr27PKAOgpQ4NQP/aSE6Jj6dzeFZOXEH7vL09+i/Pd1lc1skdUphr3dXEdg3hGBDA9yIKFjp3
NBp0OwR9fs7Gaf0Rwx5aNSxhLM5klEnyFMxaWWUud3u4OJVpN5PB02jjdXkoXeZcm7YKZtUMFc7D
Wj1Lcnyocv6zsK2uAU95CtlS5t1V0lPtjam2QQEsNpWiiY0DmZrSB97AnOShUN5hBUxCZviClseK
0k6CS39cFgNaPfKJvW1CvuhaqIQrazmEXuoBdbzb+v+vVBNSX1KKZjC1gt3hNthbd7NwkfmVtiae
3KQhHwoZcxP00zFMA90VF3/OdGG9S8VFPTHFHbDoXJu5d6Wr4devM3h8RBUfLcMHmS4aPTydi19v
YnGggTvGar+jgo9wTSXn1TF975bBLFlRuueUj0XEm8FBmJajQxcQTu1s935JeQRzIjMVFgovn82k
+eGS5QImchNbr5DnIkhj8yZrSLqwOkRCTjDUYg7LtOH3UaHRdYnSpu2i3MmT4OW6t8jAWZo7Cu9A
JiZupLCT1Oz/87Wkui3VcvBQGWpzSAMM9GEIkJDpc32b3dgG/6pT9ZsZQ0NIfqB/phiCARvLh8Ph
z6+QsoqqCkDwCv8zvxbkWN9xqiZF14QCKx52v+5PsksZjGzwt2Ojts82IMWcbcTNpVS1ko8xJn/5
zp2vPpAbiavKSAxG+Yxvw5/W2K0upFJAYmRbSc2W/ZI4v7Nxt3Z9h4B+Zj7BhuwFpejad61q0mpp
u0XsXarYX1fogVvgFNL11epsSif4qB6Fv+BB2pRNYP5E8KPqVXgoiWo8YUsibA8BIejsLWb3F5gj
Mu9qGFJk/wVX1ig50hSbgYwocSXmsLVbfNc2z5uazkR1IdtXW8jhsjdHNBZ1xSLrPQwF6Zlu2lp2
KcUpzd1xRA+yVP0QUbeQ421Y8Fk5f5TQufn7mtICKW6cG5qNlhEMoDdCaaGLF462A80Gu2qTsT82
cr76f9ckDSc6b1n7rzgX296D4n+OpOWtqN68VfjT1f6B75GM4lo0fqDeJ3QGanJf7+DsGfGS4+hw
xIXj8h8/6tev8J7MOwyYjeYQCcBPBe+6avMaoNk5AspUgmOwhlt2rZ57KnGhRJlgJbmRgB/3MbVU
jifUiuvCLXkLGvB9u+TOhF+t12+LMdSymhrPlxxs6ejKdghGdZYfr8AGKET0zebG/oZ0u1GyB/Bp
wgu64Juw/gT7QsiYMLosTCSvHiVQ7mJmhqxeUZZ0D1gBaXr9uaOrscCZt7Ijj6qdMRrAlKjb66H7
sjWGfQva8T5xznu+Hnr8zraHwMCxArkdiiwlIYLZ9tlrKCCzBTOtV1Q+Lr2s751Xld1wL3vm/DS0
dcvaT8DHJrU0Un2t/FAa3oq82DH1t70E2qLx4yC69kG/RKzDoFuMOoALYZYNhOXyFoHUONhm4390
jIneEiC896v3nxHGIWweLup0P+rVTOcYmaQ+tpgtxxNlD1aLGziVmNRyf/H5RHVO+JmXKIzUEoUv
fNOxTxLy4AHvtJRqG38FdEd8dg36h1kUIL3URxHuyU84QkHdv06pweg9/VlUWPQHSWgEObBuZS0h
1VikXA3XdSlAi3fhoA8wCz2z47x/xXdcukl7VKZJ+LDqzYlF4YqRS4kNxvJdHbbHX/xZt79AmtwZ
r4ogIG2HMJ9SkKkkXuYvP+B5rXehsHERXL+vEX9AJffQUWGb0aC91YoQEXA3Xiix96flSArEBhNy
O2GjhoncM39GbMvJH14Lk5L8bm6/sLZzkcOuLIYq0YuXrSxGxTLBZstlfm9h5ez/lWQTAzDgQOc7
tjZJ4sdNf7v2YSXfeIqxe14bGi8mPZzqACoK74wrmQar+QAg7l8pg/Mvb525ew4uEtwZR0xFK00H
0RI43yambsTv+Ij3zR7Gu0I3LYEG6nH1g3jNw0bzHVtotEbhKAczdOTy6meg3S2JaLl4o+/MpJ7Q
5apub5okkUik8UxlPVI5h0q/gPS/8WFH6XXZAK4S4vUuOBvwM/fSftOiimbVcefwc0yJa5jL0C+8
g7BOVfZP0UrWizZ61ZxHTNdA7k73c9UoeZ6x/1CI5v4z3fBjOiXQnJX+nO0nlFwBQDrDOrBdRHOD
VsaXNKmYDGyhqJLBfEKh8i6UW7cVbfDdmxVaEzeW7twNi3J0KbkFQkysK2x+M8KPDwc+2Io2t+Bi
p8Sc4zPqMK5V+ZZvJk6tNBwlCW2dYk5lswONgE0fzTQWlhcvOd/ILjeVL9OfCfKGu8H1/KftlxdD
BPCq3eG4mqRc5P4JEFFrXhmrcSr39N2FiRf+ZY/pbveol7cjHq8Ygnjp0Mxkc+vz5Nb2m6Tc0Mkt
p9dDyKHO4RNoYPRwgXXgKbMbpLD8sFJZyssqjPulCnf5MY2NoEvYSD6bPv921C0yt7mw8FD/SJ0U
RxyqtFodl+lH1GD3hYJztmF+4JUYyw7j/jUIYpCH+foNgTGq1bxwUA+w4JXSGX1pAODCyRMuNDRl
X0xp4SkEUr+Ia3t0jdpKUI3i1GXrYnjq3FE1GMffDqFM/5JBqKRL3QB3heroeyqrFjJVMrDP6TXd
VaVRvg3uwfxcGF8raB6AOJTB9EU3lbhbzd7HCVUphNsHDoTetrpzPl1OYnPxaDh8vTI6AUPS4H/B
3EJw2bRjPq8DPS+ajOAqkFNT6B/MN4H06qcBldFRTzZulgwtkoQc/PvuGM7gXSpMhrkIJ2CK4pAd
zSJnm6jSmioQBOlpnj6c3Q9mgaUiTMiWChubT8KSdHLpq2rceqwpmawrDhv3hPzaZ3MZRdUIuaD/
2aK1J00HNb3MKpE6CadAkxC42I8rTGIk1raN+FcdW+0FV4XEj+lw3jB/aNd1K+eRBVjfM/IZQmou
UgpC3C7TX9NNwHxl+nZZ38XiAAB0bonz1x9Dg6iOo3h4bHHzFGdWnxKWBEEzV4GOL7k4D0VVce0d
RjL4C3W6KwPi54F9L3lO7QEmP/VUaMtC4vixG/T8w02iWbTwty1X4mTl9qeeKgNQiVs3sSJm4O1t
/8zqgJL6xodoauUBSjuAE258RKzQdmuwgtQOWm0R4ZeIlsjwIoyIM/kMEQEY//OB/FUBinsoWNnb
PNXUdGpWkjVI1BVKUUiU/0Og+VlGt5IHs7A01e4N/nlhryKYPuxK7iVWgJyTLHq5JI83PcILm6lT
tofujD2nvNG/N7UyUtk7hwERG4/45W/CVZdYrA52+1JJxbfVkkt8rq7MeolLjuD5q80jYzeauOmz
G4yCahBsSCqiXYjnHNP/CMP1fMl/S/mZwMgR/y9zYJPcL8D7mEyXJMVUHCcZV/rzrD+7envO9w53
wYaB+lWoRVfi9h+v2sLu7WMtMDDu4rozxuMlQvyM6LraVxNoXdzY3YUP+zJyvoZ97X1AZafpa0dS
fthwtwClVL+ANR7hkdoNir2l8g9/WFCVn2CkCH9H1EXdI2Uvz/wri4L/XtPo1a92eo1tmMsDhBjV
1GeKAPDS0DJXxuKhIs5LHjls/8xaJZtpdcIx5HeOwYWWH4QXFMKd4sZiC9nIyi+3jx7tf1MbRWQr
WZMFhLkAvEy68ZNrvB3Yme5S+wie40hPAqGGlgagmznQlO6UNKFC4fNn4agAYw9R5TFThHB2z60y
r0xB73e/DiIUOtwfyETPdovHJb0honxApgX0ipeMJta0zi2Xs/JQVwW7j+3B2njKGIIPC1SkUzjc
V/+udUoUQBDm3Z58Iw/eLrl0nqSdpGjfeqCacZZ3qncYw+tW+E81ze8OVVgPFzoZSBAW3+9vszo0
3HwFNyKMD7SeGhLVnITD9LZEWISzWZkJ56iZgR6kVC7ACkzOxU3P9lNhMPUYTurwt/NNGWkLW9EV
ZbFAeDREVl8lPaI/+KPwvts3SNBge1Giginvk1mASY/tp4EoFmBDTyAzI+foeg8LkL3uUQBDin/Q
jesTBhMeSg/0qVzjy4+s4YmEhyYn/123mlm+D8AQwgfylMgTLAl3zrH/OPMMttYGXRFZznp516u0
5BulYO27UEfChrEpJkXI5jg+phnL5cgtQzcSKJ4Dk1qJPoq0a0kC64mJ/6BcfolabSDdz3FPuOne
4QX+yKD798/GZeqRHKx9htvWkzjEOEz+2shSy2dos/1zMP/bdJSdnY9DAYzm3oR1gr0jaePvOGUm
+mrhNWDve1nebgztRd4xMaEPNolakPcr0NUR/eVZHCZMT0A9dRFQP6b4PVxIeoJpVUf3s+ewJFRl
g27lG3DOKed6kvwH54+2YiXb6g2qYql4ouD46an263qJPUtQMYRyJlrC8bkbi2Eq+6MzJ3PdX/Zp
MXSXKWGD2bctWyZhPy2IUyvVPrFlGbg8RMMrkROk9qxLHF+hVrRz+mR1pxKK9KR36cGz/HHBE1LP
3C9otCgcS2/YFkA81MJ/5h9Eqweh23Oq4tnHrX7Ul1CLVOGdE8t76tz3nz2sTxysD5EcI76NH0va
rlkDYHFVYj/hQ3nEwnggNtpxHpXNMZsaZPHehyc9O0G+6mR/pll7kJL5F42phu73F86yr6I6YEWg
6Xp+Y/bUtIWqZ8HomglexVogungGlyc89ko0x2rAIZ3umSYE56Xx8oJYk3TEa365QbnKmb75OM76
Ys/vE4Y+PowRPGxFIqc+w4I23krmDCLyvoiwMxTHHDG09cyVSLYqWLJJ1EXr878T83UbEnaobsNv
zLZPFtTGbJWTT0Rw1RZgFvkw/EUcGd7LbNWyNc70so69NrKiqC3dUfOjM7mM40dAac7MbW+mnOqi
ClAhOmU8R4Pu12AFKgIBvC3sKlkGJIKayk7+NUJTeV/I7mELq9Q0ATPmpecMUhqCFwwDfFm6MwHv
vtIPfGmXcLJez8MUzHMPsPtS/16lBVN7MQMqmLA0dB9TB/IczztGh4DTuDa9y285bFzn2d2q7Uh6
oqQxsI2VXS6eZD+2kX+PY5XTNQdqAcL5doDKvpXdF2s751KA65eax52DD2/NAwO5HRA+8HbQXmdK
eGPXQdoYaZhAj5WS7cyETaf8R+C5ZXkLBr/4V1TPStC6LHJ7RQuA7M1kxF8vDug2AvM6pkh0URJb
JIk3olF9tpeA+UE2gcwnnaYbUiZ7V/T9PqxN8pwrJWzdogFJpsz17qaIE6uACyBszed1s0pqTYlC
Own3kRmPTnTV6LLuSZWPm4HpL791KEX97fyYdwTbVsqfjcrz7giIBHrywYAwKS4wIyWHslU5sSw2
zMo3l+F8zkhBi8bkBBBNIO0epsj++J1VlmNNAawMTpelrU0anvJB/8F15Gk6W1kyiiTRlkeHepea
m44Mo4bm6ds6/I2BXTOdocl+7b47NdA8yb4IHWznWx7RrgseCTqZ6GSGDMN/VPN4JTt4ygewehd8
v1HL9JmGBpJOEBNIg8h7wklJxijvFLknJVr6M4TbxWkn7mO7+bX4UTXEJf27dm8rNLGpWLljN27y
82ON3OlHk6Rd01sRpPLV3GqeRDV3o448S4rRwzjEuUhsfHp7cp12jAkhqsOf++EfXv0BN/ZGcL5r
7PqucUZqBjLZ5h7c+t9u5pBxA1j2oXzIJOABO4wDg1N+iGC/HH7j3BqFS2QZC7n8DJMIzLaMciJi
NM8KklSKBp5rD/Aqp8w4TtEAyS628CBIFA7J1zdRkuzEwvtwh/JH808pOBYXhHedHRiGJ8JaJhFz
exKEI+LkO3Ruh4Rh0f+gIrMJt/A6HGpzE2MyJ9vBFAcT/EcgLqln9e1ArPZ8KLvWd+F4YghN8K6q
qqGBbltKaWBPbgzzYFAdHTH8Sd180cnichAMWp4x6rpvvw1gRGlBNfBq4aBjfBmx9FY9MYFRk/b4
cZrc2+LlsGFG1JsKVPkiv4IMLmKnm8CXcpFYjdDOgJAAXUHIfHKioIM4hFQ1rVPjEEulkJtLzZSy
9yGGHJjonysEdpH/HPLY7R3ZBMwe42BSonjok7TmChMwLFYbZbGJXWJd5Oedu/z7TpJFDj/fAVlH
P9F9ruI+NyIEWbEDH/zn7i5r0YvuulsCIpIjG2qZV2Q5cei46RJdcjRzEde81gTTkM+l1XtV0PRj
t6Tc6N0KmD5718qYi2w/pxhpVBfMePhQH8XM+r8T02eIK4SvDztA1AAr+CXtHx3127aYJCe3UrFK
nW+eL9QDwFXBiNYxyvQG4BFYgxhwCNDcFbr94diGvuzCJPWwGbz8QTOo7iZAAbGcdtmHW2TbJf2k
AJWy53thIUmn5KqLBybGWZ6v3cSc7AyqQOMRWfNCtcBHydxn7KawHTfygIPO5Kz65aDITzmSifhU
+S1/WU6tZ2iJTh+wokMX0Oj4Pua0fhuCrwZCswSgUVpvqzEszvkS+25AcEgMPMObOgxyekQSdd5U
jZNSsuFnP6J4o37RzLAExT/E6MukoumFOJ6HGVqSEtROP5QYnMfyMzuvPkX40Za79HuarvjZNrAa
VsbSU1HQMa6bFsqXglmXUHRK/LUFMLsiKEZnCYtQMyYoDWW4ddFxNHrgguyhlCrmZgsk9X0kpoZE
QWeGmORW3gVfL+ekbpAIPp8Xvvx/EPuSeiQlYwOceaFRa+e4FbfdRxh7tlSrWleNx1JE4t7U1C9P
SBf2mo1opsCYI0dD8nPNKB8QRUQLBGPRolQP15i80d+kSpB9iSFTH+RjX3S6tA5VIwtnrnI/Gfmn
HeEqENGvZUpWnXRtOrGHZnpdDHDA3JUZa05Lcn8Q/sNXczORwbGpm3zeXEA8xBBDesIB/8IcwbdU
19VrP3ZDQL8QTnixW96IY5RyexuQBj1UrLsIZicUGqk8MJm+IneFgVGZuFW0vCsvGMAW0Cv9E9fi
EDv14da+kiMjVxPCBTsmaGTbjuqULLrFNs9+mS8nzVSjRs7rNOPge+IxBY3Zq4wOny2FNSdZeSci
P7UnBDCuQXN4CdWwKSiZ+L4SkcdV/8Z4CQpLggsADk8vBP2m01GYN4T4tBhoHda9R/JG8kYF3DxN
/XuecqofOokmywxVL6FHkQhOJcN5AuMKywf5fCzYPrff3672dpwMJLB6dLSGp38D2DoqwkzIGXrE
23NMU55dJrjT6OBrJlejiIC1NAdxjdXIqrnarc++i3LFMQyNFy0aTT48X+Rov2XTdpwjvQZB0aax
qs0asQ2N7hH8kZjelVxbTLtE0z6lb7YadUZes46chE5o+X1wwzxKNL6GDI3syVAlfVL1b4YmM7nr
aqAha0MCKLpbzoHqO6nt51nmF2FfyvrS59uxN8a3tYOcWRfI0NM5+AoqsJBWDnusFUBsxk7Z+F0T
nDBhxRKnftbbHph+07h1/8abn1IxH5/Ki37JMipb4i6WPNUFPNuJQNLKy6vb1+x3p/Ms+oy0PsVL
xOqtoyk7iivyensfsQKvKT0XMK2H/x1trGXHzAXjMHAIsTw76D+Nqm+WQi+TUp0waM8Tb4N5Fm3P
v+PUmmToYAiwkNKTO3VuNxmgi7hLkF5CwEMDogStJS1rFuPP5xOj8W5mYzcNVXXPXo3Q1rrsHbTW
j24BZo6X5QxPBSo1IjbFrXn4V8oUqHpJ5uWpyIjXCmlSgFeytFlgT4M16fHu0STbV7dOEf0r9FP1
dSSY6CbbYOrCgcmHGd/IGQTmfMG031sWQh86PTnceKTdb1IpFAtS3rMLGfmEEOcpCHCYmODb2Wn4
q+Qwe4y1QdRg3NPV7Yy/ZRpTbCiQ1MwIpTb03mwYqJ7micVGobe2XXpqkGZHERqN2RTicJKkRiSx
UgjT8MUXfH2TZlfj2rRMKcYpgcFH4i9JUwZxFUtZeBiup5aUDerfus36Nf5zj8hAVwiVl59Xl/BC
nL3vH/rPYyu2wQ5Jeepp05r3i2h1wuRXfym4KQPTi6wNzCiWsOjbez1F/cjb8MglR9oOqcDwsWef
MvSjaSyJv2EmTl3PFlx284w791XJjPpEhYjdanJ3iTzjn+QWu7VAhLxSeGFGZUCOg4BuPmHNiNDZ
xVYvpiefLcDYyg/gWiUWb9H5/FB3vmLGplt+w4AEoRiE8PYdv74bqq90RD0hpk2ZddEcmstTBj7B
EvWAC0bh7XPeYnKzTyt+n9p4EBvFQ1GYGtmdXSt5LnqNrtQo2pm0z0MX8G47tHAnZ+kjixEKHuAG
rPdgnsrebQkV9On/PizGQf4L167nMRAEfW5wnO9q11L3WTMq+0f442HKRU+bEvq64ewjMgZBQ26r
jiF1/RhlH7PKsG7wBPueHkLCgh6h9TQWPJV0Tnna4a+3riUPJz+JyMMusEH3y9F4ZtfTIPWBeUNw
aVV9+1oHiYkqMgm4/rDbz8RIMiJF/pRx0x6SL7leNu6nQunP59C6S/ehZIiUL6LcEGJqt1fwI6NJ
x9BqdXQxK7ZyesPOWv6YX/CLsYnQ5vHUvJt1NsUUDGhiDB30IG8mSpwp2HenBHg7hAYvDLNHk4Ni
OXXRpUeA7iELP4lFVTz9yMtoV2KUKUBRsjVwr6Wj4bCCYHFGTCpBUOfoGjHhwCVe5hLyd9cjFYO1
iUWyVxe3m2YSc6jIfx3BFSCxjzH+B3QPq/S6t4QUVKG+7cRKMC1pvbPig4TmNO/LQM6eDMEhtcSX
t9jXwMiGGfgqfolTbqMpyB1i4D65NOkt7J7Yf4ojaShV0jrwUDGiPqQVYrssYJ7AFfhh0idjDwnA
Lii103IRDoc4pX1ormWnGFzxFol1/ZHnAOtJlukoRzjAs+DX1fLr3LUCgX8nzyIY3LFFJPoONqp0
uvGtgMQGKk1R1qm07K3eFR1U1+QKdZ3gyu31SvF049l+V1J7JKcSAePyC/G3u8mJlZIW7Ow67w/l
VVJLBV/TVaEeSHoM+Z1QupjYCsM3n+b4sNIptQ6ZG0MX+YcygY2WSgGHyHBufblofnGc4ECSYHoP
XQr2UUxeQL8ra+5OxfsK9oPat4YKHBHLQBBnomssx5EdinsMFioFfvHA440MM0IGydTAdhuIXJmy
BqkAgzdkcQJclIqsQFTxT0fraWUKep028EuxNKV/h7SH9fdwIQICm8GmEcB3xy+vYK5NyBVAzPER
CoYb0VGGsS52qVsF72Jx4gDs9BMrntR0fa68tZkxyk5tZNrQJ+x3ddnr9m0gEA4Ci0xqvTdqMk6w
IbxkstmmcpTqTWWwYMLY3oGGK69VlJQh+z86iirQoZISuw7mLXSr/6Amk9LzeSfYblyeX6uvWzSn
wbZeVGvzQGDx+LgpY81Zhjw5HbATApQvYxsjbE/ie4w3cAflnMW8ltrlg2j006oMePB+40NEdSj0
tUdgMEZUpZ+z1SFNpzcb2irKED0dKiOastdjAF+LLtMF6ZXUH0z6YeqBjaE8X52ijNY5bkyqj51q
ctrowtZcgGzz3jk7866OKwAQJROy9UIvQjO2BBbvV5P2mgTLheHKfccBNIXdRMIv5HCTYBAt/yeI
Xcps2Uzir3iRyElcGZEFxuwhW8LjW02ptG9cUXD83pQAfAyFy+il4nohUqI2MM52P8RMnlZbgwwY
34pOr0tdeuLwW6viZfS5tRONMC6SJeUznu0zFa8WN/LtxJlWCI3wuDVK7BSWG+h+qsOzjff8ladV
8YmjnNhOmHv6yiYA6BpVUPXJZo4BaK0R2Tk4P+OGDBBw9c/ZHtawXRtSYXgeu/HxK0GLbzkFm2zR
GgWSEwQUEQDqUuPgfkQZTB1kAbIouKUTMyJ0AklYMvVFmmDS2R/XKROq+sqogfkC51JMdUtun8az
uljXOrDSiE147BuN6KhQ05cqo0bH1DQmJ8CLdlGjbWENDrGdMj894rN7GGPyXFeN/Jfz1C1q5wJA
ZWMz9ViHn959lKcFUt+FGAzlqFVULg3YiXx1NEnb5XWLPzNZfwechK89hPm7A1Smwyxfjob5Ho8W
i9Kh8tkbClTKHJruAhLyZzDkRSnpLAX2BI+NB1KE3P20yGduoJYqj1gs9aK7MxtSiA2mo+V92dij
HBLKY5HV7Q5IJPlTPVprvcS0sh3MxVREHLL6vVNnP4VdWg7CX1Sf+hFSbVlRla8NLUeuaCCrHJ1Z
t7iXiy+pSa15HJ12JTy7u+/IPJyO7vbE890zlZDqTflLo4gdVcsv8g2lpxbp2Dj0nwsXCKLYS1MP
4tPSDuAb1V8PHr6fYVLpBCNuAzk14NIRY3R68aK6LDbphUWpVFN/zmHO8YFRp6gGD6gr6iJzqGlh
Xl9/h6Gui8a8xX/HMlez7MDI2jP2EAyIeWHwocxbxBXZh/Q/zJkojvAetPebb3f/yE5ew337zKGX
/kSwN9Ew0JBUxin7opayzExVjAYcFPPCcz58+oTObxQzRKWdzVU//514ZggCjLSAiycjsFb+kfCf
7KaO5Vr6BE/y7aiANUZCkm5rwUUc0yp55c3H6NhTtlUDsjWjeveNL+0NjW66H50lkaRFqNDZBdlm
8IDB+y07TdCX5lPq+PcfsnoEut4wbwA8aygRknMA88QA7diH2YSeJUF+8921X4b96WB3sHso2wHn
KNlFQ+nsRS68hSfDFuumO9D2ApB9tFdF5phrv/V5LpXOoR6cn1YZ6CVjhD+AFwTjCTEEt1J3HsY/
nL7ZfAH8uHLXrdqRBshLWxoxn6VsCFjViLrOUt8Wic8Ic6TmBayqtk537qMalLHLL/dTAVc27VhO
n+1dBxnfEWEaY0U4dNGXMcowLUCTEjxK30Rjzbeibf2hWOzblFykBz4RSViL3P3T6FIgCkmWaLqc
bXos9SyYZFWHwbuvo4gxcmPxKuGxP3RBe/HzJOJn9XcCOib81FRsy+cxFFfcHIYAYAVgjJra3hYF
82pQpNVJUudu848ugpRFsAZ+/zkQP5MFWmqKV2B4+aiKAO2tBHrveLbaufudxCaY2ZsyGl6voScz
285J2BTN9FT2L2uRP+03P0u56cbHdDtQfH+emzCWj8ywirtPYIue6pzmQKnV32A27qT8pLlQxpTT
2VfpvTonZOH1S4kT/kqA5SElRVc8czMhVHiUF2G7wShNUlXwfL+0tQ4mBjFeejQ4Rcp8KrqLbx8j
5TPVbF09rCQcRSBXVuh7TGKt+3DbL3Sw/CXMla+BorRQAQbUUqJzF+oXvsmF3t6fbYhf5ANEvcaa
yHECfbgCkIYU7VlX9mw58zwzSi6sKbDxLktbvdb7XJSl60pmIyzBqXB8DJL/ZQEI7dhDu2x6KGpw
Rk1wvDVokSfVcWucclb9IL6Y8DC9UgMVtz44xH1TAJJJV+Ibd6MPULCd4KzC0IyVZIA1nDt5l6JA
9umC4ac3lX0okXJbX1zX5KnDokl/92obdARVDzZ+dv+Si0nI7h4fHDmX2CTPiYRW8qhAiss4D3bQ
a+Uas8c5twmOyapvBstEY7niMwFA2bzfHV38DZLyMb7zLx/nZlAVnLmSahYu0Hhs0l+hXaZD7O3w
Y+XQdtOs1u96pyvbW2ssRf3BRsiEAp+adfQfhTfIsU78giz0TFJnhjredU8mjm/Id3CmsDdglh4z
VShrpJ3hiG/MbDJbMzPevpW6CSWwusbVnNb8xyrkHk8eP7dBvNLXFVDw9KcrM1Xx6CJHyyGBiru7
kdBbXfECzGIXNDqRvEQoysWv1KZ9QlCAkmS1wN+8Xamfx+Mn55j0gfH1NahyKtEHeNnQ+8X95z0Q
gShZAKGfa17SYG83GfvDtvJ7gTSz+2zOEfTRO8fYJr53GGpsXKCC5x1/Urg149JKKKNfbW56z2bw
ttTrUyxn81uzX2MGxPjr5j1Gs/lGGFRDYUOwc7z0cLwJw3HsCPBM2dTEBmviex4vVpPyvR3nLnqY
ahYgXL0yuSbLuQLYCrnlcigeigDEAYi4Gs2N05XkpcXFsPt8ykQBXLxUyzgYaEmgAiMaEWX7U0xN
cixT3s0TyR+nujbbig+0WoxQqtDxxWtCRU8z707IaJkjOYMuYncgSafCRwQ561EdqdaoN7sXqPZR
AaClLMlAQwH3PdVj+7nkqdAJEp6Spd5mP/pY4i2NExEn5iFIHMqlpGSw9GXzFZGmmsYPD18h8Z4Z
VASYcoe7K6JHu/tt53J02Bdzk448t/mWFKy5rCob5zL195B+aBSaoiEP4L800JOS1QTm7Ice43XQ
XXGuWeRv7zb0+5UyPAeZSNupeAyQbNQlbbbMlsOUD59071TkxYW/PvLXMcTMTrebNBNfIgRX6oZI
lWJqMDHVT+5D9Lw8GBBOJzwoT+hn8qu09NaLyd3Q7d9mh2CwknYT1ZsOHTCq1JZ0x7m1FfdM/4du
gLAVJItg5wi7lLFgVkqncDJntbzMNdxWPygomI+b3CTXVs4waNi2F66loTl6rwJgeBC4u04Vk35V
eAqz3xEfFrYPY2LosPTnutimWuNlAt588RKbgcjUbOyEq8jMO/LmyTSL5Uqn4eCohF/b6L0o/o3Z
84gKn/dXaV05+MNlcQB+OgLfqkXRF3giMuS4CxY5c4tXf/rxdBr/5xZ+ajzO3ST+gwFUw1AyZXrV
c9ttPYe+X+zkwGZyAaQz666z1nU1xc3d/wf3ARPswqSIMcICwHiF7qmDc1oSbx2ptQ0Z9BPbVYeX
wapk7YhIcThXDl3PHEBDt1Bb1GMTxxWeBESU8lwBi9yNOeyKBI2jxxgrxmmM9/95bQvChbrPgXAK
ECVxSi/8epdk2tHv135AJ7ob1ZsxDIHJvxg4NQQVM8Yq738ALz+qBk3RcUw3YDAR8NPmXQus6Nbf
9hlsgRn3j15P+cyykGsJlj6/9NBP9U58sIFaG6n6HcX0mWz19bjdIagpmIbBDMxdUQgvaUN+w8CK
AAHOsg884fBLNZESJcUkwKFb0mf6rKYDzVB6DJRyJN4DtzU4ZARUUTvzcIUUGI8838pEwVpkHWO4
wlO97a/vk4w6Tn5kj9BTvNjGg0C2Su2aJ6NcUG6Grehgk4UR15HaAKdJWWRMhSHynzjK14HDdCly
spzfktQjWRaW/M5sHiYVOKyZC8pj15f0+4Jzh6GIqCRtUp52P7YyiSBIlghbRMPovO0DjXVJgiQe
zbpw56ShVlYkhunP0N/BE2J6bDjPKdm7vUI+t8X43vB08iaF4BjzAduhwSFjBx5rwChRD4hggYkY
t3ECNjzZRYYvtRDF1d3hiLqt9vGTUh1GZYxUOmEVkjQjYVgCJWHhjvheDHngZi8MTQWCZa2CbtwV
5MbA2v82FZgiOdF6cblwrl9th/RLB0gpeaG2om9SvyNoCJz8q5GPwx8nfuszLfN8smertRz4lZJw
4vmSTNWica8t/xOF6LT3ItBOIjmDxMYFsclWPVSxNzZTbACxYjFui8JfupwEQFw2t1QFyc6rp4z8
7JfDoFrxMLjSkWZLvTfxnqFWnHBV+M3rvq9ukXywL9e/xbOAzcmxJpQBCOowIH9Z6x0b8CSqLFrx
11FIl5TMQ+wiUwQuC3c5GmuAHIwQLs4cC16cqBqxYWpcL/mgIDjx6WRHwQHYR27u8rYgMHraT/Rf
8hPR2FmZvo3AAIkR/Q8WSPIAJjPtaCsVKpgnRVSSk8cp96qOppYQqj4bVoVdtBcP+p3rfWowBL8k
e8/JoNwfZAzx1iWh8HFBs51Qn+le8tawYnu5WZ0vlsvqL+DMOMliz4eaLLNUTjla8308LHFntVg1
KrF/Qq32sN4fLTF32tMEHi99m9vDc64DUPHeT1dOY3M+qx6lnNlFYu/FSH+qD/hbh0lmjv0wuh//
3ipvT5HqJ6hx3eX7HyhKXuMn3on5jydEBrDXY3yJqWI1BJJj/J5XwoMyzYI0nJYaftN7h7b2I8xV
NKXR27JhWRMNKipeuuHr26FOvfPwTApvCC0LuXECUew9XEojTM/qqKC2PFxtYnJh7EEHrJs7t7a7
OdQToi1RZXECeDkV9jvPpIQdYIZAMR95U8wkza5iIPzYqkjt91UmFhkodyn1zVRdUDGhvsCJFfPm
AkbwFgK2hAcL1S3QKjlUufTtkqU+K0FzmZmQLfNMSFslp74qoAoy33ALycM+8tEzA/pz5WVHd57T
M7bysRGz79ods5AlNBmAam2fHm9A0U1XL7tLvG631WM63S9qo8r/o0YsyZa7mu0f3uHDFW8lqIiT
MdOOcHQ88xbtnvnef9Jw6oRvbKWqCbhFp2xlnl35nPR3CD0Wiwdn77wvUWF8aF/NtfPpba07dLiq
pDTRdVR5Ed9+Asbo2bteLIG3CUrKLH8ltXiG/01Y7W5EAs2FVYDOL1rhi1rXYuHmG+59LMnj2P6w
vV+1yG4HcC4DtLX3vSTJl8ae43WZIR/lz1PNiJCUncUtActBr1dDB8R10GXamFUgirlVMh5m0Hzi
J+1I3SlueCaAmURhtBCH4SKqrSLEs/8YRuQn8YNb+2r91yj2gttwNXtXYsaL/dYuD8xUJ802B+yg
3wgEkGCqVn5d12ma0WFzpUDiFta3cHSC+kS6TOdNBC1ScwNsfk16bO43dvw630/PW+i8fe1pSMuJ
fpHteFl/xyGE+QbKEqJN9sq03KjQlhQRQkhDqm4ipdBm4zyvcp/A0IcMOzHvCH/AIBw9k6a2TNHJ
hstDXG4PSUmXyBN/fKbqDGHTM8dimLO2bwDUtFxFf+wy9ATY/Gys7REFR3M4DikZZg4zAZyScVwm
ILDgSlDZ0WcjMaG2gAme83KGCbYl4k+EUhRCnas8dmLS3TEut/SL+fd0CL86wBu7kQC4y6LRvxrb
lX1gl8NmpQhowc4we6gyhFUEIujsoeipYeEEQXnlxUiFnS+VBY2bBvgTeUp18d4k2FIRLylcWZRv
dJP/tnGG6DEmP6tAjz5M0IyZHcCnXwAj0vQDyatjMvpb5IrwQxG+YUVSny7BskVBgCTg59kyTpVK
PkKnoHtWsMDskibC4z8cOeDC4izWRg0N9iC1m86oubTM8UTxOD03w+PuuJokbWBmqgNUwV25auK0
bCWfT3BJXup3Nv3c/8sCH+xZwhbRo7WYNNeAvQgbF/J+sYcJSNbMwzfR0OTMLlJym4jOWN7EAeZP
nMGFGZtL2TXNz55CP6KFv5jpmI64PngegZqkmW6x/VAPQTKMHNkENbMBh0soDDH7urV15Kw1JmJc
CbbeYYkYiKSQOXyk4MCu9eAOmazuMHJ9naR15JNvOvPIuY2tn2051J5i6f0iDPbDpXkGStz+BFNY
ZJpChQCSNE6cpUuE7J7lZUnGHF2tbo+zU2Na1fJQM/JdBg+LX+E/A6VO4BMTYvEexrhhSMkR8f8G
2wIeEbVjXJntpvNi3U64wxoDR4Erm47Fs2Mnvjdrz8LyoHnPKhdkacYItnLPTqQKuWrV1xaqr7M1
ZoTucfhLlorRZTUvi3yvgOrFe7zMxvL+g7IiaF3uXsLxFS7Mn00TT225bEQHDhR0kIUKBIcFwkra
ixGXEz2WDiaAdWfOLnH3ouG9GHdApqR1dpWTP6NjvZqhhhSAhuKxgUSRXHmNQvW53Qy3CpLUZTMZ
HmnPZar0nkQDK+w/3WBH652N+ocrKaSG1xjU40MSLemaG+II/8dgx94NlwI7puggxfaw1iyUp/ui
pc498RSEy5yuOfi7+RC3TZmfDosQISRfA7KAXXnmh/cnthFafZXa/MLGajvhqb92pMiStVav7nv7
EZqMU5i64+44h6CxindizA4hHa6RQTr3CkP62Wnam9nbaWvUo/SZvvkKUjS7+T1EC0G8ltPcc8zO
OAN4VAV65xFUccJLTGItg3aRFkJpDfqANOnsurgAebAJmRHuUNr4Te+nfNKlUd26zjdi7U8/lWjs
XtEfS7DpYUTK7/AXOB6hYElvSfyabeI9f+UPqlrQRwKcsRxiuNfLgj5hfPL7Gw5B+L5AKL2YTKnq
9nBYiFSaVkVPj7KRyLsDeLvE8GiQY5ZMea2EKHnK37UDLhaff0N5cVTuVz35bS2LozQlQRuVNMeY
l7arxU+RbhnYLBx91Jk6MuWHFcU6KhgBvO3Ho4+YJIAKDhwIVwNhtBv8yvnIBxgWD3NBhaTCmzBL
Y8s1h5MMEl3fBLljlHuJ0HvumPWeA/i2dmkn9XJcAGpTn3LrVdne+i4tunuwl3kpKKWK5nlU3XdN
XcOIL+Fmx7HPLIzio1gOHMMeZECfjie4jIYAe/OlL9hpqieDFiRnn73HI9wbM5knQmGTGGUW4+y7
HyxAYicECY4nHZB+XulUXJo1y3ygV8Dqk7WzSVCHLvL3fbCA45LZBWBlds3BTfPQc+Sc7tfVrOKi
nrl8LVOVEUqswkBPrd61wRWNEGAKfUwslMs0GRgrnsp3SAVla1EV+cLcu9DolXs7LpU/GygsDqV9
85LgBZEUcW8SPFgmjgfdhSMSb0tPnMXt/cSnytk3QwdP6vX0Lg8fgX1ShsQJX+d032qPiGAvOykQ
W+KyROYiNO+bs1loN+1E33oxAsJ2rn0BQX46AFd0n44aw5FIrUnUPcvHUYYZMqqhdEHOTH4BpFwO
10538ItR/ktvB/wxd/Dc/3JQOaFCwoPLTQ5RBUBZ2uiA9PXvZ9ebL5vY9w/u7t1XyGb27YxW7d6A
1owljPU+hceRIrLrGkTVnfbblwmnQHxVOGuKechJlis1nMegMnOUGOa3PC5IRADzOANBDQiKqGJD
rTI8o9sd4QwxUpKQRleV/nV2brmALlWY6Sh5KJv45JjYJ96gPZUrGAzMNbcPsTXDpPizYkssZN5m
qDbUEhecxPXPAp9MXtftJw9EN8yjdb742yB6BjIFV+SPzryrIyVquiCbFqbZL4fZGdpNELTqCJMy
zIixf6NL+9AE16nMprlnG2+2XABtXTN5UPS85yoG801HGZbqCVULsgHt8YMzuAG74QBaus0NzV92
rXp8PUJk9QUsjk3V8mwxBDSQlGeIjaLjzyY9DqH4iE9gdBHklcZprc/r7ANQPO4ty/lDbBhUDhBr
z69y5+J155MCoc0huAyLRfkH4pvHXSpxf48SSFRH2GMwQkEupliESL12N+zlzNjwI31LuMBJS23c
Z+pMCPa6z17+dgf0YWavAeZ7ythklwCKFB/u6oujk5LiEOr+vbYlGLos8OnZ5OZ6BKl/IIr8QT1r
+zVaIIZ0aZnQqdBE3MhviaTmVlI6KQda/an/ar3laGawCvsylWEG1UNWB95A84PGWQPvIij+roBB
9qfRL0qgQ+Oo/t24FGmaDIAtUgchDS9rRyjS0hzL7WJurxCUVSd0zcbwniLOazX1QGBblHJqsBpa
COHJEbk+fEoL2Bav/4uzdL8Whu9d0MUCtpSJVwJhcmWvmVc5CstTz8pXFykV9RCKLopXOWKNPM47
XY3w+fsiYDBHbOEkThHHJOtLDjxWA/org0YdkqSWKryYlEC80XOdQA6eCEGD3zPF7TDQIlor3muw
dPVUwkIY7FIy1oS4oouzRNgBBeWWDZvszwXb1Y5PetAztKhuecGtFGqXKASeQ5/uiA/7wFXzY2/z
9pMI0sGj/nxg/n3cTC0clB2Kju5ItUaOuXdEUHD2MHsh2OhAWKMKyQuYpUAFHZ8Hn4HW14yj+Khu
RaEHU5Rjeh1ZmHOarLR/vm4utyWFwJ3ueSYw+dmlMdqm6xpwqpaBBvFAjVczZf4xtxFj4Fu5KY5A
GUmXKR7HOy++0ajc+vBX/RJRwKhl6zXKhPK/6lWX+X1AbLjldjwQeIsy8KaVES/Z3J89ANgsbOsp
PuQaHeFvtxB93krTq8KndzXu4DDh5Oo1pXJsmeDtV59TdIkfygnTNq8A4tfnAHarZUPBPgifM1ma
jZr0RV8XBrr+s144cDSU6aBof2YJhbWXX2tGqezO/Ib9+TkkpOFAmeZRrrs+qaD6GlPaVBwVjpQO
LJDARO/RjhZpu91Uu+nhNkFQZCS+Wraw7NOUiJ5UQVMJjXah4Tcj3nPMKenpc1f1xnEKBfCQWKC+
e7uieNnE1zahNpPbDEOLyFmKtm65ykHlpNfbJvdAFC0UcT42I66QwPQOSlVJnqacwP4VMvXFkQ7C
0ATUDxdkQCYIv1z2yggYeYU/v7RKa3ww22KPc/zcaskkJtGDJQKZCswL/JdpjTlDijQHD31ugcUi
9/LBLX+aaLJwluhFhfzJPt4f0nYeOc13za6eUN78E2SdSZn1FyeZQhM2wGIEnEfSy1yvrCLBJSD0
6UJmu+qC9BLDGCv2T2wzBuaEhMz2mynaJfUtsskqXjS+Icts6c/52tXRpUEoNcqUQ2cw6YDSfZSs
bqxWH70NZIOBycurznajBPI5F98k2vZWRqPnV1DCMXoVRm/Tz6oQNE5GUhb/5zr0boGBvjKA4BWf
d+hGyOFVtkjrrxgqqMZlvS73LbSmgw0n8wg4Bp6c88fFrTElFlLpKTHYPdYHkmobK/OU2lZ9J+f3
5asULr4h7pB5GSVE4lzVBtfvBaFxJnOZdtbqZJlXrZ6Yu3grC5CH8QX/LqopZZCUmunNCl6YM5WI
n3lwgeZDR/eorK8tyEb2kUplJlKXh05q1doLusm2j2HnE2SRDrQRfHF2rD7OLriuTBwmnWiqll0U
rsa7e7S3HsOcIoaSBS5LxJR/36vqZRICMXuEO+bYe9DV5iiCh42E6g1M1kJ6T+G25mcsvICwhvZK
W5DnH4I60FLCpE60kUgBMthOUkHPRXsn/llpXvX2Cw+IMmLtiKlAI1M1CRvCdlseqFCbhz0EWrP6
x1IFqQLz+iS8sBZglXcyBDZDVdhgI/55fReO51bJG5guDjugHDcDgMe0IZvl5HndsmPxJXEUKYMQ
rGwF2VC6IlhRmN9DoDrHfh9xGmmdelKY4tnELkymBgtvDtwyPysxHO5r1oxvp4T216hhzOgQdKr5
g+tKbKwrX0/5zbXjJ8w/U2AoQw2w+ERtQXODW2PsCRF7HGCTVkB9IgaqerNe4GrBIXnbaxXGpbHW
i1WNf81WXH2yscD0tM9W3j6hMfyH64Kk85ze96nTv/QbQ5Kb5pRIzmi54SYXoNLQIYwR7LOh3iiK
bfuMcwzXyP4m4mCHj94wfcGt5NCImxuQYk73TacqHLALt+moSO/mPiEnugxkaZMIBJxLp8tzEOs9
G+Vitr79QJ8F0mtuUq9J6/ElR9NN7eAAu6GIh63tD2hQSNejvqdQFji7bGliHfGOioIS9wKJLl3B
c6VuE78eutIcWExSXjsTPZMVDtQ19enfPTGLZ/d9hN+zU9dd/HL1NZ1XEXsPZCyKNPcm+X6BNmOi
kd4QQ8RcZpLg4jfc8BzxG8PMBF7OMlzmTS1jIJbseVtTrUG0qK5f4WemjdwYKOUZUoIsBHVnjUDD
gbrj6yDZxWz3JXR6tGpKc20Tho91EDfQZDgTZJIvrLQ/0A94mqz/62LfHC6KPKc8wIRKdLlvo3VS
2VlC7h7uYbSMxR+r6oERi6PfvYf4zObtyTFbv47S562SAganMpEo3xSmQzLRpRNZY8jTGCrD/iBJ
CNzddVE6b6Ky5nieFKQQ9Du+h9b4PPpz1vGLryl0kk2uqGTlhaJro3zYYgFjt93Oxx1NSzaR1Xw+
g8R7AFUSxHNVEl1suU6YYm/kCtsElJpJaQ2piJOBQnT7I1CSBRAdVYJfbVI8iX6So41GwN6v1Dbw
+mJ5BUNK41jewTKejAgnvODN8PBwa3H6H7EEAllNznsYiCCfaKcljr9/UnFbfOLP0DgN5mJzSL9z
IDkhu0fuPoUErms1a15M3b1KhvT6LN7rUdq6uOJwrHrLoEVJP/QEs6KIPzJe+86F0m+KLxlJhgsA
1CG0HoIa19O09f9jcSIHAF3SDGgMolNt97ljidehifYn/MfLVv9qlh0fu1c/ZP6Xtb4ak7bAqNFM
tHoNImEYllUpxAk3nx2OY5caEzEVRqZv6Ku9fF0QIbR9BRvAzN1r7x40SN1P8U720bQII1aVNSzp
F3fck/oyEEZ3GH74TCYCbUD2Cs0WE7JuWIARyJARP7vfgEr/A5y3VvQk6pSfjiaNjQxE4earnWBq
hU8gf75prUCI0LovmZ3O81Zl59ynsSMGtFyF0WRZ7R4msqajZ+Jp+nhGbEdcpEvPuzoHW5+Ceoka
5p7tjivv8xKkFhjrvvfGvj7UMiKow/veJvFMwjdNUBqf7hj4r1T5Goz6liFNKOw6wAKfKX9CK/gy
o5iiFnKPM5kP3a51o745ucI2S4tEMpSIWX9Mk3Roqf+9lXiinV+tGCn0hBiPWaoHlcx2tkQ7mTOK
wqQkFXcejKNUTOFU3FjDi5wrPqX430ZJ+uUx7UdUnnWwYrkmdnKNkf98v178WuEx+4ikqZhuBoEO
X8Y8JvwIBtQ/7j/yLzu9MC+at3Vrc/9dzVipn7eoobpEeY1EHJc2i/JDzXxWwLEUJ1X4K70zUFMv
KI/f1WiaI2pyGKgNyTRig4umiIbP6mEtWdnC/2lyKo0ckYhlZHy382m2PDCJI09fFgfBvbBkmZqZ
vIeYZCpkJ/jrTDcdrP2ecHL+UV5EDOYSo2ijQGS71sqQiMUvErwA/YxzzoKzYQyVwA0zqG8ZJrPo
uZTQTamD77OhW0vhDe0iOjzHYHeGJXiku/hhF8A0lNYCUOmC9LNCUuIJ4bjZvPwzKAPPjXFK5ma1
p08ys6vyncAR4Sor2Dvq1IzrJND6QCQo5M2viZLKGyC960hdfCokEx25D/NQiUSdh5V7LiGh4vk8
Szmqpr7A8HxFYlYQQObdBTvwuF0bmK7QcHNddVWl72UD+0KiewpomE3eWGGyXvcCjdoMAGIYSUDp
q0kFWjuKVtgWDpgdKc5U5Bi0IWhEa+4iUvv7v281ArunJ+IJOwDZUN29yyrN9xda3vCvLv4oGEFZ
WZIV6+qKG5OmBSVzEPDKsATUWxHcKT0Bw7aZ6tywVeAWqAUDa3b0ylFsuQQ/ZnwdpbbEzZO+Qrsc
hwF8PKYWfln7HqbCvRS4Lw8aK7Fd056G0z4HrJjjLID/Ljd9xf0DMjqEZwEPQPYMOM2GgjD31DCk
y5nzGkfFZVxE4QSeV3m3P+lPERe9rMBi8CkF4kdZ/Xp3mgRCFrbqCeoasGbxz7Zb2QG6Wqtd4kk9
5U3XnR1JhQ0UGlvlCdmxM+IMwFmJG8muEq2QzZ0XZQA5z1LBRXM9L/vRLMqqecVUuBN7iXr9SeX0
MrIqTEEMnvEmwatJFR89G8tlZ56Qmi2dd4LWptPv4d5NiGkZ4qlKCaW/YBwGBbTbb3rrE3iV5Z7E
blAC7/V8cv+DQy5IJYbLhCBzH0hFhplIXQFYq6YR44rv+A8Cj/2xQ06OESjdt0s72RExKTXaLsOI
KmCMUyw5zCYMPq+AfRDDiaXOACjs5qE7Dble3MP1tiv3QjBdCAV+jcNintXCirZcjfJI4Bhb91Dg
Oj9IhNTKrCYM6ExrAwBcxfiwzSrrLkEOovXAyUNIgmqE/gy31fA1i9/D4ZxoQew43SHUTPgA/jlj
IUfKmGuZsJoFyy7QBkJf4FlfQ47Ui9zZsRNP5k/bsCiS4wsxXMh+dNoRICQX2aVaIJ8lHFDqVjR/
ZWyZyDczSolwdtsl+dEq73+7Xtxdj3/YB4Rwrzk13bQzzL1x0PIxAvsGVMWJdPxLprGiXGNQHxit
bGKjXAUhrwqmj5x3xuGoxfDu0cpXk6BviJi6afJPJUzNtBhoaYcn7/tybO3IUn/b+T3P7BB9+hUm
apJ4uw9v+HTthe7r+rhfo25Sy4IFDJS2hE3fV8HNhjc4TpvKPVSDXSNIue21EBgD3HGhCpaNiem9
RdR6r9jxtRMxPhgbXRW3bhwXhgvM605kw4bBUvE9I/EL66O/LwIMo1OH5PzQ+PTiY6QQwsSeAl6f
fkMRACZYm5qnENobiJEQ31w7cufwvH8oEx5qv0EKTer1zdEa5QqfBJ9xGOCAs+eqdczFtue1eJEZ
AeoRudRio/W4LRlX8VW5H++IHw4CYfjXMu8+rsrD9z85geRKDwrvL8edW/1E3V31yZ5Qo7GbGIoG
wDlGVIghpYskoI9CiqLdx9I4iIlg5PVNRNwTzkvmkfyWiMJukrXAgPD9pfGEhitRj6Hf6RYeYKk1
AL10BzPYVpa/SneXNiAOSzqCcvhbcey2k6b1KCi9X44VlCZn8RjPdDA5uz+17Q9FRK6GO8amXJke
aLsqKazvisVx10zc+Eq0u7yy7ldJt69OP0SebwMjgE9dmRraRzQ+BzNc7IgKZeGttKdv/yOQ1eGm
xhUl/n2RbBKBBlmtz+vWzIfiloO+3mqqCsvwlVTGjni9GO4uaw6ENgB2LZFNngv33+5bQ4krVBgl
bLYJGoVdVV9VCScxujFcX++VE2h1sGVZ7wjhQSziHnoXtNMNKHyD20im1/VMzlp0EcgriyeImfbe
fzlaX4zrU8AYXZ9mSIy+dA59faURvhUuZpgH7OJeF7E+7JOgrTixsFsGFjRoAitxlc9oH9cDOK8F
Q2iG8aFLTddIg+iyJX07ayEqeWhXPTjLQkO0QOkHD2d20AELPPiUyWFRHyc1HVOPCZJq8g1UT6Ni
K86Zj0/5mG1LJT398pGPXFz3Yny4f87wh1rGRftRu3mdDrmlJTZG4x+bFEuY+Q2bADtJCbFMQ+nw
pMbvqAouPqfJRKFyuueeWxlWzlGdkMtOnShJl+9257DnO5ueRBXDogarMxnNZ0z5LWG8otcgTqFx
bMp5SNnZ8zsKXSMe0cwrQf/UL4ZBPsdl7AEEXDTNFnslLGcUyBHxStCdopS+uQe3JI7ZqfzDskee
Bswys8shg8Xu4Ws6t20o4dtCgAumo/y9qlBhXzTA9aIQr5zQRwBkzovyVIrjbVvL0HXRtfkAzeB7
PEovzOdmZ+Y50i3pQcmlM0xdo5j0kogFECJ/pxWvHQek4r83MOtbTkRqiarsiKbAcgI0pfD+0H4n
nnvcrObRtKxypeNQMUYy5s5d6taXTYBPLZ0BKFMKoHMWDUyLfnlm1FJo2NMLDO5dMxmTRTv6KqIY
mtlbSP5Cjm7tdCGV5xhOLRUm4M6mbiKc0PU9GHapBgVeslym5QKa46w1jyNkS/VN4z3WRrudSA0l
YEnvQFlJMNEV2/jnrE1dTZbnM2/afSHn4OwAZKa3fDz6B7uBQeyXoatjFv4Qa3KYfidrzLTBhbJg
F2WxeqC1Tuj2LIL3O3T0ieOETPctaXBjGX6mggX+m9wIuDokBSgqqgAN6phmtN1bUE5Nz57FyfqP
dM+AQ0GORz0K68tueAjKJPSn3Jt5stLCsVn+aQPNSrW3FuEnXVWHfdm2mnPb2LgRwD7BCXxjg110
cG8VZzo1qragi4sXBbrJLG+2roM273dHOoD8ZEBufzN6PO4DGHx7Rw/INNkHS4iM56fyg6WuPv9l
rvhiNeS4Bo45BcKJv3CTrP0yYee0NB2TMnpMCUK4eqHFOiZVimLlq53BaKGp5vDlC45i7vKnanT1
/yztC6oF1WsfSFKLk+ETUq4bEv1XLTXbM9InhwpwLz8KGxrbFyH5tCMNphejpbgwQqy29mHLpSzz
AYTiqghAl8YFDmgVixJoBUW7Z3FwZXTKCDimSvla6xXbU82k5+UAzTNhsIE78AKkc+4b1LKf5OpW
8pje3FZRgcMBho/va5+SoHSzKoGbBpmJvTg/lbnYsIyM51JI/m9TlzuS2RsI/u0pA/47fkVI51ud
6cCxltIHLjd3xVFvZALD4ib0cXRX6zafTth0evmik8bENolLU9J5+T6o8TlkwQIQfV2aF7MWadXC
rIJdNeqZRLjInrwx6SlGtlFlE9cnl4ak0Gs6MfIKjIIcaBeLTAgt0lFCgHbzgup7YfNuhS6Bp1vR
BRt1FHbL6uOesUr1kptNiDGDDPwFKXorQoxfByoW3CaTQM75Dait/6pE1LukH56N8vAYvS6wczat
/K8cwYWFDdtZKCyeWW1pZVdfragIXKji/3MwhbVrTXwQqWcFECDlq+3kxV1pr8+1JeQ8VxSluI2L
z6007fV+CMulvT5d/aYsNPvjPYqsXcS/6pKsZcAmw6kqptr5tPJ0s78VaVmp8E1Lmhig0w+Z5YOf
hJu2FGJWIX+/7x9PqV6y8D6gLuZlvMSrnGdWGoUhtdTrR46lx1pkDJBpEm6aFya8SjnVVAX3fAGR
eAUWM5Xa6MtP1bdui2RgRbucyJQngMPf8hiFMTvnYf9nwTsQAbbFFNd5l/G8XquZF7EX9dnvzN+e
N9c66cMn1IHANpEiei7WAyIt4Th7owq/gDUnU6ZUNX4QlvfUwzlo+9n/Iins/z1I3PuVNLD4Mt1f
q3WR0IdInBf91Aa3GPK1DAWuMJLL3acE2d9Gs6aR1Usv9lIfS/+11rTpwxTSqmh8G07ufWssHBVP
vWKAL5QN2Ley+4EirSiHWDtB+o5KUOXrfpqVbZbJPRCkzs6D7LRsKNapocUbCwPTlJ1oilEBRfiW
vmS5u0RTdFNwqDhohAmZ7YsV0Uw7HdcjjWOzgrp/ByIhStSsLEDtj9iWmsJL5DUhNnMGSzvli1Ov
KLpWBQAB/1IAS5vCqcaBbE+2KMskoNYBCiRDYg/Umvr6iX5OEo6fCaINe0j6Vr39gNHEYqH+toQO
eQ+eQxAWpQQY6F9qjgHwqX90/iRP7D1kCbTLxdyUGIXJ8wt/igGlNjdBoHZljsOygHOPnWXIqYuv
GX0/oat/Ik4eznvvDHvPakyi13BoE3X5LIZKglly0oldHteJqYHj5zDG3McT0+nCOm0XkAFBRPWc
WX34kcJzIRQITfKDOl8G7gIzltZmx2s/5QvLDE+9od81MMioUdAbZgk8pmQyQaK7XHdqwXqmz2e8
EKCuMh+sYQd8Hw8dRVQJgCx+YxhLh9J5hulqv/DrojP55ANUWGxnfUAyMGcd3zsQzhhA5EK2Y1/B
VuLapuAvTxNiK28YuInMuaVSKwUTjA+zy2IUMCeksVKBLwQzau5vnNPVohULq2CI+emdzBjQ8zNt
1gSXADPAPc+3wyg3JLon3axmPJEzDGA6woaaY2hTA2gOAqQI7OdgB8F+jtZKceiyCJTsKUFA0t4X
wg4KexZm6qMTboPpTnZk9HPC5pzlsEeG0mvUYokjHnHrX1F9f2ATuAiU1aPkZpm/KmPk7LkzGvEN
kYMsNiejc0XymMtUxTlyBzdJLDqAxbDSVzS4Fl7E3a2yD9TR4WTR5j7eSvpCe+Xl9Bdq2vk3qOO/
zcwjG4tI6dKAOaSBmIE2RUCgsVv3RduHgH+LkYDW7m33U+xqoCBwuwN8dP/LgkphW3rHl3fE+20o
nNoNOAjWIZRu3TmT1P52mRedygn+W40sl0OIzG7g5OvCsZc5xR9ji8cB16O38vbJD+WuU8oxNI5z
1mZZxPNCZZk+a5d5hx30atvDx67TRY0mrUgfZ61l/EZdplB5bqNiICVr4vX3FM8RNZfiiJmideWg
1/oc5x36SJ6QYEZ5dDyp2AkJqYs8LEHlOI4l1TAMLXBgio10BV1gP0OdXgnEqmdqIpgqL7yH+1ER
7EL7JhxSMDKg6cyKcQdXx3M6ssSC6ql6lUD75JZNsPa4ojB4IUVjjMqS6YuYg6kBgZYEFa0/OW78
AwfIKcZQ7a/r1RWoYcN/gub02kLie+wKGdDm23JCrCYag1nh/DchF2tuznEtJlD/zbZMgkbJzL8d
YpACM4cqWto3t31oA+EakzhMc2U1r4iGZJv0PeDYXD+d6mQo7q0vUsrNyD0KPwwfmJ7Vc4ICpAsP
2iC48/4JoXWzKrxNMF4RI+y7ZpcUFtvry8OOVB86kYGRzxjkQNlypngk88rAVVMTONN0OO8FhmGP
Q/Wd8D0Rp5eheRQB+gDcy/AQc14DeiMDBiVx6SNFoH8g1x9BV9nQ7YKJnIhZRRrJlTjeQJOT0RO4
g/kDOd6KevgLB32OPwigvHj1pcmwrRU0hn/ybQ7vjCgOuj2gBffCG/id5SY/kTX/GHYsHqdcxG2u
cB5PjmjhsswzZBWjhwTMqUeUDYkFzPaYL0Px+ece7dXfRtSeKdopGu3RsS4P47ykgj0WE6arHUnP
JGRzrHCp7ZtLahxUxttQAo6HvO2jScKymrVqyhFzaBYTXaIb/3mtiq0ugIofQwCJMhZUBYnlAtna
qhPXOLX3TLL4wKg4hv4N8irL0CnbJj0IeeKyswz9v2kiUxfKzjcBJAzOobAyhkNVUrUQeIPcvpCV
/qpgsDfU6Sv5tbXaAh/i1UviVYErC/voWXUxU7O39O3BkjQIel71LZc9ij5eOnOuNOkC/ze95G2F
afWQYlL4xGxnIYPQHD8trhLN1fu46/s/uWrQ5PQLjd9go6XtmzIktdkWshsu/9wmCXbJ4/PpbiXM
qyu0ychKUoQSvS++cXZ7GXwVqUkKVzdzEyWvqKrbR0h+d6bPyL6lNflGMYMESkNEsx2KOY1JGtqT
PWi2iu687OdATcbn1jUkfVXCguxgXFLZA2lAp20JIweV7AT9oOes1vLkQRzIg2ps2Vffh14vOsyP
edjxuCwpLPvbQ+jTXsinHoAlXXkLTH2VnZhIlQYbpACU6StGabGaVMDBfvFA/NC1+TOWLEFb8CFC
utMqQ6StyTg+3YyCJijLKD5uiVni70eCYcPa22gsGt1pMI+4iA19IXftBwztTK037BLHpYlg1u7V
G5QsKfOgjLjQO77JUVI5H0T32AD31/s/dRiZVFrjuMKhrgh5r2citqC2xIXiOuCJujz88pntvS+z
w1svbz8G9pqu3SxEwaWUO5Qlb61Pb2nPf9TChH3p+kD0k+lW7j227foy8ei3bUMqBvvOkfYEWnpl
soqdZfBzOjvMnzSkCqCakO/MTDCscMu6W3ojZuBV27WcdL+ZRIblfNarURzZNZMNzLm/iGSYj6JF
zmRMZY/MaWoGTfF6I6uK9Br9isxAY0ug7HDhxsAQkItri0/nfWaedqRI9iHDaA3RfXn2T3A0bpGP
QtmKq5WL0gkIimokvFCer7xgD2AO4ChLJO9oAspFnVzwI1stZhmCTCUslStsmH/fOvjMcPsGt0vO
pVZaqaPQEY1l22fGhDtOjouI3bCPhLwj/s23sMlOK9SgmiAr6Er6Oi5viw0a7To2PrL/T2nE1i4R
Q1BOEYkbwPK82y7cfc4BR2ZflJStnpfQO77QKr9ubpmiZ9JFXmcYcuARxVAfZXzvlWm2Rk9KhWSS
r1IvAfv5bCQAXZ0CuSHf2CQ00Oi+BZp7XSx6RoW20hjw3/kpZn5IZN+KZD1DAUZgQ4FwHAWftn3w
C+TQDbFtBgSHBPuXF3sGlgbpvxuWovEgUvF4F602NLNXk6yb7BvM/GMLm9GP0INiPonUXvFwllRJ
3gRAv4qJ5XblRZMFMalGQXSBDUhWdR7BmhqfXW36kMEJspBXg3fNwEpxOKo7njUIGx3+fptmgfts
NQy6V3+gXH1A9/baiNSQbjr7upkRdrJBb7BH/geBNBlIigEc2KATjZmL0Tjkblt4qoCFswzrSIWc
wkfGwfkZyjzQ0PhJb06+yhMjatqRc/cSKnc1mgW6hfNTg6fYwiC6pWpUBts5d++WfH1/esIc98tI
mmay0xjylRSlPRCgOUGhN5bpwsTIq4peTgo/IVlqWxrW3+hc7AgQ3QutDo6W87B7cetw6oJId39n
vnxysr1F0eQtD06vJ9fjKnFI8mS6+dhuTrwCqpHWqYNoZjTNE6qS9VgovckV1hmWfP37W8n69Xoe
LAvuN82oIB55NMH/m3x6+EZSdtWtsjdU4fJq4wZsV7zjQO2EuOq6V14bGR7nS2kQfp+6c/1T+Zi/
Uw94nrhxOMfZ47NzjRI+Eoe6PC9n5bj+cbKi3o3TWd5W+vJEFqgCfpBCKeVy90V/ow/MdZesjncC
aPHUjqCJmffHIatOCaHnFBZdGNFHXoRhgrvmS5fATUMV5xW5ANm4sAJsdmsFdzM0/dmKj+MV/2HN
IWEqvCEwwf1aG8oJPEwA2znju/UZ1c/xcLLghwLuJ5xuStpx1zI6uYkqDevDmkDfq2Ardb84GQAD
nhqIyb8MRpPaUpscFqaisQ6f87HW+4a1HK1iIXChVPH9aFhaUSACGnFLWuhlWhNVDAV8JEI5GrXD
z/5I2cYsaYtzJZCD+lO7wf9ACOW7Oz9oaTJN/OY7gELLTOlykV2vbXAmyIxj5Qjvxvi+lxVLieH4
9iu5PZ5Oa5bLDawcJy1L6MQn5AtzgAzLQa/5XNexHU1RNnySCbRjNOOA+pn5W20vKGSfJfnwPGsC
DiljWyjLZJsrVMuZxWbCnX8ZrbFYSidnGLkYAbtKee+9wyKVUlDQjOw+AonYe/vlD83COJOb2k4s
cDxpKw5F3uGZ+8zIkEKJ4biyfq5POtgC/domFe/lixLaHrY7DYrMi40ZMfkT5q6mJEzeFrSUqBg1
J/Ay7SSMFbxK+XuqA5NkpKKFECmGU4iw3VRP5ekcYnd78eohtP4F//Z0oqvkldyki/YgCSBTmRYB
1b88ti+x1A96AsBkyiq6aflPUDD+UEuo7C89V1MHUD1SkFD8Hm3H8r+zQwL4tLn7Ua7eMLSuFGlE
SNibHNN5TIb1WET8CpGkysf8CT79IT6s0sl26poHp+r1b89AmDMm0HS8pqlMMwkdgoLxKM3bqIFU
B4KoxdVDIyaGG3sNH5g6gfiFHgtu47EnMzm5bA7FIsP4utLLy8LH/cjFAUxK+HMA1On4SzgY4G66
GijVZkOCk2RHjchV5N9gwuA1VwcQhTrlKNjhO2pgWpF8lOqxDI0qYOWLu/xlfDyVEgbZaFbdBef1
9QCkAyNZSwOVXSFuIWBYA/rfnEY170GvMCGoI1OMgdSlTe5phTlprODUx5BIXmpk3sM/JNgUic3r
42aS1R2nV5SWVTVHQYUJmOiMVGh0UlrTvgVktgDtkVgnxqHmprD6BTVIr5Ug81PZ/QLJtXE8rNaa
F4LKL8vcHG1x2JwfsF1L+e3jXTOJG0x2MRPfAZQ/446LXQ8FdJpxO5DiW8U/m95lRdULdrW+X8S6
U5O1199um0XGeXrKHbetaKYnqJTr2CpsXqwuDgb/a52saWCMy+4498pLDWecX8q1T1TdWAXYb3+I
2osnHkjoFOYAvkPz3JbEckEG2dzuAg6vP4Z+z7fyi+WIOTAjpklvGNj1GvOyUPffrGtFWox824Fh
5G4bGALtrY80BH2VsgzPNgUOcJO5oAZzxIgshd/Oc/k+BKIgvglX+CH6J2shuzQ/wUZNDJzaR61v
ryUpQyqXXkcc1Rw4Y5HyKGlv2he/o77HqiMg63NIo8rrkGdJEVaCe9hMJ1ERuBYo6J3+LNPqn3bn
hELKAMApnMHPxJmibkqmpTGNVWgYVxxy+6/c06O92jxEIjm74J2s1oECkF0ZSOJ4718ZbsxyVKqc
n7abeoU1NAtgTpnNVAWqV2+LqmDYkk6cMHUm9OZouEp6n16WKhooMbMFRwVXK8RNal9PEd8tzFTZ
IJ960G1ZbX1tuhK4tAesFxH4KO6J8PLEF/a6QRziH4y64Pnpi+WQLSTzz5WCtrzVbEoUaYAbIqKo
NxLP2PTtbD6K0Y5K6vHBQfWdoMN5Dli84Pzy53MndGJFRGsjeiCRh+st6+pkmoDfHJjkl9BW+z1H
5DjAneY26vLliO+l3+0ySxb+Ox8VtSu00e7a5rqZ3C8gioApePdIghYR/WSI872bUKExl1yrknmS
NiZp2sa2IgwmMyL/YhFuTgX/hujjDyolRpQ9LiLFj6KldlklYLDY+tB5abCVFJpiI1ui+wpSi7kP
ukmOMCZIiuoneAxYQLb3a3XAK7RiIJhhILXW7a5dBzg1lGOREKfsfJTxGNbpFa04TT4GyALpW6+J
rEI4WndSsu9BmKCgp5Vik/wCYkB0Ni+3I3rz9imWUqPAWBb0/tsGJNqTQhsKC4ytP6PobK7dpZ8v
6e95nXrZ8fyo9wlj03dyirEUT5qT1XLnRhh6VigK9OhPQX0YFb0uT68CIR9vg5rxiAwRb65Cn4Pn
dBwV5Zez5biU5MsgWID7ZllZl5ZrxM8qaxxC5OYTrLtZH9tC82FWYJsV5sJSW6tyFrYnFY8XWjZK
SUbQsgvHH3xIjOQ2xCGvjRrInAy6JFTqXI7/e9lVAUofoSopR2tYxP3yHV9wfsgIateqtfBOnTh6
AbKtEmyHvgJ5gRoWcjrZSPb64LvP74oWNhy1PpzZ6u+Vs7iAjZOOXqyvjDUyxBZiLl9QngIDgRmn
QYIdTowioZMms3Za9ifPc61mnuV7xCWamCfv2JLNeUxeGDSTezY4J2+EJ/peS/h1hKiMo07n1/Gq
tdEExNlN9+Qn/UslGkFfwhWEW10V6zbRUZhsd+kZHN+gZg/f3m/vG7VgcgtYWnEwkP+C6JHpj+gI
AdvijKNZg1i+jZaAo6VpAeR1dP5OCbc1xfkahh/8uxSFubZp/iqsRAZoj2AaSMmhVzkfQsV+diP2
P+MhzxW1m2HM+H8mMY6E66xzW7ro6HedCMLzgE4Pcj+4AwmwWiZRGYE+HPe7a+J7ZW8LTCAC39KH
E6t7wyy7DpEH0DXbgp58PUDKMedfboabtpUSPcPljb2XSNIj/pnv3yccRjaJxd1Og+jcTApsYUE0
eQeWmcNOwDWknSgFwCrpGpK666yAS/hxl98EeUghc2043DuHRfb5VQ77QasaOK6sLGsyID0nOiuf
FO8eTmbV+7WN0a27Y+KBHGbfrbWDc8A7APcqQIzhJX4+Q9MxqwjkQf1IJyRwYKtiZFtF2rBRGXzr
rRg2cFgiEgLPZ77rUp7A80xt/yNOJ/V40tZWJ63aM7xygrMeErG9UUCfaToSrlwjHVqO2WoWW16H
g03RFCHM+kC0fcLHjNQ8Je6Tm8pMBrCauyhgSedCAaGkPGzeZrWfpbHSpHAQOqNYjTX261X+OG1O
CyTbJHuw1O2nFwEmX+ceSznDGpwcF3f2L+Fet1j8x6bwdi6DGQu3RosPM22V1azDQC5Ff8VV5Aiu
VQXgo/lD5/IILnWX2wGL5bvI3W4YfHj/lkjyxUpiu0ZCIIyzJ0FV3qnttP9xV8lVhMtRK2kwklEu
3WxkXPU7UQUWV3n8JCCDYDaq8wKhwywmOHFxo8Zh7d/niRX40brIiV+GsZgf8qMuHGQsgggKhAh+
mGKRnF/O6Qm3pC/xV7eGXafSGsXF6wQamc6sRzWAMdGwo93DbyWZ6gd1JhEvlIDTJne1GDJ0ciGQ
ujBSbzCRZkSUK0aUoya2jpEK49ypfs/vst/AkzKOvw936em5oNOwq4L3lanZ0kTpJd0Jath9qTCS
EGWZ50/VOhbcA5yNZNeR1DQgBfgERKkavj2n2L+1PnsFqkNPMgh2Eq0osfjD1HfQdTpp4/PhYBdr
PDg0pZxfJZekb86u3KqHHsiEuPhdfK5WCrt9UAFUu161ga5gN7tdUrWztYWWJExQl/dop1t8W5+Q
w+is7awp5Q9MHvoMXkNqzqBfXHKbAjruEHaVX/tSlfDjUy7JgZ8s2EgP8EbjXpUiWpjgBlAT3iGs
rjICj05IeQWpSAREfUAwz631s6PDb2w6JuYSc+xfQ2lj74CX3dLygNS/GQhKD9YuRQA3l9noczR7
aTq/nCLPoWnZRujPV96eBGeBt+PCQL81woXxUXfqjbG+75dhRjZl3QiB+updMSkUPUN8pYtMRXTW
I51wa9nC6sGK2U+qqACnJN+OgYU/pPv+Q8G3We3f0J1mcJcEajAWXlGAo69WzN/XH6VaI6F1fpEX
/xEx0yw39b79TSMiXwLIJbDc17YSL7Bs1nClGwj3REnQrz8C3UIHRsK3JOIe4jVTZOnx2KO/PaRO
MTqWCePNAoqljaKrWw2cEHJH5bwN+YTyBSmZ0tnNdDtyx+zM0hdTNLLctI6JhZ2QKlnqnL1ljMYs
EpgQknZ1Dd37hUjrIovdrGFz540dXvQLXQxwZQ+QNvK1FdyId5QQ1ztfA91Lg7hw4KAUwi262B1z
j0UjypBrrwz1YRfdUHgQ+JR/2JRZ+pN4Y2LpHOl2sVZbWKcfIzl1ddgaSMg00BSK4ONvZs1e5u6M
OjSGTdRM+9k4fjFheJIIS0T5mUV2Skr1Lrtq29byIsazasgh4YdhjF91DFOmY7izhsKkZRRe7ISh
LzcDXlshqaqDMbX6ZjxUBRItOr1mIwTQSuureZ7OzDqZXS9wYEFgtMMOLVaLv057g0vSeRRB055+
DMdJd8UNvgiPJ+u+hqEibdWDep7eVF/EOAJ1OUh+IUgxSxdDJSmQ9jQuRh0fQoI8bMOzzdehI9Vr
X+Y8k2DKaA9dNl60vuGHkYWQ1G0pzwlnJYKzrxFmq0beCk3HxwXsvFMBHsolegTopS95ZIUdoN6a
IuN0+4/CAGi5nmBLeyOFKssGVuaFEe+e7KmnVinoj6Gkyv3jzgRo4jOVBOvt2ZbL8Y35IGLktLU7
GKH9NStPGtu/k6/5d1+VQxfyQngTFy2lvJQcV1kDOLukVkeA0aXT6ArbyUcKxB+nyXr6NDPvxKh+
GqoLRRJner2tUihll1Hx6GotSIStvQCLXspuf9Z6a+DjgBkAcPYqlAETf9BvOzIxkPVTDHwD4grg
cqvz38hw6wd8gdiANZcHL48+8fFLU4W9GK81JMVhQ1RGTbXhU8/girHO2zuIWgDLQvwUK/9fFg0y
ZSQhXnPRCQxI/ro98SX0NnE0QaVCTzhMN+yJ2b2pM+sxBr6Lsq2D+LOImTAVgrhrfEUJQzeScAXM
EX/plcl+xKv1GECXZ7sYOhBS91rDE0ZGgnxDcQ7gIMVVruLxr/X+/eO0tgjklMVwyaaG9aFzxpLn
lwAlGZlBiQf7OC8sinpYfKg3+tH1L0R/MLj6GNWPjdWQ5jwXs5ciJhz5pIT3LmG09rPeiy7w3CXJ
LD6MEXu1oCtsVeDBOSKM9Si/OeHlSzRGyUNXlpVWJlVlhJTaHzwlvn0mJOeA7sh6fBClWejyuV3o
NKcq71blXBi0lx47lCOsmwANYW8o681yIuOTREG9YCz7EfU4EAky4EFDFRN1Phnfk0A/hNLljgVB
cq4TJaUc2TpWoUnVQSEESUYXLLf1FQ1RH0+Era3taX3bL1vGKFFIXLhNNAlUwE09teNkbJAR3wjY
gTFm8snGRs/PzE2DIDV0og2aLs8s0ok9iMOc3gc5RpSTXwVwrKniXQQOe4K2rzAGRCHhTrfCL5w5
U9Rm6oj9JRV2Z37NbzO6X+v4Wmg4g3bkxqVIzm6rjRX5+/HNuvsaq/HlCu1KiyGfyXjEGg3JmT6G
kTdejoVJ3WVrO1RqEEZQ8UABMN8668IryqeuZkWqF7bnzYrgUGy8vUCCtbarS4d7OlahkVj3rkZW
nErjFetFWE6NnZvgnpj1ksxj+ePyKFljtoxr8lwye6vG7+6eQxMhET91g4a10Jy0xhJxzwm8Bebe
9xYbSsV1+JGI3RkFUGnyIqwXYh2Z91dmyA5OnIOYUdZZL1M0Rm9aINHhYxtDMCZRkHanCen83sjN
1LjJ4qQkQh0BP6NGMzgiDLwU3UarUIMk3uYoB8h8x90dRbJdXbOhhsARnJRnT8y+7pFqTkrhnlon
gfyc/KikLzGTXLxDuL5iGmVUKXjp7cmRqL+XPJLPXisEFDPjfqvUS7LWvqkh6EtnzZdfv2xIZVso
M900ult8kr+0hQ56MJPp740vQF0RDHrrDllRGTtooYYyUEQKppaoB5nJxUMbLu1l8Z9ijPAx0hQq
jt/XKIeaRzgipDIt3WbgQlpzF6F/FqeKn4265yftgmP9bRAsn06Bc/MhsMIb/qi/KmaP9KGHQYJN
dn4MmyMYtLMr+P8S1M6m4ShqyXoN2yPupNKf3QqsXuXvLe3ogMzkHJi0P3Xj5k6Kbmh58xtYNHpy
jabSuVIQdIqWkNZdTC7UGqY138vT3Yynesnce4SAQua/rebwttyhraYU0JZlHmU/ekSYLmIi/I2z
COniB0U7T+FRsPwx2sMiJzMPsxWQfz6cGgWO1jkZfdqYl58ELpkF6c5FxiYafUfufoc34Bq7TjN+
YhmscBMx92kOO1+V5zOETjeOEMD7kPLsDCC1G2qTxdPwI2+W7ztHf4wGk4yG3CX3wGJJ4qtpmGdC
HiRM4MVH1ZFtSKcCM8b+AdU3icNKRMaRjoVTZPCZ8xSbdjg85+pibGtEr+bCjDBcZOo/mBI68MJj
kZGMJCrD2GTWF2bTcz0ZbCICdzgrgtqXVf1/ygD9USTvY58Gs5dJknY18q5vln9h9AtWSIqTczXB
h+yDIeiJ4tHGDw+m2wHQx/3orjc3tVYcGmTb9DVP5dExflz/A2wtXKPxdFBQ5EO5M6honV+gfIL2
jWcjFbeU9P2a6liz8nocqBn8qA/sxQH6O2Tkx7QTwdBSCqiCaOdQ5wvRYujBTNpYXvTVe9ecKogP
+jRFiFkk9IdczVlIwfPNjWDmXM4nRW5tVE1cbY7KEeR9gRNoMDsLWhz77UBJLiSB0AhuzYJ6QRmJ
lxG2JxZv3NVgY4LWtNcNOeO7/RRTt7+lFPRUehJv5zJZ1pC57JnG+MdwoZ1aHVqjTNvkgfH12SkZ
k9HCPG0IL5/+83jssgxnBl/ygJWWfY+4xKM0CaA5+ec/8NqO2dFlFJ3KVZtoOK7gwQESPmYUXgEh
PO/m1d0hwDxHqC4gWzE2KyRQWFQYurn0OObF6UeW0UGeJ7/dGfct/LOFjVtNrcCGoebgU9WRF+w/
BWXb5rY9Xh9cXwOGMDzhr6zwiVWChrxDakgLmZ5BkRGh7hGdc1ZPa+0nOgKrwQxqjI7zAkRWQM95
SZ3LEiVuakSBnnc8F/9oJfWVJlUManK7q9ioVhz/vqKKG4tYYJKdBED5VAWKzAWUxIqt1Z3GNMgb
l1iUIT3AySNg7QxsQ8Pp8OOR0avwYoUnsnTI3VFmlZPrN+ViT2lAzu3Y+AEHQLYDpYMPkvxqIAFm
yhooup1kioRrhNTLNhfQJmDhBX3MWm47/cwDY4cB3SzkNUBJQkRM8LlRVG6mTH1d9uUj3x4f4cUj
k7+SE8Djulel31+zYuIGjFo/gpBl1njy2h48trvw81r7UT6FD6CpYLGBKmMdYRBMiW0Kzi2WYuAG
fdBmIqgjQIhCb3pSt9aLLv6VhWp9Z+FiofSdhpbI/vpjtohNNA0GAD60uZsJf9H2iTx2SXCSVzXy
zvt5UKWmFK+tA+d5U4EfjomzIga3QXpqN900Y6bpVY5BK5PNLK7udK4GUNloGmlE2kbi4WiSuhqG
/XmS91vVu986hG9GAZ7NGhRYx23MyacqTH5FbMnxU1VLPGgEc4lOLsWkULQkUqOhaQIARbBcX7Po
+9CgR+EtLORALRZVDV/ba9usFmz0XBFQ4ztHjom8a39t9VzHYF4iIxQU2+9rF6wKwLoo464miAva
gMtytPlUOX1nKKbkM0G+MmwgKebjBxEp++R7+FqD+89MwrRJfGinE4kD28Ks3MeDmqkoC8NO5fo1
o+GMpTfqN2OXn+DeKHFxVc7pZnqOyThbI05FN4+lgPO3dmTDsvGj4bEIs/9ByYTb9N+1SWdYakO7
6Y+slJnyv3u5nL//pthz29LsUWV4gSVL93wbWHos2xoGU6Ba1pzga9es9Vv7HSrkFkukFHXuPsyk
sK0wnofpywRjPSjZd2fbal7K5p9VcjmqM/nbkh+F9TwxfSxrm2N36uAMyjiETLTgncd+hZqeizjc
0DBoq2yzaYG4LKFPUHFdIoX7DrNDPupgGYhAHJn9SX0ZJSSZUzM/+jOAGlewBfoHs+7EulPzKA8+
B845ck2gqnXdTnjM/Q37TK3CVyx+442z0BB00T4vU533Lo6bMR20NFLSYIc48tZ9JYfTkwQyoSgO
hldiRD1KX2HvxzOqpQ9mR7i+vTJqZf/z9WkJm1rwpJAqKBgl3Xs8TqMcJIWmcQEYYMP1Hp3N01HI
hcLqhnc4t/4m18qBNVhpkM9I75swp9/cEQ4w567TU+LvaJpz3+kDMBo8Qke3BR0HDBwH/DGd1i/E
5zZoCOBG/iNZRXhK02Qn23ImvJLElcrNH7R0a+DmryqRv6pek+JrrNmFB3sOfNla6uxtV+B15Q15
8pOCvqh0Bf0uC6B+N7mLKQiTuOPuMgBXs14gkHAJqH66d0lWSIzI4MQJ1Orpf2ow4A1t2PQUuqNB
VsbQzhMK4qgXz0tONNIig2Mo5zMKdorPfTRaSu9rfMzBbSlkUhX/kWlfn3V6p69/D1dDTMSJg+zh
XU++finYIcgmhxolRXd5MeIoVBEgKwhV7N9zKvJfFWE+8wbNf1W17GRTeeVg/TxaDezw2hXrMdSG
x2g+SDTFXjiA7y0e0jKKJnL/PKF9oGd4IvbaUiCaMjezyOyyObNVtR/EQ7zi/TGJYg37UuGhk+SD
V0gYQpWnpzop85urRCpmH7fKM2yHw1DIpHQ1SLB2WSG/VutWFUxYqjdMCCHEfhzss7MMoNEUb3DA
J2Wy6VXtCdVHt08iOdJTpT0yZcMLGBvzqftnlg7kErwcl2+jdrGfltGsEhsh9Y/ZSdT0T/Nk0GOL
LCi1vi8HmUiVI0wk+yQRMyTrbDtZCXScbFCyIJsZWhOVGs9AuUuFxBPKUiIoN2Ol1sn0XC/L96yY
8Bq0QV2z6nZ8jN2jBUHsB9U5wdBHtKIGmwPVvv0g3Hm3pSSmr91N4uCqt23hQXuOdLdeWgxjWJiR
eYEzpO43wbHjjYp0GNpkAK7H/stc1Nm38SPPlZ/PoLcJlIfM21zmaH/Yfng+34VtRbUn7gv0ZgRn
3Xk3hWM8xuzH+XosakmwCHl+POrvI9HUYZ97NQG/4Q5Y+aHJ8ZwMgRzyuiW31rcXI3Q1TwBQqwmA
2c3oSVeVVmPKFdwR/CBM5/3UeLHc7d7K1c2pCBkFE+mFT+GErUhfu70HUvxmtLXgyrKlFf95r3mx
Hva+NTtuQsnWS64JXZu6HWKtcgCjzJmusAZg5zLikQrF0fyvXutzCvrCFeCObmN8kL/qqYIFA0XO
hwTlv5xYx3dIuFVJthb5uoihDUZzkWT0TlUoEIatrKFk/kUyKoPvUigRRThY8H4/SBSQUlTNbWP/
kRgV01iX2wHJ7GwC3Z3gRWfUXXXkR33oAjHtOY8gkxMUA9c119GY1tG4PuNHZsgCTF0rqP50PYIK
1+qQU1UxZiEn7FPZSx1Y8piB16Ggt2Fv1s/xRoFT/nssayOWosDbPJ5kXDrBNqN+vvgKjmFemq/c
+Y+/r/oZQUNYEQ/djUh7Q1KFNEciDkDYD+DjGpQ3C+a0uQFt2jnbnbqAtlNVzlQPMCHe23W7Iqve
J6qjMe1geqKfyeNr30davDB20QtsAtMBvCyIeJQsfYj9UpeurajOO6yiVUUEo92nhpBWq7wyknIH
9HmhA/GmYKVFo7gkYOUs9FxMkg4HF2qhZGaD0cRPB92mFyNaLqmiJy2SnGwSqTekKABDyC1Hbaar
/86BaHCgOxXcVW7q05bGV1i9rqfvDhaFj704b2zEuIV4IHyJ24eIdV+6/dij7LFz+3Z1kRwptZei
yJHFRGehGabyzhTOgTAm0Z/EQ4IajF+bYK+sHcVKO+NJIvDtiSR65FCZbJ8xPTxvMINvJeD1DaSm
4lsrLI+nHmC9IWDsEL8NKdX3z/aVASrX3Xf73RTNNqUAy8Sg2OMEwLZSTtgbDA5VChtuf7uJ4V1H
zQgckaWbQy4LIQw+zSDP2uk7S46bLAnw5HDPKWkrOFLI4StRCt0wlmH621fI6dM2iLxPSGMtciho
9IB5Rb4ZoXF+aB0//1LrPQQSGFR1QJKzU/FzHxWHi0nx6qKP/+RL0uSbbk03rk8puvtwaWhaJwa4
zWe1YNvrI1xTB2RjBlMFCgpjLACDwySKDC6nVhQp5EyDtcZerPLn1NBP31Hr/az0/cCFPb/H5J6y
f5G8idOkkWvx7XqqL8cfPQynkGKYnbbzG9dKbOLafieSue1Yj0XF9lltqUERoazgFWWpm8JOo+Pn
0oc44qGp+IHNqRDABx3Q8r8e/rZcSObZtX0qFmnyXJnzRt+8wHMGYM6C0ZbkloQlFGmyMbTLJN2d
Mx3TzSF6kMoedV8IXBM5FKQjYRodlaSe1HtNH5+ev2k+f5jfVkfHiZeH/7iYSjPH10YOCmoYvPDR
oxPONWk+VXI/GPq3hUkeSnvBQ1QMyt0Atr1EngqGwfcKIljBH4YnjA0Kq4jIZs218M2JP7o0DirU
hcR44qPZrdEB5G60G83jwQcUBIbM3QO24+UFYCdaDdiVSZV/J/KwdzgmTq9h93DW/UDdwBIym0CG
FrCEIxcTTx9BW0vgPlrKHSSB0lGIHkSGX4Dkgfu/qKC2N47v9ubgCs47C04z5R4MhVsaFk8KIFf7
a4sfKzLfq8pre5QJAVIBB/z4fOrCiI9sTRcn7/eLzrTdIom3BaNOyLfW1GulLGtdQYsR4iNa083A
HhJQW1wTYNWCL5ewfgDISHdmqZ6bxIEoCRZeGt2erwxgW2G5GBmNG8mcNE+QLYg1e2JwhNcacwCr
sx1yzUWfZ89nPOym8/hF/lUz9I9uNJIx/AKaRKJRnJ6kuTYwAvdUF8xES0kt7BWRsiyOM7Xz5mRC
B+VRiVSfQGvJrh6XHuorx9G6Lz1S6v6v0EDRKHR9uYi16sI0TLMOq6Whjh7GXjKjvpa9fIQ5EZ7z
lObLXuddPsR3Y5sEzvAaeoGwPpgdHq00bp3aueJn3Yvnk7gRVPYHRO2Xt9tH39hUORqgm6oWyL5U
1CiYOznCjcgezfuaygF7dKbpfT6DBTEu9+YMdAFKhudnpSZdqaWHlyBJFCnxE3bm5nMYuNmtS4Dw
alyvDwXbfL+XQPgUe0bgE3pLASUoHZFmAL4AO2UBnjqKaayeKDeFgskOpG8oZFg7K1DXf4SJtQ5I
dAlBc4joGkHa76+SP8rW4bomrVF0iqzacafK7XNAKQjKa7eK6ZtCyJWQIIy5CM+vNKgw0DSzuyHL
KC6K/2fKlrEM5gKCZRX1fAaoHe9+dHf6s74awJpG+6W/vUGiEIQHHDoO5awjmwPV5dTg47otGrNf
SNa1BQs22FHsgOWXCqsY61DU/oK3lZ3NPaZrz//5YYXk6KvgQzwcXkdj+n02++sRp+k9xUiux8+A
n+vf8c48p8TOSWRGw5OnuOwhj0WE6ad1FiPXbKeafvCUmGzw0HOMAgEeIaEeC9jtQsDbVcBiFhBf
rHQoXRPllbRbKzkJQcp4hU7quiIpj0kvmXDsKl7Ne4rE+YMYhBM6tkFb98QrbZ0FbhvUdMJQHHm4
W98UCA43bpS68y9Z8VMA91WeDDSgnYs9AFwGVOQEF6esW+vfw0NEaG6fw6a7ev2wTiRT5oVH+DXs
J7C74MfuZDY4sVOdJpuhyIQaqkYlIAu1Otiv3SdGXvsfNPgL9aaajsk4sI88bL6x1L7O6NSB84Ku
Dhka+qB6CppfwuE5PtnRqG8+Y++BnZcbjwjm4TknN/dXVLaF54h2Y7wmueIdt6hwU6Qho/dmVSl/
irvZarQtAESDDjqKMFNdW0DMTdeEkU/ShzK+FBu9iDXqw1WGzXttg4EZVrrXogZ5ojYlb8lVxy/M
acgJ82wOH2a2sHyf6ijR+gaA2jNgrOpvI1/lG2Su3zKzwrjDt/yPpY+YR97BueFSZ3Vpy54/YtSV
931Cngc+IpE1PWAHGYzpZ6/sip+uOhGsEzYkwu7KoCZtj6QrECuMLYLJ27WybfdMseI2VgIx2/LJ
A1RY6jMAWP8aKzlyWdb6aNW7F6JhQBJXbA7FR5bsd24jN4EyYO9Po5un5o+L5Wz0ypJuY0YcoaB6
HVtlTr8owGpdfbXSxpM8A8SHGxATE8usr/8Dze1I0ChcFHNa9QvTR+BbK3rOKqJwVVZNCCJvKUQT
gl6JbndPGykoS7uKxRfsr695YwZnD3msWTs8l7dAUGeB3aLT26wPZkBXc2ln3ztRA9GD0yyeg1Jx
939UFIfq5Jeh4ocjPtCKgeLNsYjlJscbPNyfqi1QBBzwITAv6veklJW09tr7qkusx6dOvny3Lm3f
VnKjUmVLUjQ++Z88xo7ZV/A7ycQusNW7jgtOdFp7QTvoaRDDwyDWmda1lOPzY9LpuIRcN0ACYsVE
LIQjHjjKn59gnXhgzM07ODI77d6y8Hafbj56EDt2IfiJyzYLb9fAdOmJnNq8YrLh6BZmexA82ya6
AwF4GUZb8efsirmVmsrrm2A8/sq1dZXU1tbHqq3NWVfK5rgDOxz8vAKW8vf9GrmEXr9V3wlXALBd
dLEQc6m23ah70QMZEtV3yAQjrBLRUfd2GsfZh1rfUVTIc+xkSXqbqoYjnrKtgqIImCJ56x1+A2fh
dQRonwYui94zAszVul60baTD4m2oWqC5v1JVYr0f62ImiJkTMYH0c1/hlazyHjhD5xv+608yuA0A
caq5gbpTQb5crqJHT1ugNtL8MJctD2GwRHDkJnMEX0SnBakBqJ/61J2uiSgI6ERlgUMMes54zG6L
sWS3sox7sSOwsf8p8pzkwjlTDFXkiQqurbjAgv56MlGs2LGyrypwmESahNWGGJplj1RTFwzCi3s1
EvH5TI/ipfbmUf423EztDvTbQvEYLFef3G7T6OBiZFiirn2GNF6l1xsuq3RTBEBxbuoOhgyUijXp
4n9QqaLGG+csCeoYj4D4SQH1M9oPJu3n0YX8Vq9udAVLSCuJTfXB1GoadWitzhB8S1yeCuwZ22cb
tmtJEmEYUTEHZIc3iHFZZblA2oU+nmTjdRAKLZHeM0Sk7wJ6kZTgvcCLykBWFaeaZRzxBW731nF6
b4r5FCWBUClUCB2muSJ6yfhNGpWDApKiKWKrrqoYqxw66xfn4BLL1p+GqXMzmGAcRIFcOSKbQYZJ
okCe3sVeo8moNUwR9itOR+QfqKP5LM9IJOpXZcn47vx1IwVBksx/f/lZWTq1Lgr0sV66NmYfhrBH
Q5OEB+7V/ZQysmLV99kikgtYY8vYRwHIQ3cAW7f25pX9/D3PX1NrTz3UKEO20JwEN/NrkZ9DZ7Yf
ksgb6KWl/8ta3Hj5FMYo4y8bA+e/qq9j79koNjuelL47El7p/39Jy48+G9N07Z9JhiG+/PcEJh7A
va2SrdFsbQkeKlNfYqt9jOutAhy3mOTLz1jMQ0shd5Qho6UNyIagJACu3ok308yZnqyU1zSRhGq6
p75azWq+6FAiK+OWngKEDHAe1vN0pjWQweANv09148bxlI5W4ueQvT6PmOQDgRNVjEegxPpXmWbE
Coa05zZagdNM3joLNRSe4pG0dfpkeVxrAbYidE3qZUYioMkvUnu7IZ1QBvDC88HEPHhNIukH9EvI
BAyrImSIOlTzlztPXx7izdabsx3wSifqLQnLiixQXLQFicwudu3HzZy9QZOrJML8HJM8pNWjSetF
ctnFu7X3/0X7HYndlk84R8zB1tGlXczdZ9pQxqXvnSXx6Z5/THXJ7Vt7rrvEKNdHKETHeUuDpgFZ
ap65GA26DOPH/dIIfezsEnrfpI4nQH2p7FGXNWVPze7F8HK5cWS76FBxNGdBvUmqDtwVayvxy59U
EeIWHGvsbJ+bIrezvKdGaJi97PcFji2cXUG3877TTDiFGyOKGk6szNlM/obpX9ehe59LMlYOzJQ8
NLFIdHxob2nBFWga5ur0mLsB50tC8e+21Dr/TX3q+mhTJfIAumJHmPW27Mnge4D8fEtnhRrTQV7+
cR1AYuon1zjgoEZShr1UpsvaSZGylWELXdZoZa/2XwwkeDKbB8vCWHzR87gzCn8tIBBI/60b3o/L
8Lp2HIls2mhjfZDvZauMxsOmn0WrQSn27BMOgzb9j060h9xMEFVnaAytR/0DISQ35Ywslg/MstQE
uLH266TMaBFohtLTO9j1uk4AmzzK2tBRjLT5FM6thIPBf//yII270M6t2bHTz5tLR/9P0vl3FSAo
surFVe/UqFRSPtv5qvlogu6ovZl7idmKJd2WlwhhQR4M7hiJRxMFySxjyzQPWySYlgFVCp540Xcm
467m1RPJ6kqbb05dBjn07BElJieTwsE5N6t6NkuykXW2V26zauZc+bpg9mwGxCGpbMNH14SZsVkJ
CnHqmveE+Jgvd8mRseniMaLDnbqQWjwcf/7hqmQ/SoRFTv7qezWBazgkyG5at3o5CtBpzEDixgt9
JHn4cSsJs7mGReLZxrIaJah/BYto0r+AARXawZG1T9Vg5IhnvNV6ejPNabc5gveslkRcFS7JjM9M
4sdKkrbXfkuFQ2DvLRmRM5bqOtbZ4OjylC9JPIdWv7FhogXsLGPHOot+mLiLrDR8Ekrtkgyv93nc
2U8DVih3a+y0olsv6NBCfxVAYUCetNzyWKBozs4qurDS6h+tsYh6KkKs2bzMNnXn9sZF57OoIiHG
vyUeIYAMyg9lQ4SUZPfjWTEXn76MrPbvVoaoRjFCWtm85J2kyraz7DcMVpcVeqttj5iGNC6u5Tf+
L+v0lUQfKpBIQXJ5346j76fB79+03ClKtmuttvHduEw3KrHXvjfc712/RdikbU3ZDJnJoab6fpAU
uO0ZaHGjgkSo7+M8OBRoJDP9WAD4nB9FUaigLQWv9+zCMHmKNLHRYXMVLXmB9hVNgXWywhLrySFe
6qLIfbI/89w+/IOdJELIRsLNtIco2v7vqgdgU2nY094cspFIX0s+Dxbu/WrOLbXaVtCaN1oWIR5j
AzkDDX6BwNJGy/HqLZ0pW6NXL/5/LIhM9iBFu+BrRBNoLnEszZ+A696EDSvSzOzvRBHeVPipDMwC
xqayNVEjpxpE5BZx76NWut8Xfpo2V4Gvj7BcmCJj3eU2CXD6AXyEqW6qe4SJ7Pc665LGMnIuZaOC
uPN76ezDZidV3OapbPmjYXwWGGHa1gvsPsdhHRmW1DhwzWGa0NnKnB1tygNFcICs3boBm9cC5euf
Uik8SKiwkCyuK1p2MTjxUBJ1mrP29hggFKuDVZf8XZR6ErYwCWK/tffQ4UvyQmoPdAORn/DO1vVn
WAgCpHNKuvaHb/imIeFC6ave8vVT9GkP731EaHrlRh5pIH35lAdlg7vDFLro2WMS7yY4g6dI4xx1
k/OCKWalC9dG+u4Bd/qjh5PnMnLMImCOOudrJG1TteeXXuDam7ytS6UxzrysfPWHYpUWYP7JImKD
xHgdPTmR9p1y2z977cAREzz36OVqw3c9XBtQJbPR7U+Zd+moysDjP6u1mt7ZXbubl490uQjs09A5
B/UQeJ+sPIj4/Bddtq2nvY1wbSmxuBOYAS15jJz/ctqStmC23/GolrxVx+J+pcDyJqGH/ME+dYAz
WrY2z30ACqHuI7Jlwbo19pwpJxyf95c5ZVyBkiVeHTnnyk3jVh9WpwWXAp0CsldHuKuLjFcljE0f
ueKiKjHAwtuG+WH51eFHK1rsnjfFsQotNDOpTj8r/vreE2svoDSeI8URMtacCY70jiWvWjDAjYmH
xgme04U2gQJDCpUfQ5yKSIxbmlfxcPp0rnL9GZtXxSQIEQkFSLT/PQ4pilryC8OlSOnBGaM0Wsmu
WQ6QM08EX/10pby2CgH4UAbrVO0kKfd/VFHrKWof0OBk+Q+eVvfmQyUfL4qh1YhPsuC3rfjZc/Ey
znHCUft8YD0qrHcUk+1U+j2ZocIi8BdofumJDWqcqyYSlZtTZUcV2APHIeACxsJeHSOT92Krzlid
gUzVH0X1XIFfYPAflVGp9HLHlycZqC9YVN9FuNMHeDU0LMlMmI9SbnpI9fwy4X58yHNrMyDW4o84
PvIBitdU/DO1Ob6b64fonvzU9PHuUxnWY0/GDrzO9gZAf7OHh0NIzvNnzyYpVWtY28tps13AzHWQ
KvdRpd0VibsXlS0urPA8iINx3nDdeXhBJGbSUAQCnvw8bH/DlQNwrOakWKphzSV/OkREPk7zkXqF
pf5qim4P8+n3hxSrHhRJc2g6RocI01P6s3W0ZmahIOa042kL+OrEvMQX5rEqSbVoQ0m7nlDdIRSy
yUVnrlHuQNt46gjEPoUuxeWLRNquJ6yJ9yXydhX7YUV/GV4aU+N8pIp7lNHqEg9bOVwRJpNcZTR8
x7rHbgc/v+aunNUOCnj7Txw2lbne97dYjDyhNkIJo0KBbGFCK1wz6C5kjTQ9CHkDsG+Gk9qk+vHH
ToIle3sv69XtyJlGIYjCmXfNch3xdvIvPoYys7WrBFf9bLnkBB+WwZZvsm/cz5f7n45UZJTvUyit
i5tSr8cmkqWpFxvK8vm+eD2rkRdjHaxOaIy+xbIhSuM2u/ZulWjIFcaJudgLPfEskORAcN71/BxV
bPwvpgnivgLUHlp52f8oFCtlWrxvp6KciYPTeKl+ZtkqiSp2whjcIWTbrwrfFKFZQmwK7UN8pDZB
PTeiQe8GGR7vWjlY657IW76gNuFW0GklHZscpHPF+Zuos4OUkTGxAagakEfCIe8e9wNI0Eq+Twvv
Em5yqNKzkrI0h6pkZ7P9UuI1LARuBxLmktpWFcTyAK14Ir2eQuwUD5+zKQWQEedtgqOFlKylxXEL
vj0Ps1acQXIbQyYdQuvPTXhKCRSAi9spNIRt6gFhG8HGH6tHxcovbrudoOHNzBhHrYlm/G19SWCi
BaKwH6D4JUyLcDVG9396iBVQ5k2yzOaojCq+4srg4YxvPeCYKyB7JMpM21lGmo7lE8gFTVx6C7cj
QIo0MDi0mmlR/nEgDMb2ct5SYBXFKZD9x95QOpqJsojS8OiOF/sFpDgoSZuKjPWdRaBFNrKC9eJK
snlmGq34ftSz1wfg5xHz5OpAo7aWmtraP1euGyn/+zu5LMJZBdJ5zXwy6jnLrRqZw6AP57bN/USK
tnZlQY5LL2HFSlkFlNt2X5RobJAzbrsrxFXOo6uM0oBq3pDe8PFVUE7X+1zq0M31uPQIKIFx2roA
Tegd6iSj04tqJ8Aju6kGw8JzxaYEYVpv/0gS4LkQgJSFWGLDE5Z0TUBxnZBRPTyiO1cV6IwQwTSr
gbF13KabcuGK5lg1zNSeiH/Dp8eV/+mypYZI80XULHPdABf4XmWeyDEn1v+Gfk4wLWbTBowaW4JZ
8sGYTN5l37eLCge5Ly/Zqq97lO63Wyh8fiZqJX7N5PmxfPek0MGkKeDhunQ/v5RsmWp6/YXJ63UV
p5CLmwfjU9NHMg3rdQoUIL+5ESM4gqCB5HLTDhY6JPXinIX383Z6txpg2HB8Dql1AjWvgmGPwXU4
7K7OauJMDdRXReabV6aOK9w7j3o6B3hiWBMy6Hnv/9gcWIw1sGtBryIzG386S0evPM3EzLLMDE2A
mNeIcQ5IUSgvFtnt+6DrVNgs8cf+OibXaLF/VMEDnz6+60Gb88rCSlKkZiY2/pFH1zeSJo9XE8YP
sHJuSavuNsxlffqJIrhcJncMtGodN2gKfnQ+Kw4yGIHmmhjWgeCi3L/6MHNdk8SkWtUXPeRFR0VX
F92YGOfGwHuHtnk+/RcTW+oZoHVQyTgWE3PJq+6x30rwohT6Qgg6KfXuWe0tCAIaMPGan2FkvZs7
23N/i9G0w9PYAJkw+EjRxTliT1vIJyyDbtq2dpyxwdhFQvcq95eyUqJt3IiTyS7EVDd1PzutHViW
1CTfCHx740nlkQva9Dcyy75KgMvN0tBo2HJPuMja90M5r3EpYg9CTs9KuM9BfWZsawmW8kXVWNY3
Z+cjvMrE4fQFxfZTy0oXqsbmqQpfI0mfQweXO2K0f8m+DsonlTsAwJct3MXDSvJ3+k1Vhe6vKiSw
yWs3ZsDCaBNh5OpFzpvlkuy7sTo9kwUbQTO4prWSXjiiNR7DV9/JxWqvX90aXcYkjnX4s2cfSuMu
VBd84awjDwJKT1THTcwp59J/WOLVWbMQwocXQ5HWr/tTLLjcpavoTeKAPDXHjj2E7h3UVS9nI9JV
yWHoC3d8ZIh70BTJJkNunNAdtmk7qs9zbYy0oOGSyM677WSSSEaMBbX3O6QD9PzRbTshWCbfEQU2
CjbIUfmtpStiHvJKTDyvLw7ocRJflFSzBrdPsbEaOtNkPJ3q6bO4tD5Az3nLyS5CbpG+hPacjWfY
8lItx3vS8FzyJu6N6narvkhcK/GraJqiXeaLhFOfXe4ceMo44V3PMLeUrRotz2cnIHqlWY7Us4WL
3bZzbivzFcNB338tO/FB8swQrYn63CeteFjNvEExAAA9cvzWaKLfDmZTjXehLtMvkvjoVi2MNyzi
65wkZYjROTEXl/vFVSBkk1L5SnAwPKHKrLbzUw4e+F2xMh9Lj30Z2dGiHG0eEOIMJs9DBgIkGcWR
iz9WWVkBmX2HgJL1UEhbBaVsNmdhEF5id14S7Aw8i3QJcjKwBlunYGgYsINB6G+pDR1wBxBzqx28
EtnbtqWgkTV4Rf7i4zrJl92UyNvDJ5DBdZYO3E+Pij0FHT1bucF4bPP2skrJxW1efTw6un3LYlcH
zqEN/ePbx3Y4jG8QlFLnOtC0DlP2M6ubiMXmPxnbwWIO6+ocsiZoJENmghyP7h/59Fd3OPdN1G4y
qXGJAy/wRXrcwk8oFofxZN9+bB3nr1aRu/6f6LjbgnwEvGU06RCyg9boD+p5/nCMxbCxfV2TJmM/
hatk6cfaxRdrO+xMwKOdc+USBN8mRjxQxR5XSy621kSNPwmTxe6tlDc6hlOjeGuq7it0RtvnhA8e
vWUmfFouDAVZhX//0uM6RbcKZIjErpKJPfn0Pd9SIUmqLO0gVEPmZSOvGu9dW1iZ1XENWMogm0k2
6RsIBNR3xtp1otN2XE5bQCm/zP9sHhmw9KdC6dO2FAsDdjB+SmOUqEtB1L/3xs0C4Qf3P8RD/oEv
H5DtS22orDuS+YLvys73C1xD8bvp+4fHkFxxofzHVV+CScs8uknuI/8KsKwHEtA7beK1vwyMQvOe
otVJ+RZpxRV56tKfDUa0WTui/Gzm4Q0kthOQhjb+KPLK3IxP7MvJ25s3is4brO6x4W2+8w12GP4b
AAD18U5f7eK1Jj8yMoWUIZ60+OXCvJadT/w4VWeHDcB3VH6f3Yte6fEqrx89DECpdN2jW0cYw+tl
Vpf7q3e3AVpoExdPAKCBVPBo3kyDND+Ecj/bpVYAwam8eADCI4aiuRTpI/y94rggfIYagpx/eJlB
HXN6u8MJNk8T0PLRWuXQ+uKMXAXxtFZURggT3oGVOt3qWiUIjr887uPuEItZTtnMy9lCJdJaRL0d
x++V+4S2rUePUjEh+hoFJQ3a5PCOc3KeXP4P9pApDxWquHUM8SZMZnClX+O9h4mGl1ujCJhHSUXp
d2I92x4lHLDBczon/uZM6+caLy+lsMGU50Zl2BS3iVmXVGjvAy00WxroVEBijOevRo0o5JiRp2QX
lzf8HAevuMEPKA76FXn/4ErORLTEt5CEXUuhn+bUYcpjiM038S/0gOeaxEwaXu6au9imK9AWLc9q
GnWRLy3+uyRASQuSnwiwlGoNMzcuhdvKoob7m70DplAX4nKQzEqEmJ5gm3VZtqxGGzJIDDdzVsFz
TGiSZcpa/+6BsYBg9cy7DZZdybWmPO7oYVddslWcs7WCJ3z6C1j+EI8Fx5HKH44mijsi8hml/1hb
pnpcRBAAk6yUaWCnEyqn+l6tzdgdN+g+kyEFcWLT46p6qKwqD2MKlhy1KVG7HXJwxU/6nJ5DtJJ+
aFPSibErpsDNrJT59WwfZF18oxzSnjR3DcrV1UrV5v0XVnA1Cwz0lPZ8iGb4tAFN0W54/DN8WccA
3nV/t8Xe4EDJC4INBg0h3c1OQAmN0JwZteYTmT39N5BQ6VtVzs7RINLN/sTWshNUwhK7nGao8WdC
OVRjTPPD5ReQkvodYx78VBx8iyrwpspYgEj3wD6tG5Rv4wflf88xPJECnMpCg3FBJR+hwj59rsxG
1rD+gXTlOce7ZdhKfd2u7hrF9EX5b2H6MPUPe6woCWH/UPLFFSYTKTB1G7Y/YGUQtP9SVg8Wos74
l06SigUY85Cm93EwN2xu7t8cB44dmhdop+ynsYUKBQlI6zBWaK45Gpr76SJmxHTorMPQDh5KppAv
W4Q1MrWACOpq1mtPjEJNzkfN/jubSk8hysUVj+vBkttsQ6KfFrFAkBAHieXBE8YOMGthZl/DQNFz
boUNhYGxj5B5cT87xtXD60pBwhqJ/uT0tp3g70CPHW4XfnQ1Gg9uLmN91QFIZv23cKsjTrok2tEG
D8hOrtIDW5cE/aF/mFZTSMXywf7gu4a6g7mqKelsMoZz64VFCMoVg/cMOiW2YM6/UfWqZEZGP6U4
AF6KNOLuxUHfkHrjXBQXjWZ4DWbsqXIOegvwOL2FOFcB7DHd4daLkwsADbpFW2MnyksQMZ7yV0M3
Zrgrv7fX40XVckdUEC7DFeCroWdtSM/jObGJMrokl8Qgl2etez/kb1caOsZg3mW+vTh64mbXz4hY
C+bSXDgFrdXpo6dn5Tv6VnQwi9xCPBCF/oGB88qy7ehuzmfrkBCuyiDZuASQh09WetXkJFTcYK7i
Mp243RlL6hRLDZ/YeQQTm38yD2n3DHf/vSWgG64ZdiL48LNG3/iVaHR8mmeL7vxCgqrMDIXJKej9
gMPe8TOJ/m0ch3T/wEuXV5n3j39qynKkxsKlvJzkMY+TpY+Kxg1NYvn9lyyWx1zu4lkf8EKhTVw1
b+fd/UKxGWQoCC30xR1RnkRbSIp/+bfljKladckD6ex1GQtVwa8VtVl3og1AzO+kZcho4m4NA2m1
/PWoAv+Jv9+RSpgFnzydnMfu7fmoLCm7kRykXCVqELNyvfWb1clrTplgMRrVlE8TrjUbz/B7fcHu
q4+yRuXqRUIxmwEj/fuGurLmHeoNr7+0WonXkSPriez5dP+dSBMLnaTdRIhhKZ3zyyt9TTqmLxVZ
mDibi4I6rzyUkswvQbdgkbW4PW8zbbKtyyoLTcTF6f0YPqJMhbrf449CPBzONjm+OB4LNfIUasKC
n79ppyTxU4c4jcesNz4vx65druOWHRkFhqlXtAQnA7jyoeOOZBg4w9v90FlAeZaadplSTn6sEath
k2V4xH71UTZJ5ViN4OW/dCdOfjQ0ji07iBLEpU4q58CqHwDPB+YteYgfMs+Is1Td1We2aqHGmUQQ
eLtDBsCzWfDdPGETp/R4vsCfwWEbAiPWpjmqAh0PlErdKK5vjrmi4mgwsfOcllhMKkSJ9SLbuKsv
2PjcVxS61l9RucK1lTVHVCfv1OzAFl+TwuG+QzskZsnDJdNYKzgTqe9OX9ncDRhkjhpVm+lo5y2L
v1jt1lPQJhuG/H0njCs7vNBRUVjUYNBTStHS3BOlUJ0w8X7U3y54YVHNuySAsC0aM3J10C0Vemb3
sMl6XHocBj/CKuhvRxRy+Au66InTAijGYOtUL+xXg6AmrILVE0J+43u5iMFkuItZqMQFiRKU9lfI
C8p0TSola+Rx715LcWI+nmgcfoj7Zli6YkYzZb/8GhwpBkacbgZQriN7qntvwYhqcofAEftkQ1Vl
MNSfove6GZRrJCIaarGcGP4O3Mx0upPktz77kVyYzBzBSXwC7uijarmMJxCGstfgPtXGqysqJSLq
wI5ic/2f6oBVx1dOIxZ2YYj32+MPNtcLyFfBxYhcqzDRB1L99wT72WclMw8fQ0x9dKm5caZGTPUH
/FClLyU73r8us0pK4DrJ+pcp29KgADiTo5zDYnl5FjYJWm+D6do8plFlqCy2wElIrGL0iYSAIV+1
A8si+aKzOGuuvtlVynFQpOMXOqpH/TXBzGzi63lZCDqhoSwy9gAQWZtv0m8OmiR7I0Qdp6xWDbsm
dCQ5EHKcvfGAilo/mTMZ4hWqpp0W4yG1ei40NDFEHoC2zFvY38R0ilS1RvHVzygq6GnLv44ptfdG
mMVPTm6zCk0Hrhf2al240UGI7E9yOk5ngJKcxa/ZzyaG05UsztgyX0TIOJtKKUWN56WMlXHcNq7h
w0k/ihI+Vw5Rasl+d3AqOsJLniDj6VbZAdsHJlxszHUfbPz39K9DUTtAIdeto3uJNYDDBk9EDwMy
+Q0DBiSBdpjVsmJSKVicgXlL99mXRhRIVORWOyT3nou7Y8UYbJEKcYhiUdfco5sKveBuDLpShlMO
G63CPpetTqah+pafhTnIrSf90kyl4nQi9FvPz/aZneLyLrKeo0wtFwO1oikP4HoGFB7oYO7jmidh
LQLrNa3AOXi6KrPtNM0u28OFdB3wR+0+1d5T36WW7PRVrRHMCMhB/aHZno7MO3wBdRVd5HIwR/au
V/u2QiQcHBhcjJm548Z0wLAAC+G22kMPmDQIv34iv2ekboU4RLdCSgeCWlak5VfIQhju119Fau+N
q4ncKAh5QqHNTg5YQC89Rg9aZ6kPMSHqxFNd6XZ7siBFsfVCZubFuhWyyMcGd0L46dGK9flPy7e3
HpXAx3f2fx3U01nA/VbU+cY9zBXPrfo7Dbbi+nOLUpoVWYNk1o8O965oQeJNpNNKnFR7Xvs4h5/K
xYVjq8MUxB1+EPdvAnd+4g7pXYzE1hA0ryiWGBk3HXCc54FjtPW1gIS/nCZ7wtRc3XwBv4vdXUu+
AWXHqYsMh5T/0y59ItfdYdDo8hqtjKXPzfwRHR5Kw27zZpnjHP43hmD7mrMU2L7wnw0pRJcR8Ooc
dFBKeowKlaL/1e6iVKoFVRbdIyEKhlh5jAHNZq1pD2cQebOo1kNl6Vruk+eM0mCRIuVW8hNps+gR
S8+mUhfOXRmXoZGsdzISMhvWVjUBw9qY5dVyhjQPqR8aGZ19rs8WOV4Gi5DU26V20DTHelEaFNh3
Y8DLQCFiNtBJRc4hHtxBMa7386oPi1kMKNPiHrErJQ8PjTJPK9Q6JEWWjaKNRfFQWJdDb2LbA0RT
8h4qkZ2OiCJGrPHwe68CZ99tGq1We3DvloI0zc8GrwV9dPuB1u6jL6eLS90FfzlDFT6FgvoeF+sf
lhBwFR/jJ8jJ8qYbr1o8U/wEPTQQ9b2Pgn1gj6NUsX2sy+yniFGKiUk1ccp1TjUBoKyblvJ2JVZW
aOFBP4PjvNjxGfyXDJkXYSq8p4H3cm2eMJOghyjYox9GbbBEjYbwoLRxBOB3UG9woRYvY0MV4blt
R3o6pF5BjcPK2vVnfLEA4dG5i65jfz1AxkH4v414B7Mwr1aLPHqe0K0+zJDgos6pgUA8edFrjFj/
Acnk+PEdreR8ISh5m5qWkQmjEN7ibBB8+VVn7pzahSoo1hiOwVk0i4pRF+GQ6gnfNppif3nMXVWF
6AYDxp9FA2B1G6C0R8+Qm9H5aqY1fgSOchrUsFZuzBj1F3S0/zYIVybMyQwUDknBYHHnAnpD3gg8
YCINlNgNp+HPloYIqxT7iBHpHkcM2n8eJ3MvcZ22WSHgatH0Dw34iRZ41XMbbYwNVC948oYv3mUB
+rfqiCtaPFKYHMTOdF16LlKegGJojNrETWX1s7tBcqoYo+8fJrowzCo9ozgafmYgGbnh9FnqXQSK
c8wAKbR+Z0ArbigVGdbbxWTwM4ruHFBBGRrQptWgYIoyzNnna5HUtnVsFgw6VG1pCG+NJxFgz6DR
M2onFWJck69/xilh8d309VbEVexLbOzdyp6FPtx9GcZC2h8yTz7/dBrM+5mWjR0Vg+3PaIGTAH4T
O4JQDQ9z/hfcKqHUeAv7jMKTMnX+lKopZ2KYTn7O7iLoltwUL83nY6OLMRcKvUDYJdl7uooLoj93
RGDIT9rdYAb6F787coMdryVIIkf/l66yoccxFCZgZaWO0YwayL8yoTjBNsMFhsfXiDUT6J/nM2vC
uj2Z7Kb0p0fSKJTv7Z0LJXF373QB2RtnXCbZefle80T8dti1vZtpITcDLBxrbHVn3HiPqpPfEOtR
aaOkJAbSf7CkhWh5SySlVA1ZvJ/FjKYUKY51XHXh40+bQ66mVj1HAZxCRhMDOU7xRsqoTrawIhUL
2AV7f7//7Dmcm7e6selVzjELjDp5aOGPsJnVhXwBMSeN5wXfpJkebkcrXfv6ZISRUUJBDyGpiuuW
wkSTA7Bp2BaTRkJOK+anpn/AeM5UeDOJQWYyQQGxczAiJV5iu2jKPF2T2fsSoJd8WvCUXW29C0FX
UqjGlOy8ngQ1mA01H8LyzV4LVSrYPYmTITAljYZecql09A18HHfkqYv3bjbsqhnTYnOKri+wtrbQ
ZpVPf1g/UdR1m+sRRYWl62GYTfKw5Ata5y0UHpVO3BytkL8+FM05xH1JEXkVBsGXoG+qz4sy/Ugw
u/qNftvF0qDeeDPXI+OmNR/Z3w1UpBFNzP3hJSSLd2vSPso5Fxw2bSF6DmcubxxUo7PA8slfqUBA
FQcCCy2MVD7Et18X91jspX0Jet854ZohGt4pgTBayjGLJvRVP20rr5qZ2DTmyV2CQ802u3pzZApE
j1Yo0WzuPNU2ARfbB4qA0nBr6f0iC8OWlCfstxKFtrJvhX/IHkXruL40NPF3DcHopc7eHKfBbGE3
DUmweKjhJhoYgy0BCU4gJGBoqs4oVGavEc7IE/SXbPZ1vBZhPeDsCuuYikq+lr3TQh1KzYXImF/i
dBTeB9MV0Le83/9G4Veu6+00Oh27gu0sL4FWAaDAFjKJP1UzIdOx8uXcCIr7xu7JEvAsCYJYvZTP
OxP0MisWB7Ge04Raga3yyXLlPpChAzeR+LYx3FcT8wmJi6x2qDVoQk/epxKCKDMgrq5t/vXwEKlT
2X/9xVdp7bYotnMDe23SKvWQgqHIGhJ0ckrZt14bBV8jB2DZoyrko0qkrgVW7jbxvgFX//Ot5y5E
9eUEWGTCgzuDewxiCgirYsnamO9bWfKo4aHxUNkW6q4y2cNyQ8xIZHFty/F0geRj6Rp6XcpHfqzb
ju34htfZXsZsdekFcDuoVGgVBZgzkgt2fd2eICTvd4CiGLiIyp8lXkTXTJDlN0YDQtRnujMBWn0c
Vs3LqOqpPfCKVrHkvq8FotfC1b2r08AxPcoPE1p7LPnV+/gjT3mV+CLjc7UrR486NjkFY1I17sUv
E2+n/GFGQPfhbt3PTqP8TGWmVOePlWwJ5l1HTyHMHm0/+lANzuvL+9dm4qUBueR8BJFEmbemzbva
Qvl89FU9dHbIlIHpMiaLPnebQOlgbmSuRBhv6e78eH4HBZkCWMxHE4sQ1/2WYyS4JvdxHtxbBMeE
3O1XU6stzTKbA2+zIuSK9UbljoIWV8e/PzJYZDnoB4SazBwl6qmqOXhz0GBR+Bk9twrVWT7NqpcX
Rru0h+gYn4IvB3yiFKov4hF82oG305ur6QJpTsO5dInpY65dCil9f1ETo20kaO0rsynilE6nhVkY
26jmyq5Oixi0i3ofWgGZB9Tiq8FMATYvMhJJKkRvCn/mSwGneUTzHd4gHhxK3vyprb0NzVY/38/9
XqheRktzVy9TT3DvTBVWGNXflcq8NiEN55zIe/dEZ55GwNGykJ5+mSWo+cS2dfz5tMuX1bBnvJ3j
WeGllcXsmN7x9m/Yh0ixcRS6Ugt0lzQgBqoxOTgkBNJBtxqeIxBot01806ym83m8VF9LPQF/ybJn
wy/H/909S42OJb8E119ZUIVEVvmEKr8Y5EK/GaqWbZpkfbrAEIj+yAKFT+Z0TPaqtSdmj51gnDHQ
90oEo/Hau+udCogX73y0iXwOskxvzrtokCCn1jyJuqmWVp5Scn1CJc9FARPO9DkvEBwfiz5Irk2L
pHhqsH/SOqFweV2L3fq/FWj21V1JihZe1Ar97G+wrfHeYVWW2mwcH4vm3XRISOEOfm+mR+R0Tjvb
xikHkro8PSdiE6d2WuOPeaVs0APCYYPOxKshx18Xo0x45tAgh6PvHbznSDgEP6BGTVxUqt+KjT5J
waESoHdtSQirMmI0YKB9E9nJI7j8OiXXcTWbGqJCm/i0eSZ9vSnGN7XiwMdqAXfv1mgfEScMByu2
ncyHsBGx6+jyHbT7U5+WpmwWXMwTKQF0GFjVKZozxTXsnRvCNaXVg4LtcggiiIQhVbjYgNoZ8kv8
4SmJEOQAqC54Lyj8wqWoUTrxOO47hzHcyAwJlCN6TeU5o6qrjzO5KwJvaSYoY+tAuTtW12cS10zq
DPRa5rJlmCL82MOzUhgFKUyRL2sXp82J62GXgDl0S/9y0zKQgYIbpXgu+BQlao4h2OiwpPNXF9Xy
lpo455EiC2srFA1KvWanZYt8nPrHjRCuW5MG/A/ABzfFw/np/BXegUU4vTnYpHH7bl7Xdb8iQgCn
UZd8ikphqPsrtIVOdCTedhcZH1SjNKNCb58DpAMDlWTw6C0Q87DjlkL3hqDa40tH5sy8QeWZclWX
XNGYHhUAhd8CFzHssliUDbUs3iIAdFEV0PS8UiD0bgrdNrRsOC6nVAfCyzjzW6D346fH7lDo+uvr
huKyyGvkOKcpM/ZDs8KE5eX9XGZOFhT0vFXm1N/hlnd0lClQZ9o43gA4ZZivCo9rJQnIBw1MUX4+
aEnOR3pYy+E47iI9oM6yAqSssFKq4sQX/2bO4n3z4ttlbKiOrUFcuPbtYHl3TezuV/yPo8XR5tdf
go7RsMrpv0f0zboCOLLwWIQ/KlOLsPU5HC3G5v/izhYg8roXz1uBkUZgyCu85TpQf2uyojzhE+xQ
8IitcwxPahb8b88wKTtD0Y8x57tGzi1HsA89i6p69G0uqR29AQLj/rpfIIiyXDk0QEfockmu9oj9
RKX0fAudQw2X7Y2F1SkycpfzcB5ESEflyCapwu85NEZUHPFwE3iQU3H8vrBCjhTixC0Cx8+KFzz+
PEsKRGw9HNQqjdkv05hqqlLv/dHHmBG3anbJgQve/Zx+1+MPZeN2pdtJ9h9lC32oXugDV5B5kk/P
RCQ2dVpAdcEvQLgeEru3SJSzsPstORxDvpqd6dsmqS5X+0M6++dcWBAJWnTci7e+PZurhsR+a2eq
wvNk+/K7rvlqdfNdDmI4f6Enl0U6i7BDddQdVcjjB5xrtqY361l/Yjpx0pw0ZKct+DFrjn+4pAkP
aXQC21dhPbPLKHX5R5fN8u8kbzE7ltf8V53okIa8mZ/SA+gg4BHMurgogY7BcBWzMeIUE5v/NJJ5
hfTYby9SqVo4KQM7RCGxoiOUhtWisuQjDv6/dsApudNs8DAu8ISO5rEb8uSoN39arK6C+ysnZH96
LY8gJINWucLeawFxVHTWrcAQBZZarbON5BMBVV9n2BDZzo24rAkN4LYMgw7UI9SeG7O8bb+C9M/j
kRHfDI7xkGPWDyD/tpKwaJfamoRls8d74eOUvHDPUWQvPv6yMlqzh5lZnktK7wmF4rGSpuMstpx1
2lOkrijVvYAzDU7kHyZwJEvhVC8s+s0vCtnPGpiQxGk94tQyLS7odLx+HQ/Hxhz3+1w5xwYa8mrf
yKGYP9J56ZsKEtuWt+aN7Cwjdfumd5Yj+nAQZOZHT8Yt3RFzVcsjbxGk1Vq4bEiUmv28EaPc9AuJ
kgH2S6fs+mCW59LxzhHyUJJsmJkrxTWsuMqtdL1y1pXoo11CXR86RN+eIm+ir0UE64VQG7VxwBx2
jYXSDgC+Jo3I7S3I5ioGjRqXT/Inlj+8eTrFh2DywqkgFTIzc6eYpTnsvnT9Ymn68Lal56EmI4C5
gAAyjFV5BaAybCSTKUOBv8uBai4yXqZzXXJA1efUr4DQSISSkwK1eTUDamt45KW4bSw7SvCHY1Ov
VDioeGkEOXwJ6vhzCOyYLioBQgT1U1C825MJwrXG/+ea9PEbc/esM/q359x2Fm20BX63BsRj4TJq
pRmfbw/Hj6A7aEG8j31uR/pLTW+Vbrkq4rTF2OFgxSnrCxD4g+8uxNqxuCwKIrpMxYN19omhKo+C
IXwwwNuPsj7a16Q3nlIVGZdWElmjat0037n4oUweHRJlWuuvVU/4h1jOaqujYyLR0nLloJnuiDCy
FDLMvOA3LuNY1gMfKjIGEyiU/UWpHcqfpVlnNYWKKtquCtdA8L1M0TLqgWDe6i4LVoUT6fVBzSbL
KAlTWm0jO0TaFxtc+EJiWk05BrOcDOJaIF9aAMpN+YSHh8s9WE3yf0k3hYaD6AOGyoPekqMv0sHD
TYgt+26iox7ps3fKN0JiJZQevk4fqjQCWZty+rawzvZ3mWD6lK6MHWEW2BoVfJYPilah9aSQ1gUB
OlGMfPwW+g/TVtyiP1jgTpCBTV5D96BayNOTtfSC6SHdNR+QG53yr+CMR3K3iKUFgQykHhA0bgO0
0aoYC1m9EyN2d7xlp5MbbN+PAdEWTTPpUtWQtgrM/LRju74vpEr6WwRqLjxSFroPi+euW33/jYVs
U8IK/2nZaiPLDJpOxeXUHSjaMKlXbv2tSyu2043sQznY2Yr4YSMj2gKmfjDFx63yY5O7u9BoeFvH
IWD2cIbNm+Nj6PbaXcSpNxmTFr+LL/5q0ArK4CW2/VJEOcDTmzuiBzNAZ3Y7LQ+GvJ9MZM6iuDaq
54ZLhazaDLaQM52VOPHECVLtJEFCpyxWlz85ewNmitlbt4nJNEoFPNXW1i10bENQcrlW5RRLLD4t
Op2PIbchRdN4vY5xUQm/POzDs8XsyiDohcYvtURqdPUKq8dwyh7YKSFOJypnRZQ1bJY5RpZz78Os
uwS84RHNxVCz/FjrEZKPVoUV7dwRTzsytanKIs8dl5GqLuwLYGpLYD3L7fd/woN2pRraMIgw/y9t
zO4xtVa2Mzs6FQuaOI3Bk+VKgHYaowORaq2ibwJLO13B6cdhbhqSZexMZ/y2bM9afzLjiUqgGBpl
5SUO/wP1OCwsFDVrWKmhI40ZEB4Tug9bCLR2hkEVNZ2ARxLK/6VSU5v4j6P+lmoa1rWgQKaRQlqY
zW2lsYExI7wQz+8sS8qrgHafLD1NYjwdloAAxhB+Mf5TEX4waf1uZKJ/P/QmHuICgE3pCRfL3+cI
hoyLSQeV5OMxkdkeVLc/us+jwGHKr6BbhGLnw7kf9J0Q40EZWETl7Lk102YqEz6/2yIXtRPWxjy6
H0ZhyD/gatinfDz/ZrMffxIljQrTG4WoTrS88ZAib04vosIz/9A4ZxXOtbDHg/aoaJQzz1DXTZA9
c5jHTVthf2VSbHLWGU8b1UTwoqSyYIc+S8lkdyKV2FO3+WENvaESu0PA2fD+jAFUpmEsM3axo1MP
i21+4offo3MpSElcbcHsC9/c/epHk1SKD/IaDPn4Qjco3lBJCnVNCdQyZIwett8zHhmNn5VWtXjx
sNiIUtVqrhdW++pqgOmG1zHLJqxmlRZsbsl5gl9LE/R7O1aXiAEfuIkqVTdvw4oyDWK3UMdWDjFv
k56ZIc6wFe9HhQJ1DvC6fFSGmKsH/vty4+xcNdfj8KCzbCDrCDpb89pjM20BbpD0XLmqA9elP11M
ctxYuarxbRTp8tIpyA1XBBkOYWEVwt/wS+zEHNDmVQ63OZwskRByO6/IsOATyQqf9y+dcyvPpUIO
FW0/Kc79ou67PjFPe+OlmmsuyyLQEnbQLXLP3KSua8flCZMd8KXNphNGbz1H0A39fmHewsowDHbN
H09xDqrqPn5LdmvoK1EaMJyOCUvGczfoGS/uH8I7Hs0rG1+ouiTIldZKvon1iOLmBG//ecb2/1JF
zcvhJKYVhzVB/p/zlZgnBJHGDw7SXAJfsxfU+xXqwSptvpvJqoGm6zWSq8nHFFos6h2L23bC1RFA
Su7+Zf+oQRr/XSMrvYbwzvZkwXgl2CAQEvQDQnlmcyFsUXJotGaCcSMcFc0gjrZYiudj4sMbUG7w
w5XTenoKx7CdtA/v/4VeI0N3xyo8kBOiy9vUjhENuSaa+/McvNBv13xlejXVq8JnGJ8QiM+HHfBp
68x3+Q327kTvyaHD3ZcAuhchipgT+6K0ZeAB61ia4uH56xIiTV4Wj0thhv5NHIg3SkauYYAlZ+Z9
q3XeXdsKLBFq7GKdVQC1E6ZchTWJILWOEU9vf6A9v5hq7obcXw7k+Kb6ympOSWoIfktmKTRX1fb5
cS1JeBPM6BfIP9MLEFO8Ifwi/CmDyrytxDeJH8CVVSuViQJgnITF3EA8+AGCD/fwQc9AicmUOSoq
+6U0Az/ujhp1UWN4XXiH3huzRS5+EozgnhAS8keLJUHu3soGS9TLET25U7j52zT5vBer6BLir5xv
lDd+PXFMrOBLO32JZB+SCNLlitREh6aWP7qy+ZJ/0OrncvQfynxhmbrsD1y2feKyuqoVYJKvwWEC
gSzsciStgLGTOScVtVEG87VsGbBKtdsMwko5LQcPnE+PpM51D3Jlhl1TbddVIKsRnAb63i8Lrvzq
YmlKd/AK3bDOrOU5UZdK6cKgpwo4Qieru/V3cKIxJuv9tWuloqEnLcV9sudTDA3EEd3nsApf924a
r53PWrT35h5ZcO2/466q60cd+btc6KaOA11LUNoLsdUAD+bZOjvg3vep+TVJH237Sz4Z5006kCcW
DEO1l23TBxKiIaC0fuhsRFx+sE1gNNarPV6LI5hZkLp1VAMXACtixkXGs42McC6RwrAasHVuE5w3
/RYtQSJYKXYv+6pJ6ftIGUVty62sA5LkzAyASvwsH0hzk1Lwu5CgKEtrzULbkEsYvvKYOGUOGxQU
lgMtdemuDMl5dO5nu3Kb+az8xaj70KnmxWHyDj2irpW6RfN8GPbHmitD7ZL6ebbZf+6kuW7u4qYq
vhspdUz0RvDxz92skpN6OZ3Ekmp/RV83xBK2ZDYNOtPkdHEC8hSUcN470WfA+CeYQGi6eXUI8i2C
lcTefT/W4j8p+TsOWyPmUV2L4IDycc1KNuB9gfgORZI+QnAz2tKYZBcy57fjjiue2NkFrN00pfNT
Rs1CUJdTMpjfHNInRj9rTbB+4jbL8xR4396IVO0L0pSAj3rJ+5rPjC2H4B5FlJ7JU+ac0Mv6cwMf
B2f/YS6FMHg15AvVB2WPFcThdJBaSS/s0w47nAXzdqpklqMoZHrZWK4ZJ21oG3BwtgC/M63fGarT
S0DPJP2zHoHaSZKKgLmclCEEA3yh/QCzHf7CmMG2wWIwhVQYmVzfMgVCMmf9oY1aBix1e6yj9sX2
4j7bqrYsWSZwCRFY0fH2qXzUpmTBuJet417lYJ/uClG/DeGeDmwtN+G7/g4b4LadaX7k9G4fr4YR
cGjrlN4oiqEQbv9jvpXSPXBE5Lb7ayndZSCdIcPhNh+2a1ec2fsklLQmcXlukgsLNlRVZZUBRWlt
z9c095pQ5qx1C58hTDL+bX7mQMqU89Uh2Axm6i3c/PRdEi27mOYGwMBQpvCbYcK0dBws2VA3igyi
5ib+rcXZHOfKDiMn8fvQHdQjCfOAAiG0oisfKXM8a5/C/g16vVvLOCErj0itum4kmWIm/u3sDtVb
Wm0aJ9z9nYs8rspkDDJ+qvrIxK70Wp2MC5rlaXeizk7+LuOFDCD8iSGU+k0RzeWwU2shLEnnEzrP
7ia2lnVz18OBkHnbSu3XUUUiWlJDx34azUSShZkHmZwLUu38AAGpO9eYQJtFg7p7pNSw9z+pOt45
uCzApx9Ln5zdn2+bl6phooiHznWosRF+v1hMKgJSfX0Zig5bIgMdmYptrS5pbiNKeRLCyNHcW99J
xsFS1koXxzasmlXXesR1Kg5PUA+kcl4uDsM1BPVeofdxc5BSGypEfxL1EqRyj9S4zH9M2ZKc6ON8
V8if8LJ0LrLHEZ3cCxPGMXntQCE/JYvzfb931N0ZJhtvdLWpuy7+kN5aFUBC19UiFRRRnYph22TU
qDF5+Q2gd4WyvHnG1Ttk68e9LaRh/NUAvGqPuu0mokUaYsK3VvcpCSgn/kmPFj19SliLjFYClBKZ
Tja/q+++4DGomJEienK3Glr+u2j2oI+S4d/Pq8CRx5QsmTSODJ/WFednEeTNyOtukhZnliZeop9S
Au0QfTYCP4iKpmKG19A9puWb2kWE1iwXS2GzEnhlv/3ilyn4U4MknxyR4ywXlKE2ImwQhGGWrAh3
FjxaBrCXym5I8tbC8x94FAPjasJeEupOri0/smK4SP4ANh+KBm4wwtj93JA/45tgJWQebBwZ6CME
xRQ+4AydxZle1ROqJ9oYbR76ZrVZbJIhPt+9BGFHmQYXFjaI7akA1KURCzbP+jqeGypTonTHj4yd
DSs54gQI5eXc6eEnHjsGXnlwbu2SMlZckKlg7ibh1buFVufFc9TSIiXnkuEls113BkaC1Ksb72Io
YTZFP2/oaXwJcft+J5RV76hK9D+fzPD+Vn/FV6wKfqXne/4vALDjbTEF3gRZkLQAx4uqYCsb1o7z
3FnuEsNzpESBOzrTyHvucgJtog3TTMy5c7yuk+1kNTmB2aNsurCgUXDbDzlkCVbtujDBYnry565n
/diTdMT8h8lpCzMnWFScrPokjgtRBGOuLPO6t9TrEGUrX/MEuIg9I2aZsSj3JtXfQHRRX+1SJtGD
EdHT6miYszN9frvMNDBdpUvVrMYHyRWAyDqZMutSxgMm3sYZZrsOVFRPOSsmjuMbphNNqFdldIh0
/ooT4QbBned1sW89/K66cbkrWd7rTz2R/VWuCYIEPcZLR5ol92VnlVIG598IRpDGdLnTqxU243Bw
klNZJC3h3DfXYkHeGBmz2WeuKdOp9G78154JLvpypqamaGKsnS6J5xxOWIDJOhqtZmRQrNUajbJ7
y8RoGldkIfPi1lzfkZkCW2oeHi+fL8wpQaA8J8fTgZgwlLLP0TNbJiPhQhpeDb1D8VudZTTSCDWd
sshmlaIpB4NIuasT0ikj1sbno6AUs2VAUDJ2kDzuFEel5efFWkSl9ZV2t5HVT3lwU/BGBbgFK7jE
cIH6jwSqqESlRmHz3tNI4GTEfPlsrKMQQjxYglpGy5XfgU6p50VBnT4Zq5qjzBrCrlLQ84Aa20UI
3V8nid9wCFqI7YwLM1LKvBwD5KMxFw3I1zokdM8Gyq8bB7duxV6usX9MvxIeWEsLyxaHvbMInnW1
eUeccLT8laH8z6jsZLD6ynoerP0ZIbVoIl68QOQvskrlnpDn6NxPFuWMA4gos+Fj10cmraGOHvu8
cz1K7DF7+5zoqN9CFWw5u3TnH8hweeD4PanLQgjiT40f3ALPronCUl2Aiu6RN1rewX8yksbYUf0a
XYxSOqPIBTnuurCdhRU4mOfnYQTb59UNjYA3OkeqrRb132l/HQuKmPZ7vB4dmBPd4BIVJUMiyZkc
5jj6VCe4AKQNqKO2y/gx0r4UZqTWZ7m+rJ87PxzIw42EdEKAE57A1t32WO9csoMxRXCnER5ysKNp
SmYPkMVRoiYLLmAYqkkKL+btc+nddh73InhFc83x6p/koNMMd4JqCuwfKJm2KC0/KECSkkqo5x0Y
dsVfdPoRpnQ33byhNBlGsdys30e2AsDiy4adaTrdQ0Ebc/fKs4lAJ4DuOdXNeJwmQfNQeia0WZCS
k7Tgw9874HHe73SUpZTeSJFkCGW18sG7TEQEd6s2AjWk3ktnwejfdRp29vRB2hq0Kv+ZpvArX0jm
mN6GY2iFsY7pe2NQ0lhYolD1usK0DXvf17uIEf+I2A81Z7cwIagmhISh5Vgbm/lG2bvybI6yZzTl
mCVqkPUZXJqFZ1gCbSendBQ54TqKWfmyffn0g3/HnE4oZy2mQG5HDAvznKAaL2pbVnxnKDv/s7e/
FgIfCGRjgV888P0iAtas4qELT5C/gkuOtpFrzNpLeB9XbyzU+8OeNZul+o2tFFb/bKLqOnmVmXED
RvwL41wUgoG05gTiiGytwFrgR5LJX1meRnFt6XCcXQBUtpEpeg51n3W4sh6lJcgtl0Hn3Uw7/fCE
C2CPjRWVPcn/xlMCy3by1RS7o0n/q8tqAG1ujGu64aNgpt7jddiAnP1Y01IfKwU3ReJ5Ty9SnN1L
I5nyLjmZEbf+lajjBF/852e6JgNlqJmkxWQvs2lSszbcUbA8x3+TWbEIk09sZ3pF/VmPPCj07sho
+IfIaIWHgtbyHIbS/Yzq6y+KBsatGhNwP6TKSmEeHGAO6C2A7dCciE4CnVOybu+Z0St5vKkoyN2D
8BkBRhwtP5NJX1JsJW0Q53X/j8aPvW7O6bf+66m6VqZ7wIMadA/UzJ6Crg4FyFTcQ1O5Sx+NyUjt
gXM+HUDfVK41iXNrx0EGVUNdKsiPNzj88jt7O9U0muXq83LCdHuYH7mXrUToh1GhCWU4B5uHg3YI
oCV/MaBNKVH7hPGIKxKa8o51Exn7d1vxrIs0a/+cwY/pZAEI64I+J/Njl1+8cqmQJqqu55CFcM0v
DD/FXv1d7xt9ZoyrSb9heyt0jBw0xypMn14qU0drWx2b5KTNamndAjwv97MZJQFzGgoniy5fd7HE
6ewW28JjmhAfEArs/ZzBq5tseIjKg6Q/DyIuIHQl3ERrPL/xC9X2cyLWZzARqBZpHDz7bUQ+24uD
EX1UduREsr985IYAEM5i7bt+njxRcw2TbKADpJgFj5nJiflhIrWVzSILzShBfdGE4q66aslq9v+U
6XDAEG7yLYPMMYL4fpp6DwK9OLRN06OKL15gCBmaPS974WbZWbJF8ZQilaNkU+8QBhOJ5mL0a44p
f0d8lHaQ/QVhaBSJ3Aie5k6eqMkeG5uwk3wODUsPnyRmBgnw5g/RMlEySkUlNVmRqQwCNCgtwWWr
AaCtQjTkyIDZ0QCviMuDDiXrjkxCw2xGZWDL+cJBvcwf2eJ8eYkpnbeahsaxh06euBeUVflF5nTN
kW8sPVPTda9Rt6b7+i2XnwId02PcnkAH6z+Erp26Zmbb+5de+turg7YRJ95r3vaN6biQR3A5j7CI
o5XsLfZPcO9KCQa8DS/2A9Rc2t5wwEsS2iR0ouFGIdnwqbHMxmXyDoO5GmZu2MPnZJXcqcFKxdg3
PK4nXR/6TUL167ypWeBXWVCFInr87f4h+hGoBMaMvXKK78hVRS1twbaqRtnyVj2xFXv/iuSGJKNw
EAjlDR6JdTMnktHUAhl/NTbH6jtkHUj3gD8Gfs0uLNTQj5vG1gZVSaOYECian2DE4dLuoJvT0wKp
OLEwm6kGutwQpTf19j9DE6U3PmjJ27y0zUO4nN6Xt+416zU8hu9/JfabS2ZvKXEnV33AYl1Jyxi1
I/iGS/QTSl9dw2SFmBuJ7ydHJmPrwZ2obGg6PW+UTR5VLF66r3IybwoYMIcZfk489zFCBgJpieyj
eYoNCaytcnFMikMxTZLUvfKig8PH1D9hWuxtT1BM0nBsoRa1rm9jvvP5NeixOg3888WyJEv2Oo2k
GF9M0I5yJ5JO83KHeOy1lgtzrb9rMpeWRdCX6q2xH8epQ5d11nwnwSDf9oxXR7UjNYz58LQ8sfDL
rnMc+Kt7fbkP8662jahz6R2K+nMXUYmKuTF8Io5qQXBnocpqrAGkOv4tQoBKkF1oI04e0gMYJdNV
WtHA3s09feCY9ikVJJdre4JMEjUCDOPkknJsiDSsbUf/2QWpjw+TrGkCRAbYyUuiW8Jbvtn03EtG
crNr4Zd+K5Isefkf0GZdyzBLgVCUnWrYOoWNHnaSa7IQrd7zykkxTZSkv27ezPtFXaPM6XZTM3wG
6KVgTtyaF7Oaj/uITroeDj5HQs52CQ//s+GBBafek2uH8YeLUGpdh28okGDec/ScpmWyTEUoPCty
ajt948h/0u0mJPgUEcGkd/0klwSSfpXjUa+64uymYT1sQsy8L8YLYktTou7A/fiOxO+NMgsbidZU
kvPxIachlEm/vmoULufNFZVzbBUxf0L9TvQlRNjNN1DRliZKYZOa+JhbEvjMN5H2Z0CMQzfFjsZn
eysnEOPO/B21HqrsB6IOWX0IQ3derFZGMa7lNgM+pYC54FHqf13F2qiPszrqYQthTkC92eq9OKA9
SpiT2bWbJCn+TJr5D9VMqF+XJBnB/C0SoiGgM5OTDnBuEXt+Zj7XjbQf+o8oJp4Ve6yNzBL7Rfhq
zu+xCwyah+kfJgnNd4oNTVzoQkdkgOiZlKxuPDzcC2KTC2kIxz0iSzg9m+TfTKGrHHEz3tMprFKF
ynOMhDWwnFMT8HdokIjab2kEuWPdUY2r5A2QtrHrv34IXu5CJL/G6fWStjt7kWWaWQsu/oyXm53n
OjLV4e1A7nUR19MmcZlB1v0YiVeP8qFOSZXDNaq00qerBRJsPMk01wQQtfMILfH+PRwYn5bJh9Gf
P93tzsWSrdEgrBscHaDtu9nQKIDM2de8zPGNWSxGsYGI2lTAiusm8DDbtvmA980K7fH/8iNsV///
pGYvTf7SlLiAB44JU6Ly2/jY8NEngbWfN1RnLKHd9z/SJ0w6fTKO6FKp2bRcrJxJWcZzui9hLIAG
szcK2S62IgB5GyD/xpbwtBPxQZDDowJLJp7hhs8Dkf26T81HYVyuVDsgmzzTjQuJQHgYIRdfvARG
uAfC1FIV4O4s8tJKzhj8GxDjQ8axU8whpZ8kvFG/HhV1QWWH+pUXXRYc0vE/nktj6BqMlxI4xjnO
vI9wrcd6XrgK0hJTDJchjfmltR5beewpcTUtjJn7CCSGR3pVTSwkOD1XYuo/SLJMRau2B/bZeVU8
+MmT7h6bvYtHVF93SeoX+2Bx81XUs5ZVYVLf8b/6iWOlXVCBsHeb5Rl/aO8ouzmuqpvp0SjKqfNy
P0jhbdmRLPwwFG2DRg3Ygse7Zg0GvwznX6xwHj/uD4jvcEnaVTnpjLvHu8SPlo/Ss0a1j2PQ81HX
BU27HHhom7LZnbvImMZGJRlgnJlAZ1BdaANfsOQYnWvR4wLUAL4P9i1Rqc9eqbQmp4NlHHW1nDrs
dhDDl80v4z9HsjZYf28nU4Q9FQSxpj0uUldIsoKSj4QtFJsHU///pHfAgXpGEP5spuRfjuG8loTO
uqu/wOKMFVUDJMm3xYnGS6Ao6mK76eGzBHDhAf1FSgg1Khe3g8H6ePKfrTLZwC13xLAiI7riYGdO
ONFrcJXLW/YRxOLLu1NBp6ievGSoFg/ZASCrRxyqqK0Ga1L0dUkCJn+5ZwvAfuuaNrBo+/kq/d0j
wTHl+zspZiqGbP9RWR/oV6cHavz2E2D6F0sXTsEs0MQmneNgvxb4vmdwHXi6hgPhg2ISZDytLIuJ
wUAj3FK7L+fAhhEf4MrwdNU89GnGfFbxU8RetcCm87nkeoDgnoDv6B23KPF6qAtOHZbfCdkuZAu/
iLiKTBjR28YUITe7NHgzr9U+0aw/H9Qjwflt1Um2v0GDtCbb7/8PqgGnnOC7OePI784TfUU9BR9B
IN0ca9B0B7sdcAOeYiW49Ap2QSXxY0OPfTKzDb7/8OUmpjY09pODG54NjRje7rsFHL/NHYj2Izy4
9qKV305Rer/8s90iZF2bTCg5qdvYEQGoEYWCrd5XoMc85P8PdhQMm8EPGILDLMdFM7ZF8JJgHk40
LhXG/Vn6WB4s6RdOwb2B/0ZetNmt9uNhsDReE86/S2Uwclu7Tgr+ciuJ/JM6s/Qp6+Oxn92ihyhg
xll0EzbY/1VBsLaguqabPTPcxP4j6AtHeYKOj2eQFUtxeTGREin1z5Eol9f19WnzdsJ5R3V4yx7r
8IMwHJG6RyvyBv0HPM8203MlccYQZH7PrhCsZv3ytd6BGlRb7ni2ep139CZG2N91RKcGP09Z138Y
sgHUQx7u9oFAEKSNVxkI+bqe84MnPFFTaKhYYaXyqW87ncxyJFZus2aaAhJmZEXrxlrcmFDZFnaw
TA3p+VoM234BwtnZvaJp/iVCNOLKxXlwS3TCWKPHwytO56NaVKguaL+N/qOGjKrXfOngx6CsMbmb
ALtiQDAkaWnu9+HMCEoUMHPyT/Cxrulmte7Xu5A9ToOpEsK1UNNkkIMpvZzXuNaknhRtDL1PPl8S
MgJAzCJvSPz+wljbrj2+Xhf5rruFU/s5LjRRh3Icx8ILVtv/uac3M4lHwqTGwpc4xcF0ZNQMzTqD
VttNFkvumhyP8KBZvyJmAqjfLDlfbuUVija1FOoI/v0joFDf/qdP/8g69aPR9kyCosYwfwU8w21T
QsUHnKSd8nU6PuRgqvtDyu9A3mNxpn/fuZkR5Mwvlh/vwVpi3V1O9viHZxuBt0vdd+LpL2cYBCer
Nzme+YE2WDMhimJh5OOULlD5O5kkbvdstu1HXKjwuNKXPdrLtd7H2XFWRJseOXVhUlEj0Ds+6SVx
Oz9rQRRm+TKasT5QM0Y7NJbQsngy6v3RYa9mC35L3g1taS3L6+sRG0+fcwIF1yWjK+JbNlmuNIoH
j4giVycxZoZRZih/rz37AiqlRrCyDBQMGzhvxVa6r4qSDXyhqm22I3T5p3Ka06geGAPhYqt6a6dD
EQn2RVvuUKGmAsTBu2qb6aAyinZnCHrh3L9fxyELcYEUiswm1dPqXb8J/Ro7w/rNnXmEFi28fwic
tckmnkwNTwpblx67l9foWfwDRGXksibcTH9NEH+526zH6RyRYyCk+gnyED2W4N/9BIeejUgs7o7f
wVhu5Eg3JCUrLVhUSG1jbBCT1JXlMVQ52+Ilc9Xn883WYHZ8KWSVfozgPqyJufvqyXtw8m8DoW2c
jNxRsMQsA9GMk6UgZ0qTV0M/XPMIh7grLeU2B0ywZnad3xSDGEK5ribURMZQ9EoWXXomfFvKVTVs
fqUAYxZXXbCt+67+OVDmTrF24Uekonf/4nzyYkoXlnX5GeaVzoVkSLqbeilU6k9kvuuCylG1iHPT
QGHl3hRAFDVSb9NF9TFknx5AIIbEssz15XgdY14z34SoVV9q67+F7wLMeEE9zzZE9wV6ihn8HmdF
Cy/rslMSjTmkL6kWW1/9f0D5GhXmfz0ukGVl3/O4bi4jVJ4UqW4afb2D0sw/SrtXQLGVtvZS1QtC
Fj/tmBnX5ShPPdRdbEA9bOtUP8DygrjkaFmE2+atAHEELDE+CtrzRfTpvSWMYFX7pPGCwoxctdSX
gGaMvXXXP5uOVUoz09E3kxWd96770+Au6pRAHAKU3dPLfCq875OH/DPoeom1U/LEXlodqFr/j0q1
YF/MHTQVYorambYrNTgtvmSG2EXOgC9lwxeE2GEBgGRsWjsoWMT2UE5Ux8v9hqxU6KhS902zsiyQ
xvTaM2bXHOsSPoQzssLjwBgf9bHyd3IIjRUhHu5kx+BObkzuq7AqY1SnN+ZqmZWn2+NgO+YhzSE2
Kj4FuyOW2wnUZCnTbyvUKRKg/VlUb7Yx84uWYnzJ8XYy5QPHNzncpBJQF82nhw/iSSZ5zcMBIeRg
BNNEMJgZoJs94Y55v5iHkfDpiQS4n7AvLoEtgB0VHz1iL5O3avv5BIBeUXnxC6HpfVkLroMZhFEQ
I39CDDkKetCr+QUplmdjtfS/bWSFVqBBrtC7au40GOKS8QOPUiB+AXGeLsDF+RTkb7EAmIc9zFos
ufMnED5cTL7JA9xZfM8WlzbUi1W2BKZueCqwgXe1z416jLhNtmQ9nVuZV3IDxiqYQJZkbnhGa6rM
sdL+a0NoCAkFTplS7bO9S8kx00/HzVNQXACf16TA9PlnUvltBOUyw+QguEhQ2oNNj112ufCVfddv
sGCtwG1gJLS35opqGvs+GfmjBdObAorH8pgB3GIknW8WIfvTq0VmMPBYpj8nFtcDhCwbxLeR1xRt
BOWH9J/gKj5GLwM3gt7QC9L0gNsp7DdyMaipdnJG3KIQShR9bmJ6M46RnbzFy4Q3UOssLgGaEfhG
GwWGEgu8B99wlsDPBHtg7RHi7ILMeje7Wo6ndXRYbVldTgcSLpsV5TUvfUWhdekubBPwW8ewbaLF
jlMoCo+Fq4uALHTgci93bOlxn9vNNS006KwbBmMK3DIl42GLP3N6yglJNpvf2fd7KCJuw7kkCjCL
trf+cfxLwfcRyHeB6+JfpBwRgDnAIAQeq73yxrGbpl5s/t3eyGr9SoKzHdhJuMb1YwKvmOsg+0OX
l4tyWsv2eEfo5hfTmlj2EZxHfAbIEPVE+oNbSUxR52/tIaM15ELG87I1pGWuJQh3fzY2vqCHlly9
CSEVvcrYhPrMcJVetfTkNnr/EHP2ZTZ4L+RrLT7N1h3xVYNyLvLMR3tVATRbKNvdFJqfAGlMLcm1
zbewjeObJSu71vuLJd5XWYZtSpdu1pamH5A2Gk5SmHoqigj0xExKvLPPCgaCXBGS5zkTtAkpcm2Z
taXctKmLxeQOPyZgbd8mQ7/098H4LdVU2tdUSLY7VHX42f8mVE3kqwcIeOA35JRsXxvEwFLLL3Zz
P2d+ndZnkk8Y7v0gAW3p9iXNtbShVxxt+//ujCw1k3mFml3cVWJow/gGxjbtQuiNvISpASpzcATo
g5Xu6wR+Q6TodL9EOcmQM+0Uct/MKroyqBXbk86n3xk059nk08YV54kQny/xHaNCf6RkkIAwdt0J
OQW+DbTEDxLJEo+LS7holwwqPw9KDE7M7U0j4hMaqvDWLO11Pl4hIFcugYgC7Q+zupoHDP8ySFQ+
cGmWtFFiueBGoek3PKdrkdGpIsLwH6lVesBShVChFoB55cRrzsT5RjGrybvcvnFu1wwTLcvy0Zfu
q1sRMNc66GS0G1npyizFFATuvZ/vQXBKZVYtG42/FYHhOsw0AE02ibB9Cq8h8Zmm6Maft0OnVvYz
kHtwsZa9V8EvYiv9EF0oLdXAGJkwB8LBnReD1rgVrppzdRingdTsNuhA77D3W8eUo44Vob4c9ME4
A1uRymyqlYLmLJQQZnqcthTIlhPBHPzKu2W1Xp4oIeQwCSPXdS/D0kFI3zbcMe6SbMEUYKW8e3FB
c+ppSDONb+ogijY9lO8ocAVhfGfIA4LlNXnx/f6EsFSFfcb6eozRPM1v9oISBnE17MGuSrJk0MZx
xM0PBU4cv/Ufas8iAav2TAC8/i6S5B9pffZ32QJxWJmh8ncHE6We1+7ItSojTeNDXKIVnjyrn62O
hScxVZxrNdokWm1OZUJQDrgrdmV2dEeAeWXlkYqSmddts5M/uLEXC07kv03AzkGaGlLdBk43I91n
xCae9F19It3oBYOHcqFfmG/tuQrZdtJkFdbiAdSciIhxJFviTPuEnF1ZgFcMfgNQQPuPYfED4FIg
K+r3ho1+fboJYVSlcZwWF7cxQGt2YNEXq0vRoD1F9WhsVPpIaTgyFSghegfNB4VC8UIHZtLMJVai
lbvTdg3xyMxnUgODGo/xPMumKjgz7wCRzVwkpvGU0YHt6L760d6/LavtxWBtxJyWKkMpIiWnII9u
r1sH2deMcHwEOwDLVIv3HyMvl3982B2idA7/DyXXXaA3Aw7WdevaQrIcWLmKhH4053Uu4lHiEnO6
ndv1i2Y7DfGaWxcUJKZFMpSpm3Z1XlUyWYovz7B8tDBCZvHWeAMjrP4upLjPxHt+MUndH24I1WBs
Mmu6aguUMd24FmrIPLrrr/GKwjfSHQGzy24WiaK90wYcy3tqWfcs36pD50TM/x/Ug7v/sP4XX32o
fn4W+KRhM2QmBg8rGNqhsUMhK/LM8Q82tqoa3WkDGG+/7GBBSEs9cyA28bEjTkOvQWYLyHcrf7e6
iXjvwOhZe4rC6rXql2EnJMw8wWXLfVb9Jto1i5Qtx5wI4bID2TxTnDniy68U6tXRqL5afLlKRXq9
lil91Bm2VM/W31ZikV+NyqeIa2CVely2dfztM9ngHEKVa24yhBOgdK5nHLbIDv260DPpucIUt9hz
VqjZHR0SA4ahZGJWKkj+q8snDpkqV+jRCQBbO2D+Aho3Bq6pwnWdwaTwSYQ0q1VIt8qBFO3T91kU
40uVo0fr8lrdOWKMcRfc2Bh1OWltT/MFdTJS9n6SXAT4q/2mJX3wPPavpSzplcuL+0tzzQwttRxj
BDasNI8cwrct2EUh87mjO+bphyitwz7sHVgBgEVcINxfT+u5l4XN66s9kxetv7cVChjbGAsu8/lK
SNQ7NtNKjhUB/Of9KOSRQNpESAVoDG7EwHY6FMvCvUeVbzzR8ECfeIBkYEiMj2pOS57Gbnugk168
EpYBAJTaOaZ4XTRQylcF6cAxCNENXY+5tL3/iAgB91lD5U3WBYMSe1wEu7PXanfzg/FrTUcvGqoh
VtCQda1BH/RlW6x95PhKDvRt8dfkJ15Sj/NFO3wL9SkZP1lDE40UdMBa7heP3JurhU9inBCRLKgQ
oQRSobHq+HRQzLDWLF8D8/ir/CzYgSYfsdnNBjp3v3d0OfMu/hqKW3fSkkjjG1vE5DT7VXIjmmUa
sXIB2R54LAf+9ozLuiQtkG7aS6+y/mfGPHH+KRsmLj+5aypA4rQG6g03hG+V5qEjdoM//DZ8CdQt
y9FPsqSGSTPcNBgNpQLiVGiWw/aglUrCEQS1h1My+X0AEiRyw6cCTiY2YMKVoy+4dPMcZsTzvWJf
qE5fREX0ojGdRnJxKF9deMMiCRzvYGayEE5w73sykdidPa6/TxuJ7Ges3ZCxy7AjzgZCKXVwoLKL
z59y5OawpuswxMOd8nuSq+BgtANp7cC0zBf75lqDdKBFakcnO3PEtwCljjHeZhDeqZ8U1y5CfH1F
aayFsyAekhOv5xhu+bnLMB9mAjAVkOatstxCZAVgknNzt4vmnCDd4UT9hiOEbjzraC+Jwv8mMYhY
1gCzjjWjBHasNmC+m0A3KHs/3p4EEg2szZ7+9lxxAhW00UHGgEknYyytXSsmYvsOWTGMyGJl2I2T
+eqbY1aaGi04kDwRMuXVI4WZvHA0kxDtU66CLxq5MpB6UStYcCnk+leCdA6L9SpeACKeVy2qzNfl
iOCEswVx4SBhXbpNioVzaD19/NiB6ZHCP6zMUgla5FqLGthq/LYO4kMCN75Y/UY+iBnC3V6Pk1m6
oo0SthL09SqEYp0QBsBO8glJXLyk7VB54Yfotf43bfVbbuqoAoLOPieztfRkQg8sRO2ZlgqelYkE
oWCtp9cefQdHuc3Y1nmN0oJh7p8ahIhW93Y9lxruiVT8uR5a/JgC+ySqyAI4tJ3IpltdSkpkMcP9
31o60jfJ+Bk98n97ywPj2w2ZKz/TFnxVKjPOQNhWLwYUTJ9tnNzGEfGgU5zDHbSuMFRWyD0OPZQx
6dSQDiNeE+rSi0WBecst9i7GlMZvzYxZDcUwUebmE1eEwnXLCKBY3A+OXFCcMFMz6tq9HAzPZU/V
SVjWiLpGBi0gSpFzXcTPjoZa+NKnc5kdGq6QLPiKcD+j/VOkzm+LSUNTc77wo2wj5XVDfQ9GU4m4
nO6fce+wMibIokuDcZcxixHGazq9wsNwty7W9gQBJbSHYO31KP1wWjoxdes9G7Dhve4GOAZrcRY0
rPLVvPm6pKLR+l9OEEFGYYZgVgCraY7qQbfD/TqY7YtpFTJJxcisquaCkqPvpzaXKLetoeOnjOWo
fMX0G4BiqdNaKDyUXp9DYGcW3hyifOPtMThEcLk2dvi2lDpjvnyDsGW2P9wnSdHQ67O0mVa4tDWX
ILUKCk9O/aECHfTnC02dao8FBggKrJyb4DdWJVfdxZwm3YZxWY5Wlq85iMLvV46LCfBmTkW5tzO6
WRJrv0gNNjiuKYMJNSCxtELD7tD4UT5udoGmGGAjqK33WmA/6dZCAbEdMhs0uUngufQZcxEGH/xn
oABBvixDHPzJne5eN4avNCU+T+b+fAVkdZ+NvxWdkmlrBOzU74I5aSPrmXX1ocgmE4EEEaccvBSg
UyxDQ4BCN6LEQvKTTi182P0r8HZXaa8ahDtHZ6yrC2ABRL5jD1I5Svs8z8XQMh5o383eKl189uuN
Nx3hsMsgyXtkGLy8MEnzm3V4X4nYjALJqrdh6fqUwwD+jHwmtL8vnyjnL23SfNxJXv7vpp+9pTPo
WSD8oGBlqtr7u/nsKfn3o8cYISNJrcnRKvf+LhaDqSj+f9Q9t/bEl0nOr9rw30J+TC0Wc2DsldtI
S6grC6LPjPMvd3BXqAuz6htgKEpWOaAJHD/7Q1+oaPIOqL6yGWVnPl5ih08DsU378yh1MxFObiGU
JhiJCyFQWyALA76Hz+MYJWigLUdBS0x9RlMgjXyhU5ChMiKC3oMSwKH8kG7zW7U+Hhp4b2SRi2ee
byREz7mjxnqGlr8BmKc2FPMOefGANyiCds5CIjOeKrfUHQwWQE7R1JuDqDXhe65CkZBHPS9tvFTe
ISvRc3nr5qzPymyvi9MwI1j8IOu9Bo1aA3ICODc0a+u7yFSceNMyxOpvCICeDga0SlGNhreCpQbb
HkO6BTYtAiW9czMiu/WxqLNXJVVWPnY8e9FIwI7L3Pbux+xqhCZkcE8l0MHtmXk/7PzY+NN9ax97
2nb2LivOtFWB8ujSJQH9R7viJBtNeZpwxg+daBwvgbnS3xZwvbk+ysWV9IMvjj8ZkhSU4j6aP3Du
TwZNul5YKaK0mXFDk9b2z4ZJiHS0tO+FxR+cnU3wawdpkOeDf42JQj4+tPEIfVh2l8LBfL9NwqJo
xTJgRVJ/U8BSj0nDYqJSAFv7He+cMYMV2DIYb+XwlIe10ofJ4fAQuXVsVhf29xIP2gTK0yPIt1vS
em8EqjNan+Oii3mW5nMfdA4wsNGLpD6nJkg/dUVIdsIU1szMrFn9Jy4UYok8IabzsdJUcHo9FPuP
0EyKPU+HuYgpSgoJufampYvocEi7LziGvHXz5l360BDcg8aME7da+8o7yiCqih1TyRKRmPOrLFuA
seugkLvYFK8Goizii774xVSXVOGBpWpChGgUuFOQt07uo33aJ0IiuyfaAqf0ydMS0esrGL3aNJW1
MihBIgcsPj5V+MfTIS/QSgAT0vN4JJz/Rmclxr5GhaCqFxlUoIJppDI6aB5kP6vEqjierRO+KmT1
EacmOmNAZgIi+I7qbN7fBCH6+IsCZpZICVrJ88M5uoxdrJgK5hb6JmK+85FuS7mU2m6gqGqafykx
Tsmeds7AecWVdnRbGZoqDE0ce+tJAPBCODGFn0e0zdjHrw290GDRwsa7E7Kz6wXC7eMl/w4YLm6z
JLrZ0vRLByNM4hcMZMuqtqIOqVdvOV0dvPk9LkAbMShQ3SH9LkNW7T9NC1DkdEYOssTwbwFebjBK
gi1WbnahVB1bgPUw5eMlj+d8RTmgREcCJFlozHM6D/z5IcBZeAxUr/dmkPfOYUoGC2v+JQMt0mFX
mGJl12DUufID6pAUgg0gRUcZLzHzKFtCESFiTOAiFZNias7hgtLc/+u2LO/yA0SkyhA4yve+Wz4c
08UBVxgIRBpfFxCb5yUv/5yMX/TNya1dap7cFTNjHSgGcqmfcDMaUrxBs5+NDHlStgE01MxuFuEv
rJGNlVVFN00aCtJ7/JdOsM4MBaI3qy3HV2UGPq6zVJ6tkmC7d7JWQUtkknqhHjFkjeZEia+ZCp9O
aWJRGdVwYAhY6+8ot+CfVEjm5dl71DHTiZ8Kfp2C9zsxG9iZfdAF0CmN8pdx7uOaphmkDe8T9YTm
iGzzeGy9rozXK4Cwx7qevqYjG27gmsiZlP0ldX41raSMNu7YrHzghcOs4Ni/MmGiT1TeTTT3Yl81
JjtUUSIeMaqczhBhjYHZ6T4CFG5RxEJQn1ykY2ApytdHoX+VFAP3yiRFF/CLOmd2pKulflGH7FTG
V1/sfLV8wu+Y3nI741eQH1LhvyTfczjZtZPvvJHwcBq3Z8a5303ZVq7Wy+vtQ5xeo3jIny3clnvP
iGuMHhgCKshFDUWFQO5SRwxi9dsRLnKBwbEgBwM6MNd19jooeXUJ2Cx6d4+53EB3ZOMkj7EDqqTD
NYn2Bvzm5Z0g27fG9SygXryfUfwt457pBVamL9sVVkMHCQL2qHX4mceFP2rtMpccgNBCxWeb18ch
v0TMZ+PWfdZy1eulU3ZLmLdfh/M18w1Xuv/fRRTI3Qg9rgonEYO+dstH5nwKZWQkWs8TMClx/ixP
v3pl/JW5BK09Nr+CQrDyc4p1XdOzjOQnPex3QgT2zXenwlNA9amQd3wRQe8yYfgRPMdRtx9vygMS
5GnVvktZGHfXewX9HxAPJOsOrxX35phqkc9LsgJg7Emhw2m6ic62SdAkKPijC7SiRjn0cAhNSvCr
IxmNM1+puowke1ThhkgzNB8tjQjJmog0KGnBLw2cO6Hf0jbKRKJA45F29J6QGGUoe2qyW1L6VFOr
iIsTmGhgdZbo0OVdLMyBe30UzBEEbtXenj7W3oru81O0vTUtW19lwHf6y8/rub+HulYodTWEQllu
kOAE3D+wx2if7n7TbA+Cq3++EwZrOtXUnEFnAkTNGrkR9Y6lpI1vtN7NAgOZYiu/GhHsyodu0kZq
Bu05RMnoTCC/pFq2587vO1x23wFwKMO3WdP1JT9M3m8KQ6r8H9LK50NkOM8Qs0zW58N4G7+l/VPC
6pyiVQNfmlW5h7u8yu0JA8kQbbi94i+yuqUADx2TjAYA+iilAj2pZ0IhCdPGu562QIUdYqPdeEc+
dUayogjzKSZSDVY9eILtPnvBiVcxtPhX+QXqLxEbqq7eYurrhyPV8PXF0yZX0k7qDoiNiaURnNfa
5B6djpUCBFiwZuomek6pwd++fbcWTuznSMOJwQ6kGRpGCMUOapz+IZLZei55PnhYU9tDeGHT3tF9
K1V/7nrM07ViiVTTyUnA5a3+Yn+ul3y1rX+eLKFjMiZU1knqUq9zN3qnPPPaUyKQqvUoVJF3gieW
7+Go00AV0P6SUx1/oMBCFjRHz0SL1+v+zQ/qhIFsBLn16/kmkJrNpDPpaRUcVfGn9xxn4VagW/dG
peDb7hAfWBnwIOKXaMNridIxa+u5Vkze8gOZuoMTdG55H3VcX6Q/ydwwnCjaMElpGjhFqvvMGVeQ
jUV2jPOxcqcTO+myAH3eMwSQnGq6LJlAbg6l9IkkdGPy8UndGpWDdtjgy3OsfW76GU4qoBCs8FNH
PVfiDxoitBXV4QNnwgPOX8aSiLg6Dlq/E50AB7hJW+W7sGQ8h1HGeiYMGiqcnkKrWzc13H4UMGgU
POa24bjql3HxHJnVp0DRqU4IX1d8HpsAA5J4RzmBBtIXycaG8idKOWXUTObg64RXI82l4aA0NqGi
JQWHKEUbZNWnMrBFkSN/3TPnK1eAlk/sTpXXNsSVsxdj+x8DWlaMqhdyAIU/lkUoOFHzTB9Aqmlh
cS1/Wt1Cr5ZnrbaOP6j+vezBMoaUKz48sZ+LAF6Z7cHCrLFklv711WM4jFlO2PdTsp8qTLaOrQbY
yn4ItwcpwayOPJHb8U2TTzbhUc7TgTR8YV1w9/ftE86P3pHiZ+ScCXhQgS61e/EXU1reeOy4Ernl
vuV1OtS0MV4xhzOPH8VZoUp7RnxQ/iyJZqn1BVivV1lxghk1XcopE8L8aVf0XQlHQ0MSgWBmNoho
Jw+p2zzvACicWlPQD6G6skUu/ShcD6At0PFOLvRiXiEtLnpaHAubWtC7jtCF8mzViwo/sEMvVo6h
k6vGiJQwBLcLU70/BwGPhL2JfpHhEPJSkI+f4tS8+rxyW7dH+6xmEvchoxVBCe5aUVJkGjBnI4SZ
Qy2tse3o4MCnA8yPHkz+ABPcRZ3YS/vQQyaHOUn6pD0T8/mJ8EI2GtegUd+1jA5TbdgM7wyFhwJz
hDvQWWpjkwHK/Moz5RNg9hkZqF3cAngWE95gZ4iDLdp3UQDNPuVj5PJSTqXcudN2XAZOEPPxPTUq
aSEGiOymPK/2fVm4FqNPqSbh1T3pJQqAVYRxRaCqv+8HV6UdHOQb9kShD/44iOBuTlgUfil8ITBU
BMhdKf4xZclYHKI4UfkJHkymuPhKaeFiRyrashAse6skLS/eUxZOWwUnFVBIXTMOMyC9zh9bYv+v
/Uj2f+bhxaa1DzrV55lo1PXn6+ShyDn+S75GZPqlEpv+okyTeKcWwlgajHLfUq3LRxTVlWWQpANa
LDchh1XcBZvFpoTzLSU/HgQXgtx4uyq4XrTI/la1aCDzsQsrS1gxKkzIrpX46WNjdzCsfGcG3tmS
0Q7CvJ4Jbq+uikH5VVu/bl66CZwyx9wTxc+XggX5PqKqXsbK1ajt5/M9nnICliSA3vrLiCvsm56M
LUVU7P2jUXIq4zR6R7JgOh8PvLjuz9H59sUV+yZ3pQpdhR294W5BcJkBBHQyKnbnVi1Q7LGCX3CN
eqJCUpbpRDNjYhhyxhdut0y9wE9vnAjhrdok2lkll/H18mhSJfKJK21WwNWc9AL0lpKL7UUjiPVy
pWSEo1CDkQ/1wCjW06IDkRKIiHz9I3VBJMiU/wTyppRZgVDPOOZ5PmfHLh6jf/cf94AgUhRvo6ue
S+JtXt6XEjjptLzCnCmF4RUPuLYEwc3Jr5rVsGWykv6o1kSFt2NhOzynhb/OxWwULB/UsjbtjBBB
hfP6sqd887PVNTX5tnRfpUZPbNEUg4uJx7C6OOyH5txi4jCrAr1mkLT6g+SDZtdNZf7A18NaN0cR
YOqqX722xqgoNSpE6kpFSRxD3OfAe+CAuq4lbRQnaHkr9w7fdqGnt61cvbZDkeeanjEg6TiqKIM0
ZRqD2m31OpKZbc30sNBysCgzPtsRV9HIu48yTqQ3/XeDZDY6c7D/Z4g+anMEiuArQ5XtYoeXsuNO
fjMUnUxgYTIf0KtO+ThHi0tPirxdjzIL3MxkY9g2BJ9yZXim6+mehDuuiuNuoscYuqA1ahVtAUbH
2BXA8rs4ERU5/HpaMhhJ0l2afiH62szoy8yGArPU16WnC+L278jf6QY1AsKw5DiKS78JN/RbLhTe
flWq06tuTR25w+azP/QhQAXtreB9STiUYpPzUSSnncbD/Ahu2uuo+fk8qY1v7qoXE1X6/iPXoTOD
pGfXU7vBo9rIQLzzkFbS2tsJsk84mqH10vbDJ0htAdfD5BoS5QiJTiowKZtlOTr34HVFRIwAZ+7B
UvkHaJJlLS8hLIZnIfQ1dhm0c/2dou40MKjF5QnplAj4OWR+Ess+HYyAOv0OOvlyLiKdRMi37xB6
Zi8S50I2MLoWrquqlBzQ+aBuzv1VHE1aq2K78z5MY8VJYsyWda3HSVoyq18cbgBhZJNFsG93oDuC
yi3bDjZwWOCcy3x9KxalnIwM/NsUen3fEFAvGsAuErJlFv07Ryc8Jx7lfYQiSemEglIz7NcKLdZu
oliEKkkjPB3au70L5Po9boyGO4JZ0/OPwxvq0L5BZTWSsjQM7rbfgEL1UZDseUbMVqVdPWMuh+Ir
hieQKz/0sxduytQ8aY1W7P2LBuspkBB38dA5dvPoy3fgMe5Gqjk6zEOoxrWlfD23benlYLhXpYmu
D9ayLVxG/sh+hH9yp20pfUq33+yq3587vpYcfkNJv8zZBlkqLS5V1mdiJdngvlxJShvOKXYGZzrM
LnWj2Q1ZxyRaFaB9lAiZhPBiQOt0fL1cU1MZZbJRHUYI5MId2FKNJkBeFRNIl0/3/2pBBYmDRBXj
sSDUXbTgXBUuxbgfTX0TUaCNlYMQpOy/ElfzpT1Nq0QFuwConPmKxNNkUICxEHm/W9jAj0B7r90P
p1gg4SNhmtmzMqWpgl0zCQHd7Jw7Ud78QUgamAIAjoZwWeb9Kz36jObsyTanxZKwX09G4YE840QP
DPaTM7pEaktQcIt1jfUuVoDFNLNNDw90wrGqiuyBP0vJoj1fZXvvSwwSW+OpBxl44XUli2BLFg4v
6ci5w66IN7JpRdoyhp05VWLlvaLkTyeYLG1CZagaPTf4Chixl+dEj6tdNB9dmE7/tQIEhoYcuAqh
ZNfuzLQY7myiIokDAFneucQxZg15x9uea6QARGTpPN1Dza49p95N2XYGfy+cbWx/ebAVyqDvXbr0
c8LJglP3I6MbrDQ//uOvi9X/EViCo+VvKPwQdw53N007+bdUHSluWun8MqyyMvx5BWTUgEbRWO9O
RSIkHzT+lFX1Kla1j0d5Zh2WdRwrmLPwHcEmwY7M2P4DSmsm9DZunIlEhgN4AFUREZPNlhLXeF02
xmHyXNMjU1ue3X0PHrt/8S7YOaTrGLlXk9saA1RBFXGxhP2maQoJVNktu0lm2vKlCMp+egTyu6bn
vsjnpdBw/q/SoZQmuxN6nVaEhrvqDwvjjl/bAp1dQZZ2mfCPLdnMjOuJ051eid9dfuiC+P3LnuCv
2G2ScFMmZsC3GACGeitEO9fXkTaTXWD3BKKGftJuYmDJaZs5pktV6aZC3HbgRbkUyU1fNtxYfkd+
DUPcCbNRGTqsFfOTV05S/ikybtY+OmTwOSG9b0te//zrQzqsqzWlJsQI2GAF26AvjfKV5dHpVthe
hqJcFNdaXRF2aDLWrwuUznTTnH3vnRqKxrE0ABWbjR1P3Hywrh0aPMoYqMa66r9hC46PfT4tFcjf
OBR4ADlDWHXdiGzUsYANz34B9ZTKHnpxfHe2nHUdKDm7oHD+eavV1sk/jDcgH99ZX1cJRPMtlf4W
zNGgFY9PHojnFLPS+AMuAersXSWy/dal7rMqZlOteh2kvzEaI6NRxGt3yb8L/R0iVsIrEigPMo5r
RxHH0pAjagFoLaCS1N6zvK2v8aIAKacZIb8nxEBe+vajkay6AplwtaQn8ujLuYVvkEd28INfIEoG
HJeoaLtxt37qcj5zzA6gscYbos9h6H0LzHGDO43AVuSX3K5GSBCujQpGF+PBlTWCmWbB/iuXAHCA
CCIjSUKla+6Lyx6L6PApon3OfDr4Txp8O1Oo0ukf3Wgl7PUJYH2/NjuYcnZGo3c5iMDr7FNtZSwO
29uiDcMaG0L5XFHBpNNiyfXJerzK+MTVGp6Rsa7/Xslwh2PWyxYtocSZmGHfQDDpWsZa3Fq7rRqt
vTqaMvPCgHFV7vpMIX1GdMWOoqAqBRM1ffe3IMH2/TWAKfTwmYl3oivcNlU3Rosl1B21I9YcvHlG
DCTpc5CdczRlXbAQ9e8sk6i41GtwxamtHKf3LFKBKAfvLuDj9jNosrUSZLgviZ1us4c9QpBoW6AS
WtED6mV/69d+kqhkiS4YSlSQenUWq8SLf5ao8Wb1XqVp0IpbaO60gslGl17cCrAuwzL5I7UQQtXi
d6McbqkLZbqisVqQZBN4Qh+aWLf7YkbWZTZ/DP/kTF7KHL9NZLoQOwguzLeSim/iXsNVlOkBV217
XjsQLkX2afzoUvbm3Kn8alI8EEp9Bz7IndvVmi6G5fasaax/+3YhMyJqM2NUxG9pmJS3j1BiDTEr
3DrXXzwYEjAzZQ11TwjfuII2k+F5aAj1DlBfSrE/sluivx8XDCZDSdbubDQwqnoZ6kUD8a16Vb/t
I3ou6KNtRiCjXnE6i3IPDMgvXpHKa+AEBcDusSb77aJnLFWMobkEgzKGLlANSzzA5KYkToTjdzPA
bUoeqTb9kFsaOyKdroM+soS2wMlJgXdtpS+TdVjKcTXxWXTGspop+czNHGtrdCvxyNgFNTw+JLqh
ojcNxa7jpbJaGHjlHK/0+CMnXTgTAiwiVGThrCcv87v2+SZPXjjzKGB9ttjRaMK8VW9UH2G5g7Ef
U4XKJEJLkypAQRvGRaV8RkjqIwR9vjPnG24d0WvqBOYa7NEiNmUsyc8sOm1i51o34PbQ40BGmXcc
8t8ZTOVx7NrQlIL7Yd2TaatZ4ijN2supt1yq7CaT/b+1nAixUY5e34/hL47YJl6Odzq4Q8XRGDMt
EYnwSV/3RX75IDvP0LG0gncVkTghQewXNW2mYUUA4mJdkykfNZC7gx9UUXZoVk42Y0xjr0qPc9i8
w1ADKQEkS1bvpz6rt2E5bdyvqH6hWN9BI+YH7l0Y9Jm1iTW0Qa7om7IW5qdJ39NEkJmlPAA15rb7
bYCTsK9JDfUfXNG+PtQtSEFsGUlRcCyyLb/q9WwYeKthSy/N+RfRDlYV0r1FKO0/Vs1ETZwCCVGZ
pcfUsvtTMhyjZSQhXD8+yGWtMpP1Kw46fg5YBuSb6488zZ8c1hQvYAuwksr6Scu0WhsjX2rN3ro+
xOYYKGTytbQed/Nh9x65cYzI3dEgSnR4516b0PZg6v45A7L5iCLy+aLu8UJDoBbCv/v/oAKkMQ5Z
/zO0ApDAJfrAm6EMu0HgcrO9QOZ81CMxY/0X4LeHw7hjwvbkX68MSx6XvIfbIjj4iMaOMpEQALuS
7oOkXWW1tBzHEI2dSTC7tmc2JY6eE5UxYsJpJSeb1NAmJMUiufKXWCtsyqE3tTqH1HgAaTjsRBQc
NWdOuhj0nZLx7U/j26GejmqppZkN7Iy8+1hHXQgPEct9zLsRpbVRag2P95uOqLBYjT+vR7GnVsQP
eQafC0pDPK52/IB/+i+WHxSZwqsMbFJt8pW+mOnouIQsiy1bIjmzfOjSpvmnHssumyd7lqJVmxIS
WUlVUmN/NZaCh8b3ZSBskqMsn0b/YV97rfVZH8g2FWx8geZT8qRT1Q7DMRIS5yiyRv6SZYdQ3LVA
KcbFjfQ4GQfSPjzY/b3i8nulLZls6+pujTEXHRe3UNMs0WFVB10kjVpD1+YblPJE5eZU9olHloUI
Hj/fol3/r43pRE3Gipri5P7UaEXuELaoEAHcOGhjilCYl+gE2004HZguNuAOnZ2BnrhBDkjefTzn
gjqkIcwhdNVCntbXS1XojZwKO1PXhDGNBbRGseCeVIOqLvJSyu+tzOcRdPsI50P28yD/GLYcDqrF
K1kinL+mWCTjHHrYJSUMWRb+a1NK4NkcVI/pVKWOULcf7GuXdan5+E0TLnJ5Y08KgZhgNlpRWroI
vZ2+wi3UHWWNOUVBH2uYoFH2m7P+2GNHXnNCYDH2/7rDmkHtIC7vx40TyuXqo9lcvOLJYfHYSDh7
Y31XPV4hwZDkmi5p+yAgQ+frAbufqYC9Hht8pt1oN4TOi0LNlG+rGdf73qu+/ooQt8/gTMF84Af5
hGvqH9NdokTnANcXfKuCuOXuj4oLFgWn3nGBYlKE7b1gcqz0pkYSHHCTHbB/wcj+jP+JqmjnhrRF
+0baI6QXaW6OiPdnrzkdh2jLGfie1uaC9rXHxSyqrHRQkybCJus0i5305P2pWZaUSiRB1+byJLYD
HEXN4DAOkV5Q2sj029g7cBS6Yo/V4oN++RHVaoQGYTfbz6wOEzAiPkTqv8zND4HL4mxylqZ9m8vp
ny3OcZr/TkUHnVmhc2nUZjUJj6xbjp9xakTHdbIPSbf4vPNnFyoU32WAPrclWbwbftohAkvu6XgH
S651L4z8ggttNAhufTY3NT1KHEJBpiuBCZLrauUpfV8MxbZRsxzRqADjzVlcGF4pEteIQnsVyqXH
Q4j3RtVxhfqJTXO2ZcJTXu5rBzEo02teZAeiuZ55FWT7fMr0d2TpLQCMYl1rlSombxbG0R5OS2kp
8pspEXtYjOdQhcyjlghaLny4wH2GZKS2N/87ke+Dg00LbFikkkDmtvh6McSeU5K+GCVltNWhuU0N
oMcCG8d/nx+tlFdEOAOAaGo3mRl0brgKhuL8QERFQTi4xDrNQNgEm4R/4mYJOYemqZezuZgiMuDT
ehn9lWiBzF89QwcvvWUMv4fgcmRvzBa9TMc8iPCMtq6jfFLXAGnopaGD4Kp4bKltmeoRCcyhxYG4
qjROQI9KM4xHc4BHNO9YIZ2rlV3AI5MltzbBUxnQiFNhoqCnGYozqmd5RRMg3jKl+zxqRkF09d+1
NBzDCgbP9QQENXQ/leU/FoqYoNtWQ4gYhB0b0pTRCWs/RHEzxpuQTo++zpZ0RGtkDrmFZ8LIPIsh
cXVEBJwGfC9fP2u0VTg7q+m4Ec8XXkSVhKg1uA89SenKd7vjpBR3w4fWAeTEvvEXYazs5Hl+qsR7
q6S3GqFQ0xXq0ksoOpGZTYDyUfN/2nMUErVt2Qs3IYyIEo/osjcO3Hcru5fXayAYg5kykankviYO
IihC6AJlDSU3VD0fSLGUdrQ4DE51jvNp9Re+FV50zECdZrVfQXJn4QrnDkFBxcSVIOH+lVHvDN7Z
mP3TiseFu/ZuIoFvfNsOBulSiZzaY+CzYM/0PZd+Ec5RLPYdRxFjBE5LFH0a+Ou4otFuz4t5+D+5
+uMykG0tn/e1+e28dXmfyByr4wd/LAxaBgkeZWtW9HlB0zYOdbTyEanHw+O/iBpA3hNnxS/hSOUO
McpfV6gD+RwcWjr2eC2/6Bku5Z16dY8WvbTk5YuCZIdX44/2G9NjTnd1aZ+XkiKazOI9zCGWZfrh
9/67wK9jmUAYIECdqnStUwVP2TKul9EkIz1krTfSSbfg6vQoC0mPh8g1oJJ/sZSPD59EEN5Wt7aK
UVprcHZIgE73X3+bgqtxaU2cMzbODBfkWhLoVEY59zYmNqlCyOQcqCBbdvvCA8s4bHPaRPf/z/SI
XR5v8JBpiodO35g6k4m1b0NBBKMckMH8A5Hj5R7XPOl/HatYd+QlT/4tYeo2uc2brNDufg+2Fv0+
BOGs/CmtmPd70UxRLBh7EOQUTm09ddI8RuTiEPsFhrTsLB0FwirPtMllJU+Q6yqhIBpq9O4olULA
uCMwT0ivhLZbSVKPivHGKiXA6r2QDhA2KyJUdy7M+9Org7JAWiGdA9Upd74IPJhSp0YRJohDVJwS
tAnjjE+o0zxfeb3pMeEuSHTDK8CUxH2UwXxtQIyIfZGxResdvqNZRYF7nou9ZsGkIvJfcbIMV9/7
d20CcLhiP7Ssw7SR+gX5UBcRUAULdoRcKNe1cVgbdRslmDB37aqL/we07crSXGy2JtM79nLz4sZd
SKucemn5b33lk0KYwTVss+MTc3qYNodXMeRAPWM0V5jriixZ8GMRlXyflHzLF7OhLZNntTGW5hce
s1Kv1f73Kp2itM26+O90POozFgAxlOvD18MtOOLWYJH4Aka9TY7uNDGJyqLdLFiEv7GzS7nxYoqZ
kHWegHiHZovCPUD7ZNckBzKda47kFX5Fr9T2TBjBYH5MEIIO5DgWD61DY+hbRNZMYaRbyYUjacR6
K9LfvCwLNNuEzhXy6SKIseAUIqrtpMqNjvGQcBmxShjC6rv+FDhUNeRt5q02aMmH2oBorf3ei52g
xFZ2SSPitjx0/Ixv5eXPcYnrdTWBwyxqRWEnIKux7JDP7nmnbRvgOQYd/j+flgxs+FAGSz8v+Owg
u8Q44mn6W5zsnIg5PszwsFQdq6MX6BNbkw/MTO8QpJ/86Vetr5aB90aWNP+DBNCryisc6fgrGrxM
ovDPP3qtfF7HrQ06LbeVy5WsNtpAz4L9dREhQvMfJsWuoHxVo3ngKGqNaQgeqgnRnOA7DuXSpTB/
YLMZDzN2ByMlRCmNA94gKo7anmJNuPqas1v95Mh9iEftxT8HfSPkwqrYGisIU2Z3KD/kjsv0lEyZ
CtdHZ3as2Xu7WpT7SyYH3Mo7KEX1OQAQfncJix/Elzpu8Us874cTJMmDp4cTGH20XqWdpoPYfbKE
CDMknLTYg/JWUPk3YzvERZy3eoLJzdzv3Rw/eq9mBvzK43z9sAzf8422C/tRsSyd6d8ttjYhGNtk
Be0sKZhDXwZvApP3gEXYDeJBBo/mxYI0ktjslmAWNvV9chgtEoHaR1F13uyH0ekfoI0vlcHeeG+z
QkUAbhTIg9mQeRagUbKgyn5jc5VYWxXrNNmkCA40L28L3eUBol40Rq4jZ0MwTP6Q9shTH0Ru8inH
B5meJ5LI3Uwj8bAwzJryt1V3j1Q1dasWyjWR8cPoJj9mFQq6w1i+rFI72taB/NXR/x5qENvA/uCG
McDdAlz5YXziGYSe+b/YfL48v3sVa2odYQHkZpoVzxAzFkY9Jk3RT/3R+pLjXK3NcpGUW1a7jJGv
zGuM7mtRcO3YYa0SMszZ2IeFkpxVB5ERLIyLZ1GQlpGWzB061zsYRLpOBsHQJo8I5pbFL70abDZn
3cGghTwmuavyREvGTXiJEOBNhWNw0UoD9nAt45VMJe30nxU/0ttyW+rM7bpqa5cfqeRR8LvXtbjD
iMCE2ffXr5qani6/AGO1xU7PBSeVFmSn+c8rO8cyWyGXSvGz/8AFZKDq6AuIShBGz/Jj3E2QTyum
6E7eaFXEUcA7hQfX+viX6xoRTAsWiM9mndPlVYpHdGmvzAizAcji9VHI7luyBBTL5uCpxcWBXOCk
SCmZ2qO6cFZG6InbLMpKUE383KqIHTM/uNhUkwr05bjg6yxAVJ/5ac7edcebcExAwpQujn+TPd5d
IuwOfD6PrssHg5ke9JZMHKoDyVBxMAk04KAGwT+GLTZ4X/tzbH8HxR8YN4g+LvsdJMZypydMoY3W
iktYargSf3bM1dP7HneHSmk/jLn1uYl4LdC/KPhUmSVED4bIJ9ZGF+BO5l6Y8HNG+FNoQ0LFNr40
bNQDtDK2W/tDIYpEn58rFOK2vZutByH7enrkImDe8024sVTirpXTu9o1H0/KwyNkLEvKqDqG6qM/
DmfT4PBO7/0TN9Bal6vpGFkyrjiPomnvAobBLH3trfSwNrdeO407fSl9H1nMJtnr5uJ5SmyDQ7Qn
yyKwC+g2NwBfmBPRn/DG8bic1obHZTWBdL3417JNOnHml/dtmakankAKXmhTd6wL+o6jPqeDemIs
15kE3f0qA5kYk8T8Av0PJHBtE2CgMIVgMvNBI7tfBu+YmJcIPGSLVl3fHcRQvExlZGe5LK+Wuca2
COjWIBJk7rT6y1oE4t2PI+57cB9Ov7Tdf4VjGEBWrc/NZw9FI9ZFnPA+UPO/VNfDDlzDSNyC9Wa6
g9SlV3Whdeog/J5cO+xe1lTXHtCPS/fk3S/KpQTqJvMZLVEga8X8uWkoFepwlPPLzm4yKj92KGEV
OaiDaEleFH40/mrMpbHS+q59fTX/2NiEF/b5OzbEFBVouJC1AkpVKpFy7VEzBLc2YiuJLXOcC00p
SNSxrEve8ENuGKJWw1a/6sUN1Vve3X2RxlkJJ4GAI+NIO/+R8xHvGEpPhroZWFBmITMfb9zqiZJB
OfMgppSVpFpLPYdUgU6OLh1QD1WivHve2BM6v1RTyjfgUvk0PchzEuenMkH0eJyNURLnZ4lZkJUs
zQy3GB7HecUQLw2lwcIBoDG/95/sx7CtqqMGF42S2S/p9+MS2iKiomB7xirqi58syqv83PwFbQSe
X3PnhIv5oxqtWELpguT0naD0uSEe8zWg8Y7sa3ZAWA4pHUewSzvQJpEIRFqW8JTBgW37/ov7hxG+
7E2hlMb88j0OFQa4t2QWEORfB7Y751nR1aC0sV0TWQTH6f+wWTILXqTh7wVHl5HvyhwMC3AjHnol
8zfUuxgP5IumjzFIEc1+DdzNkLq/OaI0Yxczc9l2KsCMc5Iu+dp0aRoZ6qJnRqbm11M528hevzzV
7dGHvu7BC+eb02l8YjdBh1/Q7d8oXErsG77TIsvr966Hg5ZWXAhtSUZMJulWShGTXZ8H86yl93CA
OslqZZk200n3TZzQbJfjgRvG0Ddw7ajQCXEA4g5fzpG2Y1TmuwGyO+ouGeH9yVlruoYKWrVVoefh
TNKjDttNBqzTqrOCqJreDrXn6ddpRBCudaI54QmCzctT4HgK4Kj/bZPbv/9sPiwDKttJhJCw6Db+
32q+mrxk9IV7tWCc5zaXpq+2AZ2XDWsJ7gmqEdilaKVJVbUCtlAQBvN4enEP8VEogNOr4VsaRW0b
5h8enku56thDGNSXjkXC6v+lfDrkjhlFl985k2iaV4mDaDpWV7/GgERr4EOhy6AY4gstaeGZhzMU
PmODGHwWg69G+Pbmi/4fZpJYtjlYCAIRTpvBTnc6Ab5Gj9l/M2mI9nlKzI+xmFrobHognBVSryJE
KShQ78Tt0OYYB9U0CpjBNUPKGRhpBznvkzQpn2KEQlOwJEHZvUT/gDh0rX4VeGeSoXV4ARHxObw1
G+PoCB+YRFiC+RsRrIubFNgsPJ2nD7JCl7uZz9kfw2wcxJCf3P+51RrErsEKQIfOfEvrGsBY4mNG
sIB+FP0lVHGJ7hBeeVC+ojApQPvjrDHYiGp0j6ATH3g0XSGXmPt2SJsil8wQO7uEERtGZJrfPLmT
tuLTJWxLf118ziOJH7k4OsDKLcZ8nTNDQyLfjHJTV9SWlsIcD0GoPHwP3XabmAxLf12f10HJQgPQ
KqGQBKnD04WIx91NOXaQljOGuddZoGb2PV93QxamF3sMYTTKUDyBBTEXZkXJjomUiA7q8rGg0dde
JgLoNUwxiVhQw/aNgVxM6EoOXCSP0glR/47E0dSP/osjIiLHkR8FeVffrZUW6cZJpQ6CCb69Bwlc
u6mj08FeJBiAB2lqSz0IGiOhk6w5jqSozEtJSi7yQoaObBl6gMIvi7hpVqP2/Hdkjk4yNBU6Haaa
gmgVNoznXPr7P+Q2aBbmxcGkZTjb6vCf64gDJH/NBn/JkjRzPg0gKMt8LDDLW5i03T/9phLf+weB
DK3y6r9eQ0Xg4b0PnbsHf7DjAJKo+nX5xQLJTI8qvrZE0LpUqEIrDpAoIWDgjl5+CoVeMjUeOAyx
xu5LRs4r2IufXPMqRG9iOgP66FVh7icYZejZ0nGVIzY3EC53pZr4RJWiG8TsCAXzLA6FyP6ZIqOV
etiZQFvbIa48MF3KOfupmmYyTGbmUoB4UV0OccPGmOcJKc9xnoGmWP111q5KCFXCb5TkHwSR6vf5
O7hFs1H6w9rLl06oNo1ccIUmcxf3AntQTNjdmvf+DWL1L2Mct9Q+IyZpqLVulKxvHCjPk3C/fPir
ObuQkK/ExThAf+4xStn4neBoVC+m0HHaVdmo0mZR/0mzkxRHIlA6wp2djZ/0MNqeY7Qx3DTWsNtu
K+nuBqCP7/BTSnrJlplcwcpyI9Nwmitdlx8O7Foo2wPytQkSIHixFNc1aOn879wyoN/WpoFwJL2U
S/Avq3O20xPIl4cQlYcqHqASOFiIHADpb/VXl4VXAK6tE/M61pbvf3POAvM6epmiIbVBgaFCkfBZ
+Xz9B/4q75nevsAkmLLfOAxFm3ZREd871Y30fB+guOO6HwG5PASQsa0HwFsCMKlEkEiCKClXZLMV
W3Di/AMYS8c/WR0LYUuHZ3WFLw9sUtnWxVF8N0QcBMh+z/H06X2Wh0w91uQ+ZnZO/LrX75j0BO29
xJSs7O8sGrpiURCSnlJjCSamj3Qrubwm8ArcoyATF5oiwJS9lH+7oRm+bxwSQpOszslgFYg1TppU
sWcveFjHeNAEDKwptAbzRPtFG8bf3go25smtGmM5alpFXjFxmTh4s045KoVXv831G3Pb+fgPkju6
GOylGzZ32nXKzzMKbKKa8CleXF2OnaeIZ6z45lrRsT92lOFiF3LL0KXQyt11nOK1A2Lj7z6Tb2rT
0izrC7Yl7xSZktD1yo470BUlCwQ4wAU7+W8YX9zLNnbv5tkHf+h3wqyvsw6Zko1K1q6sbiQo+aCR
0zZ58t1WUwpNKYR+P8s7yPt/rKLGJmFkHjn50AJahenvukeg3bW2O1dsIKAPhK3BcgF6D5d7k44j
yd7OIDrNj2EJd6n2i3ZUTC8/LpDFP+RO6tBDDres5Z8RctfihHqb1QZbsEwhdQC255dF97Bq02ep
vYl1KlP9Sm7aLAiAzYnfXPlCEp+rW6hrOLvSidPXgOaqsOVVS7FA/c9vJqaulKfDhHE7hkRZN9iA
yeYp/riOQEJdG9MmVMJVBdpQcaKy/5R6EG4qiEfC0BfcskQ5kjPbYyU1WJgn1V1STXUsm7/AnHKd
+a7h1uxOEPcPuz+XecRCBZhC9A8WflLFLK4FrkD8rmlk3ssRuu9mqx6rbOlzENmSvmnhRI6AG9R8
NdPrvdFtRvXz6sQJVOK5tS+NKLMNvozpIllM/3Zs7Zsw+fCEK94tGn9Cu+Rg4xfjZaZhxX0o7ZT4
8thi1vR7+/lTDd73LaNm1GeuQXR7f6fiYhnxyMLfBNlquSvMgMyqmJrKzeJLmJLkVoZSm9Me5lLm
Z0Iwgmp+q1j7nAIDHOFEl2x5n07Ed1NXzJdw9EzNJBA0Ydxtn/hqqkSL1Y6g+c1DCs6BxasxHkhT
ySiT2pbFr7b0PWjZflPuz48Uxte5hQ+U61+3QbHZojur9GFsEHZqXBNRARrzqeEIwOxQ+TQ74WIU
w4zVpeHC8jw2m0byXVkc+CVuBqqOkdxKM/y9dXKG5QEtulMfoDazKzXFnNgJVZzTJOT7tSmfVK1l
sCVqvZuxTR94dTfw2jBOKhXJ9DvmJqn3F9HbkIjwETN4SsVyYwMUteM/xHyWdc5kNwuEmgLQ6QQb
Ucrgs3lNHOkHnGTa4oUdCynaUTahu+IZsqhM9YesRH8XdC756Bcj72ZeoURRJzNnFuOarvH8Jgwr
AwfHLusMh0A3/ThGmSpP5j+z/jnxfQ6W7ualIVjB7lzGAOE3kmTXmg2GRTMqGNVPuJpPfgtR7bZr
VLrgWiDjmvuUny+nHaOct9QpDGL6lMwYZRsbSz5RHSchqtCKyIF/ZMQ8eXDZyovpPQ0sWTXm4UNa
ciU3/chUBVVZd3lZHaFiEWuPN8exINOYsPnbj0SvRsn4cpu7vSMrvDYMlg3rOyynbAxfgyVAyoOF
KNgSvVJJ2HdscrlbaHcO76G10h5WUCaA7hEE8nk3SZUEe/xAndBTuJlnMJWl5KtzNri5oTgTuPRc
3qHzDf/YapJnOkPc5EeB6vVuRrhfKfPeJ6HfP3j37MrzK6dcqxFsG9N/lFM4dWBUngTedn2XYlHE
BvjK3NsZ0Z4Du8ZmmPgtjblXDr8A6680BKmo6lnfwrDsHOk8V0cCHc5giYNZ8hpftXbOCMdskc8p
Ip07sDOcHojMTalrC+1EbvVag89kqyl1J6hVP3nQ7NRCNbsvHpCK7xRxcmgQ8mrVQnemFiPFujdL
Dj+LybBby96RPRpw8cwUz/RwqpcIouNDPRQyYExcYyk/WDO97IwG6OZrj8nWhXI7yfIhmHvg6/dv
iA0lKn8y0lbSUJu4yOaUIG8KQu4sKCgrxE+y8TK2D1zndH0VYGiB9BA87swxPyp55p1m2RpSawGx
nTtLY01RbHDDBwMScqEegOuhMimQxmTjrcu3nwUWU8YpNCqpLTjzGzpmycfLW8Nlv9/jq0l+NWbE
t+gXxftV9Pr/Q9lfNkM8sPhfrC0iUzaqLzfca1ueYgHD9BAWpDvxVEs4T2iGrR0FJoab+cIANGbx
fVvCnJ6mIcz8w29OzNQo9L2LKTSdRx4Hc2OvBIm2hqrpjSNHP4JBXlqdxsTPEontI4x04nP0Np6+
aAhH4obzatQ2394WMdX/o2iWE4ckVRDMHOBbEVQNnfh8eJsVoHMUnhSuhrtY/bi29V18dTUuUWny
Iw1qX5OmvyPjV9Jiym4RJfhD8d8Dw3Ld6gu1tTtAzGHTczXELNZeX36DB+2bHS8+v1l+9rwCB5O5
+mo7qwLTR2o7wS+lRmof93vDZk9E7yI6E1BZujw2alfUMcZCJPcBK/Fpr2kxNyS+bRh/urDZHoaW
+w3lZiqAPJnUbBgz0cn7Huz8tCQs3ZUfjVlpEFuOV/ppPDfwQCjtcuFCz71Wlwt93bfMFe3YZjST
z2i4hiUDyNvTrTwgAVISz70qzEFwimgGVjVnP+0OPEKjMw5eKW2O6dbf7MqB0vd48lR9/i1VsTPG
VT4iJciRS+KGiZ6lGjnu/IVlU3UjXR019J/2RUchBZJwXY2w9WJw9mzDu96wd9trD8v/oG0inAkM
YcmbgIbYB6i9NuT0b/V+v7oyj3O5bnrccjeN+xGin0POJD9+U0F9wOmiFIFMNegk2BO5RYQXiktk
K4fAixHTUxwdXQmkvWOVoFuadz/7BxtSBetkKv/gMYE2M4OqUWVvTT0ojaPqo+7w1XuqgINa3e4m
VbV4CAbA5vjfxIuy7LNSxbjN7Ea384eDMLIb+zta9g9Hw03MyjoBvXNAfqyS9AwqGEqebdjyu6vw
iKcbYb4xJPIDXZqGkmUyt8GdlZM4BZOrgB4JqJY0Yk7V45nxe9ZPs4+s+FAHYdN4745HweM5Cfkg
BWXPP5hbcQ0/sgKSJyNIj4vrgwPAGMUaLTPs6LpLQ7h/N0kYu732Gm456YB4A1cPrj8G0+as2nyh
fVcEDmi72w2BLVF43YODHzT9qDx8TR60Wh1zH3q8e4WdjhaK44Xwo8eFgR/M7wEvIY1hk0zvelDL
V7cr/vU1niOY6YtulawC/53iJIaGZgSOdR2Dv46IN+iUPUkXiTKz2kdYQ9YA9QbSAIS2JuL9NhWD
0TuDxTAwCv26zQT+9GxVs2PlbN/Hw+HiIbwnsxLUi9v1fDnxOt/Rucbo4R6coOTWAm/SC5HviEid
zLE8DQoFCwMsHT5mapPrRNn+Nio3BAbd+xG768peH5on+liG9IZlGVkd+ITSpVRSKDy9JTzkpRE6
Nx1dLoKe3r/QIKFcp+IaCuazAM3Z3OeYdXeaLzDkAzlZ0g7XVI787Z8bB9ULEiw//Km6wV9BUZxZ
sTf1puG+NbUwZ5TdqntkRFNMykDZ8YFlaQ/8wACpamj6xYfLN+1Ex+ySXQILna9e3XMHaE0H5LJp
Wg0EpWqP4Glv0cib3VaDU0bvPenfQbzNiIulTjj/DvLfkLv/mXT50wsehuzpLDoUUTFbrBkWoEah
jVsHyZcVvA3pgcrFuGxAlrUl3vlNFNt0mknYZXUyOa7e5+EGe4itOfE+wV+IihWcgdTBgLSRQHjA
nMJXaqh+U+W0+g+en2AZISiD/trGslApDBkvRgjQ8ccIbgDnxuMapdlZrlpvdYXm/t8iECC+OJds
KmPlCQyzljhgWmOiA+tBF00WP9kjfBjGTngIx/5ICVjQbHVoMIZ3M1DTGThg84r6sp/itD+OEJeH
z2mr/F7lhA6wWU32Jsg0Ntqzmd30JIWjKvLZT+6l23bW9owOkiocpaheSmDKvtNz0jdTisJz5+MH
MAmfjDF3MDTHq8l6GCmAYgpi4s9OoAG3O4J0LGau47Go6KL8fOXtfySU/ips5GYOLgQWJPagaICF
vsYeNYCNtAQojxWBxmXvKcpPr1BRbHiDjBri/+v8oxY/g4HdJHyWY51QmZm/WQrCwPc7JoXD9kHH
Sb6VzjGIZKbjQu00ffZqqWA/w38bJxu4mjbE2g0as3aoHmI+JLdxXscJrzXcLZWySRG15Glu9e1i
16e6YwjD88kh6OoJ04y6oLST/Q+gCOrKv9inxjerFNAvRFYguLHCpdevqB2hUNquyzBl/OSjulHN
Qk5w5TblxYP73PHNQwkRPJgtajZpj0hra1fIUecmdtTxj7NILyp9Q0hZGmWtSyMBvVwEvmPL9ZyI
8BsoPZiFMr9PWGWK0a+adaQ4wYMY0N+7QcmaBsXWMkMKVm3ZcCILUcPakbKJcVQbVamxfVnwG0Io
cBVe587lod8EBI/Bt4zojnuyui5TGkpI6e+b/w5E/Ne/dfZXDFHLF4hZgozuLqyfyVUG2THUXMsg
whI8+ZfL7EnJFNZdJRn24E8+TXVxYu0V1jXYvzOoI0GEvZyi4r1ddNZfIVLTJ8bgURzmhiiNgPLk
LuYA2R4DkEMxpAEk4wv4aCr/P6Vdn3FMRBh8nSdWr9tKNrRj4j8B3DCVLwfzymbyM8FWoW+PZ14d
iHiBSBU67HZ5BkEt4YCDBGRibaEKdhx8GHwYU7rZ28TXasnfvFvvec5Y8TNmZo8XL5LWzxgEKLQQ
Pe7cKrWgt8a5DLM6kTDf/s28V/KQFmiTsP6qpJL+J5w+Y7vkFz1lVicXQyTWW69ZCNFyTp2n6FNj
XkaCW++YLvcaiszNleLS8zLE4+masj3vMzDpa9kc6XcQDBbPbkoQCBqAuQQHY9X8HvmJG7560RV5
iR5gIn9YnheAO+RGimTC5unGXaQqtqqCl2KJyyM2rtibHZ2dMMDeTENhof6sIYTSiXjuoHh+RHNd
WHUu8SC25KmtXqwm54GL9JWC6KydAQvWKVzdvOCiVnV7JGeY9qkhGwYeXY4KIJtrjAz8V8ELoRVH
DEdHtGk/1n4LDFpctBY1qIw8lfayn/JeULVts1jxRnRjHiJQoLf+Eu+31zBCC+DCKRbiM47EhJyd
nyEbrZKAzoRT6Mddtl9AzRl1AXjOdx5fIc46kay1XLhVGe2c3nW3lbaj73ISjLara6AWGpqQkkj8
67lirFxY1m81JmZhooTTTkwfzz3/a4sBypUT4zIpAPBEkeDPiVat3yFyGSFJjj7mrKORXUg28clp
5x5lHAYebFrj40wrUrx/tbr6A6UV0Ynou4gKlW7aTUxUG7scWB9WKu+SwOJXIFTZuYN+ymLfZcYL
nY+Z2+wUttslzgFoiciPU3+gb/0OZBAfP9XtAFGezggACxDzTyLWba1XAeplf3oL6D/Sne3UmA6+
wj8RxY71ikYMlBeZ/qYinXSbsW4TnkzpV5wH4g/dknBZnvHrnByaMMOuUDwTsyZ+7YXb5TwlMxPd
I6iNSkYVZKvaE5An/cNLLSHSBapxZDwA2Aa5dzuyfbIbfj37ylJ/I5kd7d6h85i2Ln7cH+m/5A/d
oovJ2rGsJ8jsA7nGlPlTPyE9uxPj8eYxbpjo1xYDdRXPYtBufMlou5ZTEn52rpJCYjzQ64DrVa8Q
vFdmfaEGcCvT8yw+YZE+kHsl2GTKc/HnMGG0K0u/vnSxS3hT+sKt1unfI/icOR/lnSN7+AyOMMkf
10VO4x7An+eKvJWPhMRxob1K5AHrug3n4dlJ60ixO1//vWBReEEBuW9uo45LV/T/q9FJ6ObS3zPz
ya8svXCZWEEHamrJUPHyLqUvTwFzmQxm0V4q5DLig7Gik8FPDM7YvdqddViS5B9m6lA9q4YdTjSD
HvXIAFQlI1UiLsS/ziD3mQ4L0vHU69lkwusmSPnYxnOQMHdEbiSl/OJNIK2Ce6DWaOZ/dRw1qH3H
HW4xsBXar4rCbf9BWl07hH4CqjlVBPJlrkJDnBFrA6VMWPNOoLcxAy4FOilyzQTKA+4W2VQPrG1Q
sJDIm9W5mO17nEHhvX0ZHK0EWSgbWbo9CH5yOcjhyuXQfiixuk4yxnzgXFu2cQGRqd0Retvz+FRk
UYYWQpl1cEJXhj3GKvdeC6B7oUTUTpL7bu/uaXrX9De7kdkOxUWLAJ1WlPFfEvvZtFhGGT08Mwe6
u0apoo9esnWanBwTxcMDsH71fjTyTz7Rnzf9nHx+SUk9ywarANYjfo2Mhl1mR9rxHCxLYQJoJoOn
c0xWDpVliFVWL5Pr86rlSw+mqvHd8Hrd4u0xVLGu0orCap1v/OULRZpCDdcno4RPHK1HBWgLX0Zo
FcfLzry3PJgKoftQT5fEHcZ9vI1nUZ4MYVjhQMQXFraRP84Dmd6YwsFdIpQNy5pO42UVc9OKZ33l
ObgO2b0fOFE50pxWrg/rx9pPG0cpdML6+veVTKZ23ulbt6sESPUReH38zqBYLCLE/F1tPfmoPXQ/
KiqY650YKisbEVE0iEtOibAvzPOqUngKqpN9GdZGl6wpofta3x70q87ygc2RWJquZaE459GAdNLN
WshLme1JLqtIorfLRRKKAwjLKcxmFW/Jdg+51+45OHyC0Ellr+q1x3p06ssRVZ2f4A1n//GY6PM9
8TuZK5myuRjxz/IN4/dZoqQ7XYGJe0kHZsD4laGEZhIbTbZNxZctmMnBMyWC7/DvqrSJWylDIq3f
LW6I77yae8INb1XgrWqhyNEuziSAssn8Opkp6THv/Ha/jUvyLYxPm5CYdB7SEwnCvwSlWtbZun0R
sKkc4oMngNFdaanQAocKNDqfjsJwkaXA+0O9I/FGfoxUjo65B63XM26ciCwe2kU+x3LgjcUCuO0M
jKWp1Au/4HJyEEetQXI1+AJBI38AUeh9ZIT6P9gyxSg8UXxsvC1VBo1oKAmz1MZZxKFIDvNqDamk
IwGMKkVwW95TH5Tw23XkYMXaGOCgFlLKbVEwIY9KLAf/2fLKZAHV/5QXs8QhhssHX8LahknJ0Ugo
3ErdxtMJUZ2UnmevGvXG2fMs2bqLzUESs0sU3Xyeks06hLMrwvbATY3iIIifK9+Tm8UqVdSV0lt4
FQp6uFHBv5Spasi1peej23Rm6PXH/+mMqTgckCiIxt3F71HEToqI77hDWmysgCpIUxnPqv29vSWw
NEFEFXVKOZe1HelKdn8kQCjoD5XrrNMJqFllc07cJQcxS2rkj5ZP+HB2NxXnY+isKo+Z1qBJFbwS
+pwYnpqgrhEpEDpUqYuSzch1ZQsuC4Wmh/YU5k/flPankkNWWp2+9v6r8kXloNgnpkHSukl98exF
IGD/ogplgNMkpvSayEGTmHM0FxMjqMhfWjKcRxGhJmB+vuujnL1tVqR0dT0ztXXW0fRB+nXLQnD7
1Y4aUQDHVSS94QX1y+fZoiK4ShD4zP1MzqBweDCq+EjJ0WiWYNugj4k9KqI+QvE1YZ6BoHCLl37H
J3q98BZHYR8Lxa2pB7aFT9d9Dlzoc7HFP/9q8aknEcN3g2C1VqznfWP/fgscjVdyorEXQDuekO7p
bUME5OWmvp+dxynDPI4tYPOiyT0UZqcV8DSxo5kaP0q/JUi8y5ruCb1exDaHprKSHH+66YCwo6id
9R+bW/V2WAyAJnnr0e/HTJ8X3rI9vX+pttXVPwoa3B0BY3DiADiz4qVh2dr7CTQIXMh/wdt2gruf
HYFZAZT9jKtMYumlx+dQIIu8F/unrHP7vWcNLrAhFceda9mu5HltM6kW3q687hLc2gdBGo+1OBD8
O44ijyeHQmld9m5b85DRLuDFye1IAUIMU2pHJkFqQrvPLau2p0wn3BeC8Xpz64Mmwlq/4TD0OfkZ
XBEgnmCw9PIxlxgKw6tsRNazsueG0NwkJBg69Zm7ITZ9WloSmhdu4AEjOfDfNWs+qce1Y/9FwZ+1
5HcHXO8LmN67GbIMKymuTsoL32W6Tg69UAY+bTFmTKXx0THhljMsdqRIMAfvyuExMFa9Hv//OROv
ce2JxlszB8g/9FrXLiOSVCfay3TrtMwaskerwNOBepm0jbNWG3cN4CITiN1Xm5oH3QnkpQwT3woj
0tYCEvnvpd5u3T+sdmgPCaK6LrY3rP98T3ltBBzb13k0aEBXpay+lzcFntq0j/KFiAxw0DV+pFLZ
SSIyYFKfmtbg9DEQ0IvRAQb5eWGxkMziNuVO5QHat7F8b8/MawPLjGtUBu9krI82Hj5t0zD50eZj
Hips0IZV4y1sBGrsqnU5WLZmvogQr8cAxNFxZQcvvUkKD6CtXjtn22edxW9n9yMoNBjNP5qnoDVS
xTgLXRpsis8L063WT+xqNSQgYkEiU60vpo15T7rZ34VUCAx9WSeF4ZEcMiEK+khoE7UoMoHnfJ6v
zyrCIRoezvM2TLjaajWyqSthSbgXf7508Jlo72S0/HF9DD7bRVe1u/vKTBWoPQ0KbCbLS6JyDt4p
En2gwvsYtBh4m8YM/xoKYkTadWxC/7FGNN4IaJ6OKyeweLIcOiz2dK9mmXMyWeHLndc7MLKVP1pb
hxUWZ51nD7vCOp9HYqfrzdL2jfbWZ1UroDZXz+HYgThj3kROxoV8Fp3yXroCSkO799shTVjO5UDr
9VOVF8KFnXydVYFdn15XKxiPiaQYmgtQpKqoF9/S/o29ujQQ77OUOAgNaldejavGRggBsTY2Y1lF
ivRoGa5uU3wqEDRdhOWwfF+hWIblB/s69l3wWYCSsFUaZZ9p57no8f6ayZYhX1ZQXmCCuBqh1FnN
1xVknoCRAQuDHzKeygxaRH6B2IysTiPQAoaYglWMtB5zkc4lBWQ8mEvv2rF25pIfzp/finec8lAB
dq3PBKrj7M+QRsw+H40IInU4pAKRSF9o9Qducg8y8KLUUAaBL0Y6qD84HHrLg3cwee9Yy3x0Dbl2
SVAoJgIj2DZT59DqY8sMXAQdPpD5Dr0COPNEzB3djC68zBRZ6KHgmM0wYH/6RyhhXi97PcSF2onc
i0vVhX61tPNYrmJGwLtYDR5xzbUoV8Sc2/uwxUZSXbXjoyMhrXfUpucRoDYuQ2Vf1NFdUoVxPStj
GCXu1hcdECu00s5zQJd8ulsY9S0k1jHk/3hr9PD7SrGR+I3j7JBWibdqLkdSBG88RAG3SrwNXe+q
BJzouhEurBJNcQ0gGxfWTxkCVr+lroKl96YWYAlS2ukxcUv1D0iAiUF4cYr4oEOkZOjGSsWg3Y3K
0FOTLM6sVtSVLgtbsiIEsClNWFqTMGOj6sMzCREBTATgxsEMjmghmqpEVCMYR6FemuifN/n53sMk
CKyqvVo2hEExjHTeWeHLnWPrz6MOBWkipSzX9B6sgXIRwpm3+qX/2Cvzu8pXqrzjfzn/11bF9Krl
lBHdCoVeeaElVUP+aYpxU0rDzvuE3oFh2t2kXn4rFNn4LWP3lM0f2KBTkZUUsFYHaTU4B2WupGEA
8rVeG5kMKRa8YjcQ5omDQXqFMRIFrP/PXYZDzfJc9DaM+PL6lQfFDHM14QTZJeLK5efkAEUP+/0P
lvjo5iugfaBlWmH+jA8AWfLHx1own5aqJJdeLXn59xwXUNl9EoEvAhPfKzn4f3zuidYvG3ITrUNe
3jjj6TWWMp6JSP5br1IvqsEp9n75OmL3VCvyZ7QkYggJ0hf2c7uvRsRMIZs69XgX008GKrXA7brv
8OsAmgzvqUfz7oENE2db4e+ECE/FeE3UjeR65PwwzyAEDjPO0TdjKWjV7naCN8gMsH5n45Jbue7l
qBWg52tJhHgzPt6n2LgVP2vv32XUjFkE2iiilrZeY+cyjW9OD87ejot+9V903oQZKkkaCMU59GNs
H6A24Udn5FDhKI1ozRM2qdHywcoLxLCt7ldRfnzIyIPi6ps8B3AG09hoE6VoJDtZYmvhlJSBwaMO
zLKuc5GdafJztlRvG6dAxlp9Un3mCVqina698QIOM0X90Vr5Mz/0a5jplyYH7ZFtNCFA4efUA7JU
z3tYjAzR1atidCPxHj33qipAv7tYmqt0ZAhtB7QfZNrhnGG+7Xx+6ToAr3ro4P07apz4hwOVjbxU
T+7oetWzU1Byk36ce5aEa28hhdCLXJ5leX46AhYZZ5y44Zc0SxUhAfUBc9oXZvWEwSMbPEZQn4z0
AKsHG//O4lQTd+9mGeVoubJrgpSniREaOpwtZ2uTL3+6g2r6sr8EtXlpK8biJmP7lKUfvtn6xuT1
dHoZWA3jmRzht7wN6oWtYT7/PQwcbLH37NQopDBZNRr6QbHnWDmzKd08+ZDQXEmPLyqDDqw1j9Af
jgTuGHaxyKl/HjPmwrrvz56jc051JsLG8VktGwRb0CgKc3Hh9a5L8eWM9WQKav1N0mzjwLljA2S+
K9mlFPLRiiNGCggadDw2k4GNfEWLwdmRua41ELbNurP/aoMwdfTvYFTPifLt0JSraP0qPuxIMZLD
3mmDj1sbG/GX8IABSJ8oYsxcZQHAVitRj5fKvZChkOe8q6Ya3lCCxPFiecQwbBXwrBTEqMddJlSZ
Dpfeyo9aUOSLlpRRbwJE7BWSXnc8XvyawUggqA9rnAQ9ST0Gq5pnNBdGI5tLlHnA6JvU/wr9oNC3
LczZwMZcL5HpCrK5WQfe+tj7bsNNylo3Jdk5I5WDgPKU8eaEzC8Y5NO8EYBV8eWm7HDnG2J8TnuZ
eG3eUaVE0yWdixvAZERhwiMkqVVgV4qmLPTrkntC7+X39oQzEbOLgwBm685zohulDUl1u/y7cVJ2
yd2Joj1qG3kzF22JJaJA0DUU6GMgfBXAtK3yOshD9iCpTpoaNmJ7Tazzq5gCZgMhC/flokkJs/Nm
3x2Z/Q4Sp2yCEqdLrxo25SRQvIzBvX9P9Si/Oi0XIeKEDu0Noh5oA/S3kqOW2gl5Ilpsza13Mjqt
0rBLvc3wpD0t2wxeeYXJYIwRqpH4irXC52itajoly1fOM25dsFmCcSjCmn+xpYhBQq3cwRLB96t1
M2YSpUD/TvAm+5Nms/jq0sJDfc47bVYBGG6BPnPvDzDX4m0C5NNc6NBKDLcwjA2r3ZapMy0JWb78
o7RTTrkJ60KZNCShqPq9mIz/txcLL9v68CM7vwwwCHDhCUn0iNLXV7neog+gqZ+BdN8bD6NBjVDw
l1VmD3Z9jtAVQFZQavAD/Juod2I9HL6GB+Ol6qW2xN8dFrfKEkEHe/ftaqaXWzPrjdDfz5pvLP7Z
1+CzClztQVs35mAfqJ2L4YuU8FhhBNFK7xQkNNBntLoaxZxS53blVGDjZIWYIiU6xZpVOrbaGiuG
n05ZyKm6ROvQunRX75U6MvkrNDXCV7mP3QldXMNTcfTMtAmFF0Osc901x30IgaGNwvgNhraymvxm
vkfMy+IqYQ3UhqztGA8NVneaFgbMcN8ipUYRTz/EkBPngrO+p/V8T6vz8IvrqN8Rvxhx+Avr5NP9
EJwPysRb6teaHNcBfEZ60wlqZ8/Sx1snlWp0H2Q3p0gXJB7YoebUd5GJsK7cOR1VjlFKe0n5iykc
q9sxha4wUQzrZZPhxGtj4AfbYchO3sBxy6H1niP3VbPJfscfIKuhitaobvVj1CpChV10miTQDYHa
E+tAawWBTkbLmR3ZlaMdwEYxV2bCDWnjmTZAECW3y45RQoEz7+MBHOc5/X1c6ut6ZSKTWg57I/xd
caeEnZcaB+rSNtvj9mwxJy5xjvyFLIq3HWQHHw1LG44jptpuZR9X+TVFq4lYFtczaRojqbHwJHl9
Qm4ZGV9uLGjdkxQMchPAnL2e1yjMfiLOymWSN6uQLRKo6wNbOt+1O4nSKSPgmv4xLmrUsHBzCdul
wrIpcl25srsBxCWqkFYaPgTtvdQbZm0mdrQZyww+WjPLqvJk7+QKKHtdB5QptSC09xY8hiTgTiXY
MIi5lZetnmfPFW9U/ZRIenCl4a1G0cqm+pLI9RAPa83Ky1ppduVOkyKxdCtIOBdadFlL5lk2kBaJ
pr/t9z7cXhuZhB12cnhYsQ0QjIRyz5USBhu6JnlsXHZxOkfvN3y0m30us1r8PO7eFN20xgk3RXtt
21gxLIWkpUMGLmOna0u8tPHE11uhKimuAH5GeEwgqBOlRbboNrE1ER7YlDBHdoT3kTNsr4ICLAve
uUOeRba76P6ibCwZ3+ta2+IskDkdrqcZWuiNmvcSLq1RrbECYTnTQ8/weN5d8KHdbMvgygcTpK4B
8dKzEYA8FZHwWtH6lzqSXLbkVGsHDFZ/4Bw5jhxws+ElwcN8IUEzKXgK/WdZPMwbkBwsernVt6YV
A+vE5Q4NpPaRoAzf6TmW5/72cy04ztVYGYOxH74uhrqzQdM4R0WqL2nlCtrT0jaiDbS/AhUR18QG
ohMqWhJvQUk+bKpxO65wWWjEUY2zWdh4tLN6LMS752FPxmuXg/uy2r8haNxnIWHKJw5DZekuUo+P
Db2VImS+4s60hM5q6V2ESH7O1Zou7WxawbvmXAwxFyPttCZ946GXSemZd9ZqDxTaGuCI3y0rdGYa
tMYbkX7M3NuWlxaD6qhHONyY0xnG9sbeU4Mot2kEnlSCdt7YEBuE/iWV32DL5krXdqxmfw66OFfM
/BTvoSnGt8M8Q0X+VqiOoGUkcft2L/+izrYt4PQWWX2jJyVFtXv1ff/WVKT41kCE7+5A+SNye6wV
bmmZTrCh9kNZ2LpGjQgVxMqmC145nEihvFmH1m49WU7nnxDYM89+u8giLniK0+y1QKbQGsGcMm0y
420NNWontasWeM66zJ6Dih+8aFMiOk3QEocLULcq6lg/hMWzY6FQ5G1z5Zxin2RIjjdms40DoapD
tAh/igCP3Vb9aJJRwyEx10Cxl0f1Ni4Lau6uiKsInTK/lOWQlaOqiKWq6bqBDinWMqveXfdtY0u5
LBMFZLIGckqj7YaNBOUzkOEWO1/avOnx8dNG3kFDb8eO3T8+b/g9oa+0xbXURRGeVhD6nGbhYOym
3qtwqrQPVlOX/545j+32/crRloaIaNYqeWqtwl+oY+9yxfA4ZbanZanoHBh+Obh/0H1Jm7dieTtJ
KjxzwKxCQsJWwqWeNnnG/olLgtLpng9ZzPvZO2W8z+Bwu/FmDRU1s0sMPd+l2ENFKJ+3o2oGjpU4
EOyRB+i9kSU/MJvAg76saNJC2eYWei6kEjB6xontlfka7N4bxdNk1r161rXYrW8cDj40UegeiyTp
3Pk5LU2t+3nUf87XG5JRD7Dcan6c53ebYSfghxNlTvHWJ0Q/dVkA+tnFQwqyQk9liB6mMe9CwVYH
Z1KZACDS/3qHljUwnPl5gjC26KBAKGfVZHYaYMiQ4d8aqjus+FkRq431aVrlJ8gTuIiKRBNh3QQH
wrmclPNudEVkw3EZakRenv2voyCh9DjoTcAhdpVoHzWSM8TMmsKdrP6MKe4E5UqgwbBT/jycQo1i
ftHU/5PUQ00JdXIH+gOKWEhq+U4oEEYmmqLRQysuOArO5xAaZK0IEEcuBTRnuzHun0rtYvDpddnd
PCE1ZU12QNkR0TKlYk07kwqmPJVVTeV8ONC8xWWIBrO8EM0PoHitqdq2OD2pBK4TsiIqh/CfBegw
TcpOCh4fIRfwUBgF6qNCOd+JnoWzzQyGsqpLMNiFRa7e+f98WoGranRsP+TzoU3FZUtkLsik5CVd
YgVbFuvw+B5qbzKC1OPfuwMVokJk6ZIovX2QOHczsFCHcTzE8KNMfdfTbdCCKCxR3rWxZ+FF5Pho
A7iInqY34erMBrl4B7URAKJc/VOQvhkcYdxqFY5Df8Sbfg5pLdo2uU0okiFKNW53RWqs0wgadbZ6
kcHLi/uPpogDNXWZema6JexHpz32BKCLC+Q850DcdelxRy2zqTethzpM6V0+q8ymcAo7oxtN8inp
vSIV1PNafs4ulLkymuiNnpwOfNC7HUNlCCivOnOt52nPoazqathsVzIoFSgDKAGD9WskrSjHmEPL
SU58NTaXNDnV5IczuZGT4V7K17qagjV3F9q+HpIfOyysl5R2ugYeuDz6wPxH4CcCEF0e4etpeoRs
7OxC2OqWyES9asEov11xEO5v6UIwnDE64zlvBHIy6PJ/mlZg4hqVJkZCdaN5/jv73+Mz1k9Ci3VW
LAhDYoVtZJEcwk8P79VtarSvzBY7HkrIxiStoTq561o7857X76Ii+oSQEgttwrEq5dMQgZ65LodQ
FzVzr2XdeAQm10yofIkvwgkzRIQmpzYbXPyiBlHCdFREQKzwmISVcPW+rVgaGgPPvbdLGaoCdfCO
jOU+zp7DtHCveCYBcVSEu5pWJdL+yggffugpHrswfJ/8SBWzIM3NFUpHo7kxbbBdX62cLTxO3pj0
Idff1SEN4oXY+Zkz3y1BwGtA4pyBB6iwAa2Xt7GUSGrsWKd0nCpI5BsEBiL0Xy6MMGR112Iszop4
r8f3v/B3cbFWCt93Uwwt94ro36qbox8Q1vqN0CChZFqajOFay8IX9VtiXqFYTNF94k2gxbrkf9Lc
QsIo4lViq1Y5ApRbWiezgo0ZeNPAN2wWeY9b3pKAVbKHvloaP41dg84VA3TKt4fcv4U384duYk/H
hpLTv2QZxvY9FviA0X5L4I/r75gzYMA0Tj8OkOqc6ee15/8RXtLfT+PRxmRCc8eA2oypB19jGiPB
VHD1DuzVjYgtFnPazk1sHW3avoWh+w6DiQRAeHZu54PTIsZC16mA1vOgt/MyeJN/arxOCAYOnE4O
WqKncABqD1gbLyejPur8CP/JJzFpXElu3MztnqSrQ7/xo/99sRwX73SLfxnr/m7dEMNXxFgQF5zs
5b9cznWnb6dbmjR9zaEJm/CYBzJ67LjpU9iDYk4rYzDpGrq51ew79NnM9ldMDi+fVZrek/dd1cSq
fpCsdwwMCo/G7PjnbuzliLSqV7lhklfX8EDKbmvzsdLvmP5A21CjdxVnbMWYn6eO6UR2DHt6iNB+
NIacD6AN3tPVxI/McG4xhUBOuILUzicAAkW1LQqAYgC0IaQSlnr/MlHB2LZ9CNBxJ1C1pm3323k6
vkhAiEQgFwgN6n4Pku1nDQ3KTYfNEQcfppDbldKtst+d3Kw+MhRLwkI4YP1MRbT4UAbKOG9BwQNy
nL6+83i38Eh2utF1WizgYjx0YZ89nxupOu2FdyJflGZmWUpOGScMM2BJVwjDuxlIcYYDPVG6t9EC
+3BVoXuFBJe5wG3Vk+UzXdodE4kJ3ge5KWjRJKuXo0tA7t8B90SZDnH8ePluIjIBo2BgZ59r3ulA
CxkajO46KiRAf5R7X/xVt43kYrCWKn044G60gIR0l0xWWqL77hNdJrDniDZe4zky6RJXnf35k6cn
RcYMwcjwhiFurucaVDxMWmkbk6uA2tgSf509MY1zlG5o7PXi2PSJvJeh3u1YbC/cnPKU+WTEZlSe
m08EIqgJL03dpYu3CM9X6PUWWajs8OGM74RWsgjzgSljv6W6woG4Q8mbnTKcalNi+JFvFLZMy2nB
YMLizF6sl2IgrzNY8LJHJnqk0GTjcoNLLdGkFoPKCoR6esgzC4nYiAZRn7J7JaqRA6zCyioVyQwF
Z9/JCyjopUEIM5Xy73rY2rPNybHEMVSALn+Rrq52q8v9xS0Ev6TeO0Fjr59lehhdwV15RI73OvWB
5J6TxE3FE8tRvYXqK3b5RdkncDOtyJu9MfEyCahHrXeMdVp1TBbTKlHzgtDbB/YNTMt1NUyIE6kX
/+VNGq7uAI6makDhsMI2AEZArjVCBszLjWVrB/jRlbQPw4AP/vuGG9/B7FIF9/x3+MRyRjH9MGXH
bDudYYCmpuFqkfXS44jdeXAEHekif/PCdaGijpjZTRXu6kU0XL/wQy+lZ+SwYwrJv0YEE00c0S2Y
giFkJgpJ6OG3ciSDaYZZptbx/2wPTy1RahfJL3B5I0aHX1dG7CH/c6jrc/gk4k53hiCQdq/LPqip
+e1QzzOxIbHlBstp2jHY2FXpP8pvM3tmKTxAtx7jqClZNnz9GzRTwd2YAk4Hc9UXCW4Auyd+BVPN
MmBbxq1osvQRjlz/J5rEq10vchtr8g2+DrJTd1WMlGq6k0Ht56Vx6jR7POu39ojxmPnBY70O7Mun
taPB/it6LvfgIk/SR7+O9zO0U1TF6PK8NNYKyuLKypPDC6ngaVpa/zsiDxkMX7CQds36YuEY/yUp
MAF34JM6S+rPBIC66uzDLOKU8OKZK8Mz3IDZKPc14umxGfrNbVUcr/djQZ5oidq2MJIKU/skNTX9
eLvAXEENB2/1T3B+7+k75Ul14OSy0lbM9e61YSRgao1XQC/st07w0thb8/XmKqs8CtDOCqPrH63S
Q+EFwMT+cW29s66rwvDIVpdSh1Bq6kZY22GCpcKpI3vxqPZiL2T9rLYL5z2AvqZk4YnRraKYNcR5
9vZBx0mufofGDi8Cvi7Bz8ggPMDqAF/D8GssmqaO2d8iao1/ppl3NxSWRq24Ixaa9zQx7cJTpXBj
RfyQg7UXt9C2Cb9cfYmrPTjOuqbkTXvlWEITiDbzXmYeet+WtxmZjfpxOzjMhuog6EnwZgVGH2fG
yKBQCZhuYOo8ArgWK4dHvvCs73zRc2PW8qJ8qGAWtUPoz30HOPoPPow5BSNVF4FFUkcLeyik8SIr
PPvLx7amIGHkYa5a79ixf42kBYS+yVK0z1bTJgrvXYGoZnIPj3FBD4FbyfH2/ewfhg1dF/ZLWnsj
Wf0Od8eZAuARD5qgddBJvHqxMBw8dsAYY0kxEudY66xfGcz4FFBX9b7M+QpA2lA9odteWtBiq0u2
YBWMW6JLbPU+imddfhP37UaCxFSUB0aofsmN7DYaeDu7RjPs+oFiIVsRvUBlIr9imrOBbVhO4CF7
RK9ggVuMP43njL8fJ7SeH0MIUeWHpWsmQOWCBTHANbAOS7eF+Sa38ZBfLgYunqghBrh+vKxPXzBC
YpR/Kj3XkMkKGIi3SXCgbdeFnQgXtKpLQHaRH33hug5+7uw3kD0yGxvH7cuWFldtQob+1n2KNTk5
yJGuNKjijXAEDS511gZlKI1+JCjzTNUPaNG5Owkxct9EYSB6JJrcj/dvxwWfpgScy3VAppayn4ZW
qEWHn9K2C9ZmDUnhNtABoHtJMJJmtXKzoILVvxmA2RN9BnNk9IDnTVC0RXfqJgHl9b7FogLaVZZo
q8+JmkR0cdhqk9icQtNQSSSg97nMkkgXidcUTKvJjUgB92ODp27/8bympoANxObumRmx3rpnE983
2SqyTI1dgLzP9zh8O2+SrAVkjqSikeq24nBCeBGkZ0AdT8/N3n2TordHLtX+4xCtFYJhYmR+r0PD
P6A+nL2XoftRcPTzdpBLEBOYRLD7iMC5HElFkG+w+HE3VZ9k34r8YLfxGZUrTLzKY0k6PI8enkKn
nyYhYRyQ29SBkC+QsC3PNOzSUKqXgtnuDHURKftKfpfIizxvW00tBSbRfjka1fqbAsypPl4uwh0R
ZXmolC3EQtq6KcWgJ16UXpwBDum/ZvNC+6aqJqFfOa/pcIGzj6Y5jV6YX3CbgtKC4R2IHhKTAWUu
ZeB9zUTPJM53hvCE9dRPgZ79cvR+9Gu3UXcRLf4vVBskFcfjGPzexz0GGOycyx78EMlvCRDTpZtp
W5amTAKuJGV+Zu/bmR6XfxtkDRWb2wHptvu10YT6YQ6RhbpFMRiQ+YdhbnCfV0S/54YNRxm8ZY38
bkk3VDAbbSE7qQfSrB9zU0jpekzxoEDdZIrY7B+Z9Nm3lSi6dvTr0jlCphS64v3dvjH1Nx6BsH8w
ALoieNb29zFwImMvi/xizGo6bxBU2rPhLFp0AKbasv8p2b3WFXQrEYJzonXCNmKz1IZjnZd6mF+W
IavdRObVtNuHZ5hRhq6hRIIAc6Z/YZzn5i5dyXm7tlS0edw3CJx7RgrxB3+L5VrAZqITECijBigi
WVcMaKFwb+fDcnqufojNYhWylhz9Eb8HtZioMqP5PqephVURhJBcWdiGJMP58dBZEkdiZLBvM3Hn
jXNsJ/pXlU9AW5B29j//RKn6b5DjMI9EIAP8ZSU/dzxVKeYYqbtqRYv0xjMmMc1myj2adoJF2nFK
Usu4l/VxMZoMkcOCvgIYfmzUaonpFJ3Af95h/HvJYZmYUerfCpVtEJeNbCEP6ublavPbn9CKPGRb
BRkYYIdd0VcxVX4LG+14EcKKuyBGL92U04LkcEXYBZfDGkEQ4UK6nH9W8nyLcPlEsgh6IU4ZEboX
A1g1rTz0UQP1oAz3otZoYCY1EeN7YjSe40Rbx16DXt+pdwKrtff6q1dpMscDgYCKGEOjSdijA6ZI
5SoaAd35+6TPitor0qNIIHlH8LxCK3p9hdxR0curghHQJ8hhVXFNyJthgsVCIBiuQkLwqw9w8qt/
YVvyDJc7mMPcO9lNX5i+SZt5pmNie/Zxnc9UsDvNCF/Ypj2Oypn1YO1L1wYc+rNxy0HyBVMDrTef
dOwguOzwVte6qTsgtIJvVObGls2YR2POGjW+CsgVxq5IawXxqOuholl/U5jFQbs5Kt/LTORgrpXe
EBQzECiSbUbIiwx3b6gpxf4JcFPu7BalIUVzrZynyw+TXWF83Qsr9hqZlrbyOyEg30131tPNOPj7
2DlXOij5i18ETrpMff58sTLebUkIP6IAUcCD2Cg111auDbaMvkdqs0X3Sat8w6D1t5+B9ZCC7fPm
sXsiot31i47O0Ej6gdyM54kep4ZqSjR7d2x6l3uFf35oFwQ1EYaxN5vL+ZiU2wHPMzMONtNXnJMY
s6Sh87WDKo9s5V6+AylhT0fXcU5ZstsvpY4uOGtQPbHrs8r8wvGPKIp5r/SNVx980TPeSrv0S4v3
XcC0cIXElJbySzXuop3VzJgTmToTGKtHQnSXqLBmKjfqZPwcHTfqSBym1LlgSJfAShftUBCDhGBw
rlM/wa/hPedC3LJLtrpFZAzNoOkme1u9OSWuRMhc7UYCOg3xUUikZ3YmwOR76hjlTEy61iI12/U2
2yGOm6nm9MN1VWIx5qOi0O5JzTPuRmv8F4Ip5/rJN/k0eX3UsKK0O/NDXrQ0Gvb0mAHzPEWy7ZWp
lXuXXZCew6KCi47yk/qLv/3udXkKHN3sTmnpP4ngFeTGyLySof+TuItM2QYZNDVHftg40QEisy97
NwPe41dFIuwxRY7IPpD23GeWugoU6m04elDahg/hjj4X0ZjTlEypi6fnPAslrNmpbzx7h8isF5bQ
Tm9q1bBCC4X318+mGMIyrGE/pq/GpGeyctHXEq8hJIXLNRWInl/V5x0+EKcqG7qbqoYjaxp+g1PC
acJ9TqgoOEOOsJwUaxAt1x4ikwXCTuCznxQuFje/JsKOKXorLjIun5oJoAWn5JzKdrCyysjIdK4o
+neVdOEYyycqkT+5q8ZXOtHfCEbk4uPm8kLWCuceo+WrYAcd9DLQUIyxJG3ou8Xh9s2xTYgLtA8T
hYkh+MSB32it6GCw5oLsXxOAultMJoXR0sok+rpcIBZRrS5tCSGqbQjJlGAA/BLzLDTxNkeRUYgX
Zs591CtwwoOk6cVe+JOvSbk+ED0aObL1HnB/EZLKzHXL6Hx98cU7QwwQ7ZettFYuuKFPRIFyQOtw
WJOh9SaujePzJq+OUqk9qJcOxqCdgsf+wpBeNEZtC7IXFTG8hwLH9sjXkWQn/vShyc70c4OxPECA
VrpUkU98EAR9ch01CDVsNjl6BQjWhqVhvbaLYeWT3v57MjQTjYbMNJjx9nh4qt4ZJZ+Ap2FZV7on
H8A/OKuoDT3FeZYvrZfTzcJxxXcenjcz/MVBWpLhQa7boJeXgDeftWH2DiOaresqig7hmcKov3V5
li0x710XdqH5MBc14q5BhhAZtkwH4oFzqvBfo9QP00azbxDKGQ6Tk8JmZgtyNvNkRKCCkxfYyJeu
yOFCoxvVZSe9Z4inp4klquucti+vR9ViyqToXz/YzxIxOewbzMveE9KeCbLYCEnXbP2CGvi603SE
SfEaYvUTTgGpe5CnamKQXuCiZfhGOluiq82yKNLDZaf/mnSRGVioYQwPBJY0HYS9ewOtWeWFmn+v
3rs6T6vXDBB2RaQ1afp7gbLytfoN20el0tFpY9ijfkb4WEtmjxZ6SCnyr7dGqFe7ER8vIaoV8YvD
nr20rqJ5lCMKa/cIm4I6doky/l1fFhWdvxJHvZILBQ+1k8J3IoTltsYH+xPnWSVb1Bc/q6tT2jhm
QSZCF0fTbgRPC+HCSLWNjkNwXwLp957DRu6sPE8MFMoebcodlS8BRw0K66ahyRb7YgZI5HsgEwxi
aJySXGPpVc2pFBuZiPxphOSeeB2TFE/LcU0n26V9w5UPflItA94HmHaz93FrgNwloriaBgDYaSc6
LqdonFt89wW8uBYmk2CztYA0QHiGVi5srLjwim1+vXQ0riA1lxYCevxfmTEqkp4TFlOpvV7uVz+6
+EJNKPoBEkGc47+ZTEvsP1Km5R4zzPDP9b+aN4POTnaKJPbDaT7QpgM0PnFN2A//iB6Y65DedOj+
vkmfzhKspH49HtAlWH37LKJT1aZwr0Gj5GtaY5wWVUFIhyWJKNhQnJh0MDqszX+yolpXaVumkiZ/
6gpcZf2jMo/BHePpPc/VJMDUsr6sM0VRV2v/G8xFu1WvYN3U5ZQ/beDy3frPe1k4DZsbfh1t/Wwq
8WCabMd4l6VCDtrCineYwm0LhOZmy7zAZQpaI4GsnCRRDfvAkIaO3Fpu3S7J70xeR4mwk7OWQiRa
VsGgCLcIUAVMbPoCEjzFXDKExPN2LBj8kx4LGO8HevhZtjJ1KWTK50KXqHL4GE6cv0KId2sgcgCz
jVgKkeHFjvDxegZ672s/oZhxfoziu7goLZd3gii+5DmEHA+v/wmwpDPIDpE/Dcac+mGt9+dWRXvm
BxkDGnse4pb1YFXWEqaYwm+X3AAn671dhYJEDGQYXAdv7AkmjKMwrS2OEw2eD9cnZ8YfQrxceesi
kHBSvPI9E0UxxK8AImlZWF4JIRIVJ+SCUqQIHXWLbFEEDOJbrAVRCbmwuK+r9UXn+8XvPTFZQTj1
b19r4rot6DgcKa5VrdFPv8zEc83s0r7n5MTKFTfyE8gBSshNr/HTTEjoevRiVq7Oo+b5qYEyXWby
T59FVvxnzvtBa+1PVbqmt5K38PlugWlwnB3YJ7auzglm0N27gFnEQpxB2IYu0KKZRMJ7LwEqjr/k
8UfdmGvP5vtK8cJjUDGtV67mfiGLXN7EbiASwQyuTSKxprPJ10LEyPZsUE0tlp1k85AIRZYfqmhq
htnIQsuPMfSgM1b2/hETszE55vD5wqgIbiF1YFbw/1NZUsOLBp9bg9EHBVx2e7aWUMsC5WydgY1t
/PN5x/jjQCedZEzbDC0CsMqjYahEIyXnjS2+pzfqeHbXoyogFeuiAosXFhsifXo+z7tclOIp1/Ia
FVvgqTZUlVR4YVEWLdjijxosEwp7xjUBX2YFpY07XNF5z/IDYdmdt3M42+wdyhrwUTYjWqqmqJZR
Bp7p+9HjvetUt11fI+kzmIBuD885gPE7zo8NcihjUB0TD6kv+WANeJUXdQYhuB99QeTkNfIEywxE
XTO8SGRHNYZ1ATvhg2HPw79OhiYXZGhzwTgbMd4fmRJyFLhqQmo8iHZOvxIVvGw/lf47AQQaUb8q
fwOmE24t3qrQOv4pP+L/h9Oei3hI8l6yUdWcN//JiOhGPo0DnM0BAXpS/Qa7IzsiCZI8w/Kxx80Q
q8lhCzgKNhhqyHhAiSica0cl6XWk49cTiWpRUCK3IUc/JaLUEXiCfVxCpR5ELs4RVf8jdgg6CZNU
kf0sU3gFgbyzxokrWsjFZL20GcCz54vyI6KINCuT6QT8XoH+EYd+g3vlxD7sYcIWEQTT2YodUD5Z
L2fVaUBM7M/Y502AUYj+uDfocD2usKZNNwG12bZv0lyCzWwjNxxdlZDB7hkICx8KtifozK7O3K1u
Qf/LxHEnPmZ+uaLc65UKwDTnuJ2P1tSXkSSEm44Mw8lfZgA4+PbVYSSTRzwsZquhmrOtPS6Fy4fF
q4xBxEA7J/wwzT+V3Q5PElagCSkEupG/6eKaf7rf2k/Y8ylC9zD39ey85W2CQvg5T+UCdIjERbtR
tAYPFSWgRbPPEOVB3VVOlyU0EY+26+6QA+rU+dUdEjI59OVPAmWna+bhBSxPJRnsyQHu9t6pWBEt
qaIkfKvduR/+mDGgj29m87YX2Ga/1Qn8vI88bkaMo12CG5yIP0i1m1jv1UFL/dXAEofh06gtKXLP
1ag8AvSefhZy2NZ/MKXEqzoEBuejmV3AvtEC0ELva+SHIiR+fUHsE2gBdbCRorLjZmGJ04wFemTH
duFRMsJ1w++6kExo1ZGcf+4+6u8nExqjNMuMkoOM5v6JYTNjesYF8JKqH6zTmHvwHVRzb7fSlmSh
9NAhFHdGOlfG5gQcEY34+XkPsmLYlCFetRqCUFmS7lzvJzttvzQCwMCeyOW9Jik56JB/dDgGcMMh
ZjMJUsGRD5kH9S8EyGj+Kcgm5PkRA8dJHqAZV4FO467LGJ5yns8Qn8l7k71HwZkUzmqG/k1dTBx5
21p6SfW2o9f3Rs9uY+sx1/sHjh8C9WoJy+kQV9vk5YfsRa++0NG7b9phkNeIoSaFXLWHLGAHByhy
9nJywjgUi99hgCLdl84HLdK2RecFvf57UVSB8LdrkiAedbGlWbzRyv0ETZuMyfAsDdB2QEu4aD31
37QNr616tdvTx+qr1+lqnI/CiK6SpWUNuYFcebHax9IFVx7+MGep7tHomug5ONs1by5F700rsfSr
0UVZq+U4d3spt94qHFc9nJ8oVMsENJal2v5oyyK49mZ+LYu7kuMgHuRPEqegzptuxrzA3NiLSaZz
ULKLjfEKih33We/C74nloEL6TKm2fdId1iLuYFxJkC0k2MPDX0l7XiaZCmJRCt5X7rXXta4HjJRe
1ENrY9aScUo/9ONG3InRmDFnnO21a1lNV6dgieL/JDs5Z7zDBc7SqJXtThL2OlexUsbJFtzSCnX/
Ryaq8W5tjayqdAH2yCXEyL3/5QfjUkDfTiJE+q2oQyT7W3+1eRy6bvvl8J3YcCALyIFTIP81XK3u
A9WyRJp2w7jXKlDeMZUuMxExeSwRmjYWNrq1d5OPnwF6wKdxtLcQGxHevY4yC+kDKysRjGv273Ap
Ap4RAYjI6+i/Kkm4zT/O7xqG3IKur9fQnb1ZBU8WolY9L1gsNlXioffOAsm8apJIiHO6xVpC03xk
LBPL3o+zPG/kNqYvTVC26C8uWDvU23DMAArHvxDdBLQoJattp8xeGTNMR1BjEESrK2S0F3hXYQSh
JTPcIp44AroRSXZoHe8QXTLqvwvumo64DKGTybSMCTsNPuKtwULq7V7edIGe3HITM0wcmkZNOCcc
DgMZgdYiMPmb+KLpdMd0LzIFH1BbQgpnqbc7tCPGxIgreEDfKB72Xnqisty10jOnPSaJzpAbz+AH
+bZddc3lRIDanUtfiOL7I410Ow0XuXwcicpfbdOwH4CIm+sQg4V6xX32rb4BC8l/R3cWEhSB51AA
caG43y6tHg1D+qcx+fq+1XmmIiOoBGopcqO6qT2NR2yNujWRVbGDLEz8zQ5hIVyAhYXpMz5RIGW0
Ff03gdDTZs3ci1T06r7BCqYAc06MrVA2knU7uMDFlQLek02TO60qP5TVvYXEPYwRBhG7Bwv2tR0z
1tBpp35Sqagsax9ZbVmItEvk5haJIXTTnih5CzAv4m4BrQTsGodXknCDhXgNatLS1EMkymUFUiFu
wSSGk8MeVOnXc/U4/c0xxhkuwkiC5YujxHET2/CCkfMrCzrOtxbBFo3NcUvWhsW8wWjKLRxw6Tog
4z/k6+Gfb1s6Trk/N3lLZZXtohr1sjgt/+LTQlgBVl+4XKP1EWt2EGS32K79ozWnbQQoeW0AwyIV
Jp2h37Fm4CgBqGurbQv5NzTivK74BQ29PTSbPUiFbEX+iJioeiPh8lvRKUM8tspDUXGBFDff3yVY
OJZFZa7j8kQNd90rzPH1HV9+8BjiQFjiwau92/MiqgVPmOVx5G5yjm9DXcSXqEr4h7OlSxKq9Xgi
9nTwDjOP+Yjd8ZAsYJLYc21JXtSpkf9mKDTcd8CeeRHY5n5DCrzawcrmL3jP1iuBClpl1vsq65N0
uqdcoG322z4tQDYLzELTx/4X6KPuYNoCx6u4u93SvrIxDIazBbFBNMpa28Z5oziFTApivVwmoCOY
+lOPIEqlpB0xs8/bd6DcGVEbrVoROvt+uwNM4TAHuWY7e/BdAjAVGaRNLobTPpF1EYW9OsdHdhZx
Ds7ZMLNR8E1r3uzO2LTpdB4c+hdzuALXLoCNvVhvRiot8SiGMdiladd5OzpZJqBw0ZBnhyMbwUry
X7xwhksc0kl+VxEA3cNc4yyemgLo6vRdzFlllNBWfHheIttGAdPP7x+ttxjwtmsW01rA3PjgMtOu
woyGdmAs59LDfZu0VGgYLOpS1GHUvESpZfeYrrT5f4cxJG6rh5Y998z2uQRGIzDvH5LaKQZDuYoR
ehFlp+mjE9CzBXSJNXwwPVZxhGRi7coyYqRGSLhk7l9gSNAF3GkzMJAyd7Tg6rmfk3uUriCruNWZ
HAJeaoIQhF4dQXcaitIXG0C1B4kiKulz7nezWZeocOKo8UtDSgn+HUFIv1e5gYouw6sMSZlQg0j3
aNnFFMiytHEar9GER2ZrAUJ1HE1HQ1A8kYVUiuzyqbSdo11nnchmrnUyuYn41GNEeMGNzfngCTS5
mHmf3l1z3QxxKhiYw4v48cqYLNiKm6BUoOXypYeW0ryC/kyP8ywfDiXrJgbS8GyRidvAjiyoNWkF
4dEXJt2qtQ/5ExXx5d3BoNbAAk60TJhY4zBsL91QjeHB5YjAcMu/0RbqW6yKBVzOFMUYqriwLMS8
GT2oyyOCnXClq3pJunVaCn/KBEKkj2HrsDn/ghw756CYZ6OwoM3gOeEujAE+70yUQwo6Ly6pTp5r
IiNfhVAm0ME5tBkXXW8AyUdMcH1+cLSZche+UFF0v8/z+TmZTIFcfdNVSbehx9ruJHlC//cTMTIn
EIiDVN6fKWRCm4oqVxZdBEfghDwcFdzb83BO+wdjWrJD7uZlB7ffVzi6bmhNuRPjwOE7xE9orJ03
INKn+RwZ6jU5Ki09HovkHuupgDyIZjsLNYipeWlnGHfZdjHyVySDAQPE64oSbu7rnuxUWz7WpM2M
9o8KVKDFE2GKiNkoBhMM7C9DmOpLNwvprLoBODnW07c70MGLUOxUYfsgh7sizXezf3ViE/AfjEyt
5ggmpiG2ZH1z59yQBmqkxsqGCDZ7Z6gMVkNS7xHeOVyG01G+6YMVG7HoIUOehoKaUjGbwWXqcYF8
BW3JZG1t7Xb2n1eByu8LtaLORg7eTApuuoSSqmkGyLQCUZU3CCimgN1H2TPAta7HOK2Q7RC7ELTM
l3jHImjndl0d3q1wtHBPIO4wgwcKM+0G85zhW9mJe3ixEpxmblD/Yznot74U2l5IvS2LNDKPfhO9
xnDljVLbI+BENLjycXsoXVZ7FiefVgu46oH1eNNxiv0FzVRs78P79mfvNxu3rija/q05ecR6f3IB
FISb2eQuXB+1wku93fa/OlCDkUfPWK89MQTqMRsSmzZSgtKrOhG87XkrDv238rFeeJBaI2aXSgAS
hSL5OFg8cuPoSjTYYfRtP0oCvbXbfFbz2vAQTDogRrXtqlZLqP2Y47iN5UkEpMXf+22nEyOOfLId
NWyioNe9KzITOztGPgwveORLyFgRFjUK/EBgMFJbQYkqtCJ932FyGdAkhr+kIZf3EUgYJPhcIvwl
w1UsgcVdKbR1Puk9+URRVkjL2amgrd04mAW5Uw85cRblnACkF8KASNMZnEVROyB+YELYEvB+eLXa
en8OZmQISOe6dldku5NyjhsssWf0mdOw1lNQaAFgWyA6UsE4JtIAJGEgbRmxStfbz3oyWK1JJc3G
iohgXWRSwiSnyvqdjpAIYgdXfITjJM7eUH2xtUQlBfWtPXdavyHCrtprshNLthVoFL81CIaT35RN
WnwKRWKNL0HG+GQG7ROoYu7ZREh6KyUWsFXiLNgX3oc/0SYXO4fAhhZah+zUzRknZcq5OmNQrg4f
b43f4Q+cnJftudMqt03jZzfhJrYZpc5PQe8ITVp2XrC5AG8MBAWCV97xjJydO3Kg7WHsOUz5uYV5
7EK6onz1vEbg8ShSZuyf/HGVkmBqgsVLd5gfoF2DENdcQlQqiblirW8067AFcB2Q5f9erPODJ/Au
iqSCDJglzWjpe+jlvXny24g5WLrkm3uYX3B2SJIADzJq/v6rWQJFZ5PXCCdoBajv07KtcKDX4d7s
r1l0llEWzF5l0j3Dfmn9IGUEBAd4ZUZriHKrIeE3IATplhS+ruvsv56x9Hpa2xNeMA4FNaEheOsw
CtHvFIHkHMr3VgZp96fGf8HlWOND40xhfOn7op4CdumD4CbWGP6FTvIeDztDdHu6jtcpmLi3a5Oe
8+r0AuA/IEtbPXSUgqMSw4ZfkvOElVqqt8Np2W1JI5o3FKB7DnVS28e/4tFoSseQwqkZ6+Xyrepm
18WIzAjpjkpXwHkHb3Vn0Tq4pSWzgfhn9wX/eTPmPHy4xWAuDhkLIf+bGJBMmz9BBdJX67bfa0BX
uTO1ZRNesopE28s9Lu81OM+HfJDKTGvboyGQHOj+QLj4L/hvKS5TCSNHLQNMvrOvCslWi5QCTaxI
sHM1S8II9g/IhjGoMZgxENZF7Usx4EDBUY67prUGZ3ZWQDjaOLam+OxuJEcl/bucZCSOWms8nvSE
lU4NifCV5R1TMc8JM7wXnWgw88Vu1jmEtW4uiK9fGVLLLNlxE0+SyQY6bxWafZ9knaAdx+IEEFaT
Karc2I1kl+RQwiVk9rFbbbQzGu6zplLAwGCuiin9z0dmMfmV556gN6bjEfNd2EpleJydzfjFwN8M
GxXflzMti7OUz/5AhDv6+KAXwiUrRePLS7VIDIhetqEDrtKmZoHPJKZAITnRXLoVmCSV/juCQ/32
1MJWVnNRsC6zkMThJylKAqlEOZGYpwYqPkGwML5HR9p2hwQMrdupk5aE6etrQdd0QXWYn3p1kZTr
4+nkZa97lw0KH3llEew6hrfypKYRgd3eDA2ZQABDAC2YCIMc6UcC4UDXbdPprfqJ4pymowj/jGFf
b1+44Jq9VH4HJxEKJVUWkYdyUMqAFEvAT2wLqeXq7scHM7FLRAGWM47ZxXwDr0zzOOHKydBiEtq+
Vql1Ezi74BbeINAznYMWdmqgirL7+Eg2cFP7O8ucQfiLlNsIhtgMqly1Iy+Xs/kg0vuOERQIxdAY
81T//psLFd5VGVKa5wTP4V6aMP8gTNcaQ/r982wHueibXCwWSF19zSub160zst0EVfbrhhwCLsr0
u9GU+4fqCyZF2DHL8f1wSNT9HAUuyDvp8uwEdFMXtLDg6/eYPuVcsoLo4gnoJwIgAxwMcrfa4Okz
zQy0kqgxP34pTZE9m010wMq98n8aLoiLXwyV3/EIbWgj6h+XHwAZtipqJj03AQxzt+AdjdU5tyJl
8tZRsgPU1tOj1puaMDNjaMm+27U9QaiSW+cp/dGNOAI70HE/JL49d0CA/+lhT4mm8MqomkkvrVGi
kIAEJg3oliBoSRlLdyoCDMfvviHuDFIkfLwtMwXp9nKz95NfMNtuTQ3fY1XyWCu85zoZwFFYxpUU
3cvNpmFJQN1JD3QF/hdLPHMTA82YLYzHI7ipURAW5adfgLf55Vdiyd5jvgWFwOnYnMWO5Rz4/1PI
ALhZMJLKVpAquJbzaL8OfnRVOj2kJjr5fZtw+WPj43A4zikYU+utlIhsas5GADIcrPqe3Oy+9zSF
tQ0xCpgkUmmKdyBvjiXlAMhMBB/205jgJabxZ2qBg1gLsytPooZecLE1eqoBw574qGT/GIXX1TR6
aojYnLMElf2y4BOaHzcrpJA0/BLccekQ9B21pRfqA4JRiqYmlgMQ6mq6BJxthhvgFQaCQkkh53pM
Vtvqk8ddRTRxanebWRJt/KkLJzQvXe8xPeML72S1QKKCKRaBeNAc+o2XynGesebGy01YUzARU48f
U8hw6jwEfMaRRoBL1DleKpKSC3pIqKK3JiCxjKZc2inI7DGY3CwJOt7+m7LekWcC4yFuQkCryidX
c6OzlSwNsrFooGQ2I4i1XvOdwW9BH0tnSMenVVaHp2ExkjxYwrE4DOztf2n7DAlk+vf8ff56AC/E
Ui5PHh3GjJXf7rDK5YrUeJzYbV6bfxUg6RxN7zEayCc3MMUoFjayeCnHErOKlBzrcOHaPwnHG6pK
NZPMFJi4LYx6Bcn8U6MX2LeAkK1q5IW6u/c6VaUlzmGBkNd9FUGWvOnaFrWmzTUsZQleGsJYd6YC
uDfEk5vnE2CYT6aHr8oRpDJYL4UqGroOnUH38TwwdNIetTDCcVa6APTGF/QHtm63vOKtAhlCvoT4
DAHuROCnA6Jj+7KZnIt/rk/lNF1aeC8Z4R0hOvSu+2HiwQeOK4weLmP2YMdyYP9wnRpSKHD65irU
mQhLUemusfbSUc49zKGSK4b/McxVQuxWFCTqYK4/iPog3XefZL84WdsJ4eppeUQX62RSxKUkbyoT
70/9Wp6Ad2oFSYXwVSWVUUMTTP2u+GjPS8Kns2Qc3yNSQu957wg59S0P8BBSMz3wfKUM3oB9EKIT
RQZySS3JVI8B/iEcyHKCbEOSJMPL9I8Y1K6Iaxrg4PxBvRYyIFwR6vtAFTyL2Adaf+/x7469JPWa
yUrY6ud+9MlugHP/v7U+zz+ulFFpkmjgA8v3jP3/Q3kKY4/E/aYjsAQSJc4j9s7T4gjIOhpIur/r
eqn7mvfrHKKWnZg0y1T19jKk6IuTPohI2oz8JMIp8O8yvERmsCR34MiuODlMmREUeKbNwLw8QJdm
U+dxOiFyOTif+uTXFFVI3vz0MemiJtkCgRUKBbFTsI1eD7gpx81NGar0YrybnDkurFe8utghcANv
/ghFxzs2r8u1moNvEKzzCZo0Sxpnp+uEE/RdZ6AgBxAboBicQJkHP5ixwL9+bClTKy0ssoyAY7cy
eZ6C3IeitP6s3mVU0HbehbIsfdoy9udt7xiyY3fW21bIfrFSkAi3bj4bH4dHZYT7wcP7u5u1/vhH
Lke8CKXxYoNgvljq2JmCPpkeNC9zQ/ie5Q/lsmrvJy60HR3j+ztK3H/+NJ0UnGE8jHJhiuqTG3+N
0qFBDddm1b7KvGrxIn0DN8rdTywH5qWqoaCaX3BvlQe1ZEI810BU3oo8t/xhHdxvyXDf+lj0MpZq
2kh85oLD7NRbtC6TUYzQhhz3XFv4iTlKR+kE963Qu/QVmVq9Ikjo46UI3I7oupPdEkwm32ERlji4
+6BOViS6fiX5+DZCPykDlEND877g7yE7xsRLHlB5KHp3Fo9PSmIU2sSKG+hN924s1OxeuE/uuxGl
wuzrLHbvlvhD/K0FEQDmGUNSOJEPpZZYTuFRgi3S9gudDrmcGbZwTRayAMwxs6cf8SYbxIAK6n2u
o6clsWdiAvV1J0uWky+Fi4zP7b3oU5+aWRF8DG8TKqt1fuBEaysblddAWYcCrv/SfqdLGH1etUFF
KW8V30RTcf3cHnQnjobkdvfuyCmHGa9SU0jqrRdd+vAtopy5cxrHlPH4gXTrunwJQq5kAIWMlNUq
HDRXFNpWeXs63yjUJsnZwIdeLY750xWA+Qdc5BFMB1r1k5iaOIgfvXv3yeA21206vhY2bL7PnFak
zwZ7fSGo+3z7ftaxOj06XgYVElRCJE4hpc112tW833cKWLAe4226RAZKs12wqvVau9ot+eht0wzR
G9IiC3c0wbQ5ijIorjN+w/gA8NXMIpUWlP6cIbZXRRk4SVpNEFmhkVA0xaBHNMZcBTLd0wzSgMPU
jnpi+l73ZyVbqq5yVGekLefeFVRARzxBT+aNVtihtm5FcnP5W2/d9XkWzwocGAfMH3ozyS4azMBu
kRlVhKkneNvNlSGNdc2HiFqUPiB2rQVLPTSAdVh8e1xx8QTpOqmF19RtoRumvfSIRd3RkD0TALSe
InX8AdQNiM6XYGxBVWti2nhDWs9TXr0A1X9W8zacq22PYNxHCjSQUjXO1BcI0RElkRa4KOnvsg8v
01HEWOqMQcX2P7cyxanSmXQD8GOvFj7cRcOLZr/fVIGLUx/iHgkqFVOrSBrfslZlDX+n4vKLgcTo
iI/FpmAttRqekE9Wop1TcFjZe0c4qUTlbnqtrB2JOBlCr9IvVVKbVb2iICAjiWnWpOkhFjO6W7OL
WxJF/iPQgLuVc+xlKEasuLU3V0NwLl6rB58SjaWdxEwhLRfyLa4QCCG4HVjpU3zYOPeY0w8uT5OT
vz3BUWcXvFF6wibyNW38gXlDeuJZcraEbyT0f6SpXxbkSWWBcOaYVGors7fQBorsC2TcdNne3RF4
BEdu33VzObgDDRAOBgeasjX/wSB6viD+yHf0tKxBz+Lylt6YckXG5jtMLve4DiBBQRQx5sMgmGjQ
wAvOW4be+4Ck8QAkmwU378WGZRQ4SGIyL0apyV7JHdMl+IND3uhWWdTbBZyyw7j7SDzVRo6kdedZ
ieFPYRsdpU0yi02o8AQPQ4PUFE8ORDBSlXiLhrjufeAUwgsJYOYnSvOzcb82eRizOBRr/KU1QWR8
8JyPBJBjkHs+qOTUhoBFtWAtQ9OR4oBx86SlEUIYKGuEwKTw82o4jXmDFgKPPSKuG60dgX2Oh8i4
osGv2ksZAWFQ4SwmVoMoY6pt5BVDDZ1aHwqdjyOVYofZczQdVHiyFt8GaSr36aqFnNgZ8XFZfmHK
dfmcAmbhgQS/xCf7+yQ3+Y7S3xo1VbgXJHHsmaMwn6QsyIo37N+Bp6/QD8rffHtPeWYTE7Kgt+84
ZKmZcQnD3VwqTEztISO2J5Vul8dj5x2+7v8ojEk1nF/+xEx1ftdwjyTB3p7bLaucU/PwNFI2pbKa
lW4EWQS2GAZVBdKDV75XSsP64WQUE4oVtCmIO89rOWa5ZBVMmO2Vmp1zRPu2N86MawU/Rsvm2+eP
1xzkdRCIInz0Tfi9aqpeqVteHvRplpYlJGQ0Em0mVOg2fSkHOoUFzqoCyLhDDPAHtsYW6m10c60+
ddW37euxT/IDFyqwDsdGcSY3EkLbmBedwlF2ybZqT6Cc6AyXXQGfV/Ei45VkDzBTBuQHDPn+pOp+
VBabmN9JxMlEf/eMcNfCDCmoC2SCYvSAAjwAnlG6PvASIeTCCug+aqc0QP8C65aJ3HXa9flyDarZ
08WbllpjGu+vBHoENiC/xh5ZofnNVdDxIQR8nFE29dj9iLhCkd+B+/5w5hv/uTMtReiGkOT7wEUY
/sH54N0CbrJmIehot6tErsbVILNgz9FrWwSe/pSe1dWp/FaSqFya3KdHMz1FnZuDZmDXK+QpBN2y
aov2Ptu7x5eZLrbZflUms1HT482mD9mMCG0sw15BR2YhBYGFa6ulfvaDLMwcdfuuLtmQjUUCmbBJ
FPizCBuM5r4Vu/ArjrnxZ/lPWJgKWmD7uK6xj9SRcyt0tr+qkhM2Y1Y0jZQf0LddhzLlhyyw4OuV
/GD0PMmoSsSx+zwiQVNg58+h6s2A2zOZ3+qgXb/dTJkAM+56r/iaPlwm3mC3V/dqbyFt2JUTEakx
b36TdZyLPuP0hF4KMH0pfPA9VWQbY8d4RvKaZPgvOqTZHRE2LnO5yWuXUbMKfGmCokyQw8Txx3UN
Gf5Qi9GvS4yvXHxhS/ygiQql6lf0POKhZwFvnN7/AomXak2gZFVOgzf324VI/XZP60G84uSSAG7S
MbfXY/rcCyerna6o0tFjzY0oCJ4+xJ0DDSzlLN/oz87Glajbx0R92myYrUGvGdBgLzlMdLvhSyFb
16YQwgn4MxKx3R47ZxU1e3Rvdxbe1dEUVEIKPXvyL9ri9yOA1k+HHzrmJ2P70kUkQrIuhRpLDL4v
NAmK0dUBj+QV9nM4pr/tcR67kruW1gmPPAKMZTd1u1DQCg8cvsUpNzl18LCwb0KYPF87aO/o4T4s
y1DrZshWrDHR60eRmc/BgtcRKgugquPHYF14iz1B6Uhk2r4waqsqBPlWikFg+cDj+s+vBYkch4M3
OEB1bfDJhisuduSiXldtObLZOLzTqj59X69YZ+sOPqH4oyc8In5GlRyw2GPVVLr0Rm8r8VQCvaBM
iWoffa04XofbRoNM0PZ/8VOncMGILHIWHjRVzltFPRzTzRFsVQVgemk9phD4le0SGaDmoV+n1tOF
V9zvLeiRX9oDSm/5AX31VdqgZ/w6hFL9ma4N1xgsUq15jasZ3EOMEJLlsX/1q3gXaJZ09rwEgeVx
t2NJZwq7q4/7hyyzQ0uBf+NiJJUdO9YJggaCgPn2Un2xCeOCnHdmZFJNylr252VzOzwMoKzB/9hp
5K7K1144BSOUy28xyrL1o38N5TOiG/NctC7iwHyopTDpmGRZaruSwGijJMn5Qe1KXZtF02FaAT69
Y/Vl6Z/pVR5erjroYujLf3//7Hf0f+UUGsUP8Ee0GkCkqcCtggsa/BUi9OJTNTwIXZzbrtDkCtpb
oA7rCWp9jO8E3wD65peHZAobTdBlDvrvoj4AWXPOGQhO7tp2MKXxP+r/T2288Fdr6fg2nNEdkpNP
KWQBgYWt2OSLRvco4HHk58+sQtc3RXx5UxgSkMC4mdA8xnbZtNi6ZVEPlmfvEvwiA+BsYzz7IZGq
muRJnap7ayYPPcZSo6DEJd2Tk/8OZ0rauefFtcV+T/GiQzn7ljaPmo7V6hWZbdScJI5olbnOHdiT
Y4tmWbfHP82DPVyXsY7oH5Hmpn3urYlZ2iVuk84Dn+T/kjxFfPOm8TxwFJ7/2jp3z/mFG/7UDxaE
MkxRvKNPtWzKB9kYU7xTALhtR0gVhqSMupIEt0a4M0lG5CMbGiMrziAat6rxdzFqCwgR1SOi8CRq
ZdrzcuYlbv9jSclWNj7GoZ4VJjYuzLvb85albKWMnNjWwKmGH3nOF2RE9lfUHitYWOFmrwpt2jsf
JE7xCnhq85/Vmdybb9Mstbs6AKbxJYUe32vDIx9CDs9Uaovprd9F3J2z17VV9J0jfNi++/8SfWHW
ckDmKt07zf2fiR3hyGtjO7ZUuwvPKiKv6VwcKdqXSENBhXv2qLq4rzuiljQvZL6+bV+ue4H+IuZ8
bAEjcWmVQEcRNWtIE+g/wbOhIFt1omfsawk8YEvdI2xuf0odSDsX+Shoi9qtawdkcbd11MGRyROx
g1Oz7dGTST2kFZkN8LzZc/4NqV4rUclbswCA+QS+2y7dJQjnZuU0jr3EY7oiq0IDqmNQPOrozgtx
YPgc94bYiMCGODTBUebJum8fXi8oFfCWbXZAGtsYNS/4mUGoQpGL3wAbxCMr/1r0QPuUbfgBVb/q
lBCZiTTevxf6kR75duqFfbCDy9dbu4a1gVM2t1bFxIXTYwMM4vs+Y7oJ+WwGk91B5aX8mosr0EiF
1JGYxTb2XfqzYRs2ZnhaTHvIPjJ4BIsL4SWSqYOd0JB4/CNG8TQvhJfoih2rf5Ta5pfSvVZTU1b3
rV4JhMNt8VBrQ41GW4KHhNAChDMS32sCLfVP1JbdEvAkd1HYXTdt09StXpfVP8dBuyFvEGKLLsH6
ONBrQVnx7pxy9oURzqKqeGecAcSbt/Pe7I0QhNEYACgQZzJkhHREfZZT9MsfcxvKl6DgwOYyPWbF
MfOA0YgBkTUZGUhVxLDNPUaxU6043sXY3rvsLXS0qz30FpWC7xL/WrAPewJhDNRQsUjFIsOZKVNX
AXhBLSaWaPN1L+T8YlWH67+aI78PMfDxe/gBrUbb47HdlcJvx/Ysk2coI/S/hogrzxiMde9pxXhS
ZbPWuKOrDx3wMqmtijb37Y+piu46504RUfIq4WalEYrUxQqCIwIXlwOZPPMOmIgd0mV809iRyPHV
EDi2oFq6kdF5GiHOBPX9jQzU1AaHK5vylSsWMN9+8ADV6FN6Yu7Mu0qi379KxEv903ZctBq5ml0B
DEWZ+NEL6qEf6+mRhbr+yufgHV6k/rCO7wPwWnkLIFZpADpbRVkRybeoySlU9W6aCJwbSa/ksjt+
D8BYb18/q9cRNABa93wiQ6yGsx+RtZ4JvEaRV0OP7X+om6AmPEzKF++z42gh9nB6zCo0agevEexy
zFcKXOaRvEFoHGmKZ7XI1sSJ6lYRYv0nifboneLRORljJdo5ysBpGlYv/IZy5asiGiKcvRSgaD90
WenYYLHRyHvlbI6/w2m+RA3pXbKvnoQevCu6pEuv2WTrbhoQX2ZL6X7I7W92CE15u8VDiSS5s4A/
5vn70rVdDfqCLtHqGuQZ0bGK9sNXZbl2rDMrz2FOMhStE9bigLPJIo25I1ah1U7yUWjseKYoE7j/
OXabaF4L2Bab/4J1iDcygpCxjWGPXceNqKE7B1VTip7DZCwJpFMxpPKszBMWQ13YuB+F9GsdP58U
d9ArMiHSZV4WNsnbPe4B4FxDVCiqOFKhNMgEWqAKxDpyh8RELdWBz5Uu+Vyf/hFbWZVkIB9yoRyl
vRQ8EgXCEYghXBQFMd0zzq7F5dGEpNRH/V2YtwfvVPpg4HHuRupBmARAAHKxkNQ3WNm+YvlAW9hI
Lx1Oh1eBHrB4/x4RWPH9St9yULD1bwFaiO5BUp7e9PiQoNL92xqef7U8jY4r8KfnSq86b5YQ1pvx
03q5GqjlqHCG1vtLw4eu3r9tV56i5GS0lKp7qszDuol41v9MdEnYzB7RhSka0vtNlfEhn23Hq8WH
PkSRc4b+1mWIO6J8EFwo9wna6p3m/jjghViARsqLcbY7LCOF18JEG83Oiqxm6MAuDH3c8MvzBX+a
9fZXhybTrgbLPxImbMMVQLBXCLHUcTI7VvChPM0e5zAuVhtogK51jgYqpZ0ndFjDhMUvI2/AYAxx
h78WLrUvOB4tgVg06MhlW41tYNxO/ukEK8MkRBV/mpbo9Wku5QfqSPvqpQrcWwE6CwihQ5RGWsaC
6tSN2rbk9evM9A+T8g+EA7wLUvNw1ofwjjXF5RBsjRI6vDaHkM7UYAzbG8t1uDThGvPSNVJbv6sj
oei+1EeKHt50kWL/4t3PNEec3PweQlspwjGJiic3eM+oetIuQneyrwMe4KhOTJhogziSCvSjqG5p
OVKzJQO6jnV4TYbfipSu9Q2Veejuxr9vF3py4X/OtxRJucpj57TAhKpk7EpCdJv3U93QjykC8f6j
l1Bw5wwL8faYt4473bZicnR/3/u78GesYs9p0tJR1Dmo8lQ6tHucy/qG6rTIqL821iAtqp9BjBBD
2FvOzyJ7sv4NK+htZ53aVYRBPWvfMS2GTKSx+Zpr1zK/Sa6VKQGr5JYZJ0QiA/Ko7vnYZWjTY9pJ
crKQAg1UYuFJ9DIfrnOZTZf8hqJT5ogjK/JVmjoV+Y8u2GSOO7ZWcWhJx3up7JMCKZa9CHpZ8WeC
4uGt3hT45smfHF6HGlN6RGyRxv1Lo5AkHUodNDusWVacbrU88P0b6FLswFCwbzVHEwXFkP9Z1I3G
RZ/MRDbD5oP2/BHI1FKW1eJYVjW9Ow9gZDQLGS9b/A/9vjGG7ZEYrnMjdWwBfB/3GKBVy3Eql2uw
MBNUbSJC1IpMq6U3YD+KGpSt3vNWGSBXm8dcBhsBPOkSCXEl2x+WNZIju9wNd/SggtZ7wqYxsOGM
T3mdlRKnjjpKpLzXiSV4fE6mzyH6fe3MMGV8q7gDBHVM821J3nRLGcw3jz8za7UIKcKYWx9yUQT3
W2XsPGgqH6jKPNneYwAvHuklag3BU9RL3zFk75/NarNAEb9PPoXMoTMsLqUlFvlhyH+tMPFtcQ5t
iPaJXfKpFxnVAAGVjIjbZk+zf6lH5LUFVmMgURlvx/+tFneqZimrSe2FpogsRdRrYwT01lp6SCCs
UZ565ILh8d9/6F9mXay7bVnV11UewatwLTaGPS4lFiQHNca4vlYxejwSZU/X7zllVR1QymHUrUKe
lusCETEiLdgTXBwEx39kKDRVHKOHRAcV4RH3476G80gCuaUhPRyfG03WSOn/OSv+P4SScZbGYXMH
77FB+9WkwpTor3/Tc/OkejDrBe+BXBXt6Nf63IOeoa6rpAT6qn67M8eXQy0cPS96M53fN44OYv09
5rwxnBxWYzQIO+ny8tzB3agFr61IHI7FlbwXdW3VSVpq5TrbxKS9dN67nvLOC7xpX1FiI7AH1HoW
KWaa/mZzV3OGJVFg2F1kkYp/+wZ7BS4AgKbeR7XhLx9M9u8Pieq61uL8xHUJVYVE+/t+Vaq3n92J
33Vd0JedhLX4yTY76VTZvfV4/Gz4N4lcvvahXZnD6WoNxbDCTHTU7ujxDxWDSNm3wwQnVJEhN27p
MQt+23MDhPf69fFO9SOHw5TfuH0YUoF/gDtbrZXH1bG7eCGf7SRW2jcS6LJYg78WfFkUcmLMK9Ry
wkkQ2NWOTSkzXL1njJTWfaN3jBIvo1uKEkGF6uWt8kWYxUumyXdBekZye4QRMGTL/K+1moeR8/zU
r2Th4+3fBvge2UDKY3Nb3/9CBI0V2KIovuuklrObpiMxi7sSS/gMPEUmZXqirS3ZEFU6aR9Ak2EX
EPrbOn+HOowUUdszsxbwVmb+cqlbp0Ja7aK0DNg3KPThjX1eYk4JeU1o3PblzQxrwUMmdY40jiOW
9z8WVJyROL/4dhFjeUexdHOSXrcM3kYVlCNpoeGA9e1VxE6oFeZwjzeCLgG6UtAWDkKYEcDlSGW9
CJzTBunU0ihLlqz3XxpZgzU+YzJtZnRDssLLEp6LHAnZ7k0kLNDSbJGaByiwl+HyHK3mAqiDFq/e
134kJW1P4ZcnUGYxwDjFrebX4+cGxgUhfn+FlcNz9alwzlB02k8sD+cA7zW/O9lF8faFzMwdcFwY
awX/pOX/XvElII7B1tWRlfmlac0Q8oiqk/ZUokfqNMvAapvZiipWchlpuvFZpOSLlADR4dMFfvvN
Ve+t2uiG4jT4egWfdAMFXTvbLutzOss65n5U7Sp6TNVZ/8O+096JabnZgngUspnnahINknwEefqf
MmzkleHpdIuAgs231pO1M5TUVKHvwaNNztrhe2Vg/6ignouMgXrjA26wOPxAfaigyKnMNjt0CFUP
rpp9OoC6NprNiY8k0ptok795aXefeO3El+BEHev9647mUzbikV5s/2pmk/E2cstLHmgsSWhY/qhk
5/CnJNAot0fgz4CvDWIvc+wXt+MIGh2z2QiOjKxqFPQZPZg9HGxDY3ohVZXsFIYoTQdnVmWDdmCn
FLmuhWwOBAPjsTdiGx0zBA8oiWBQhRWyJYqOaymegkMc6RR2Ow3+pOHJLL2j4DarO/OkXSMl/H16
WyswtJyxcHg8ep77U3GsPbbGRSMAmRtALsUn4cuhv0jBX5SBoV45JXS5ehOw+WcWZJL62woeSpym
zltyXskUU8x4AOWIjZ7IA6+hh4OpoUtChdyEZBVz9sUf0k+II8bYd4r92HQ9yEwrt2OKE8xRshCn
wI9QpstVaYYzO+0JMkDlsu9YFXiQw7UU40VEWXUyErnuJBklqhmizpIjC17hSKFs9KsymjJZruz6
GLfEqe+mViBx+6sG+M+8p2dOFS1IKkz6uVsErDxGOjq+HJpTSYbCmgrmXcdrs5eNYV33Q2puPkNo
0LwuRWKIp7wWk9OnqsJVKxRTa7CFKO3vjrWd4j4FYZc4v3T4kKbRmDShSVG5SkL2AvVfIvjj2pEs
x5i+KIpyo2Ao0hhZmHR0tl4NNrtvwep5fUNDB7XnIhG5NRG0HQ2UBAqirsJyD5ZsBrJujI1idphJ
vyUianH2zj2vTikq7SuT50cmZ4pY1hhgzyg9f0qxkMTVeNISW7SyUEyQ7jEUOpclIrVIkCPByIlq
7R8v+nE2ANQDPMmtF/S8cKEFbP+mBr4B48vGeNtk0Q9lJzbPYsvVPfmh44uBqpjZFiMSCocwQslP
C8Y1enmX8kC1UAsAI1Nw+yx+4BwcmzRnTeK5oMyzyWqu0Vyeot7VELifbvffYDQmhklQBOUYY/DO
1wrkMnBC72yd3CtFTJinzPD1hySOtpDQ5oFquE8J9gOPArWcY6LzI1e59/dMulwqYlGx43ldBm+w
IsyGZvYcytS1uyHSlICB3OHB0pDQ7wC8WS4RHx3tuPkSSdmTd9RYCfJCkKf0sI4qJFC5AiisQIf3
R4P/EHk+NpMl/LyBUGCSM/1fCTYFj4EYeRiwJrTIFpOaW1+eNOhqfboIaISTSpjPFGb6fNm2wnxJ
JNHR5ZZ1T+clbcEkAmi5wu2qSGbW9bCKhxV7mc9DyBskZ2CMvtd2vrZ9dcoxdy4GAJIcv5VAmEza
GdrJT4GZJiYehDxWJQcUSImIyc0Cl8GV/FIKcF2dT1XYh1O0JmGt95IZFaHNm7b90EwqVLw15K2x
sGQk3RLhTSON7Xms/adpRNp3IuOl7kVE/zTbsYS/F5f9KSU2hkzy2PSCxbQw33vUPpDgenFDhMXS
zLG4kuTV5nMUdY5F/4zcHQzJfNjIrdkfNYAmp4RsTLM4aJgA7i8DmwKr4X/4MnXrhYW2Un3cfcfi
/r6Xek+SE4dTSUr73PfJ/f8kU4+fK+Vl2rizEMzykssU2NQDMaM/uSAh9nzLyvPpq96CAQOUsE6A
WaHVUFKgYuEkllD4qdk5Akljp7NRuRKmWdAHZzO6gtWRWhpztz0ic8bSc5aStRzjclnDgjG6uwlH
oaAWtSOlvLjFRPDxEUQJ7HlZHQPQeW2Xao2fVgzTkVcLdKDoyuTOa7g1tiWLZpCq/3RCUsLzK8u1
4smipBs65OpQCO2yH1Uub/7FuGh2A42Rt8XcQ3o83qd3IvocLcxv+3znP/8uHzHEnNJY4zLHXrzT
azm2qJLTVEzwzQjXCjxC7iYbMYdMRnY7XM/ox7N+FfDr0bMyOND/xTKtdHmYqR6NbaComv+uKlmp
H2/lcZ4AoKLms87v8J+DwwCcTtTdBZ5LbbPIjZ/Ck4ldEGifEhbSgRdEp4oW0FnwaSH/iixLN1eM
uhqDPYW/kfud0SMlilLFuC46e50bJv/Inqcarkoy/vnzAbo1iWnH67D0BoCPAniDWgBJQsV0+mbm
eaYjALOVsj8w1MyLn/mhTl0AMCVE1W6RK4TAlvjLPR0t8dIAJvYouC4U1ZSvGrtZK/9mOIMrw01s
stpnGP2/OUcLODGWLxo7FHiV5dFTLa2xW8mkkic7hqo0i7zZLj/iyx/6FIJafG0SFNgRdgS8HDWs
6VfGajlggC0ETdJctT0cWukrxvScxvHgewoRgO1YEpMynhEh616v3q22eLXRxGrP9+5slHCgDwhY
+Ws28/eyrMRSA6yubqQChfMEmm35B2BMCT0J5NRbbkQIUKLmOqKH5wIJXi1ohIP6un7t+b+IgxlK
aCYWIkhCcOcLXoUcebZxJ8LeXN+DmQcNpssMVtPC9eRtIw6H0l90z6i1hnjya/eQmn1gzty/ZwF5
+JhUD5UkXv/R5Q3ibcVNya4UEyBBGnXakAlsZOdMwoiTVpLWZmFgI8ZOPZWJJTlwJCudY0QnQ4yJ
yBsBQP+Lt7PmW56J2rxADI9axs1stCaan+IV9rUPmf8ec//uPso6fBtZ6Gzzy5JIHpKF0MAFxu4j
lPM300R1L8VzhzbWxy5TZTTSF/caAoT4xH0Wv/lMPcdWNysBcxaRtviBHGfNFvSelc08YauIq/eg
fTiBWl2kVQj7Fh2kemJU2Bjn1pmE1F6F2zaSQ7Um2I2GEVVvTbyAwE+q+63Hx+CJ/V1wukgBQK68
LnB8B2FTgfPiTlPliKZSW56o1iuA7pUGUTpYtiL6g7CWsRsBprNrl0wffIvec6bxCBh5kAaGhquF
2af1ZhofLiVVHy97aP8oiN76cM4x9AChLPGxcg5MZsjIK/41uMo12srD280byKokPE2znjPaHMFd
TvD0B4eCNE6/mPPeHe8OfVgbjWq9imB4LWFD4t6DRMt/QTY+3c/TaJGGFHuRvKcZZZkFsuU04MhS
JULQh85uFSpRp/SARaIhibdzrYvwtuSRlPxzQnHuq8BvT0o1QyYUgJPqKKNVZXM7GMPu7KBA/23U
4DVNkaNNiev9EtqttEOcaa2nrTOz2TZ7vhDZHaiB0ZSbjXH4Mmwo//34A+YmD5wcBUtUQreUcrkK
OcLBe2xT8rqByeM+9PGTufJNs4BHyIc7TwMzC1iUPzxu7vHRFXrFDBOnvwCExyPuYSotB1l9kWXe
VeOC1KDBGpbTh2Z38pbH6ezYfERcYYwk7KHlp5a7jqlaSxaFVd9KpJfiFqUM8L7S6FQ+L3JB+qEi
FQIUZaJbY01w3CqScvyj3UAB1mVg53/V4hXUuiOg7h5k4Yyw8Zp5Vd4qTlDFWwscO1DFAjIR5jJq
qk/UImUty6NjGoKCFk9oMjM2EQuelyLjqyytkShdI+FHLVTDVTACM15S8K/D7HSTARAzf9YOQAwp
YrbtRZXAo16KYssXtGCywe5PQU4eZIYJoOmpukuW77LTe4J/UsLiEeFYY9rt/TRmYAGSr9vY6KeM
B6qSPwk2d/eY5lEiQnHVBcGrDn+SNz4/SdRJH7yfEY3FlRaX+y8LeIkSkSXnNY4rRUsaE6Mn2hJo
w0Ip9NUBn+NIO9ITiA07eiOkfGDJkuNkDa4IZYv5WfQoFXPEcLsMifgdWQcAVFB01BT551N7dUVu
UuA7WxvbDAt26iYp9NjOX42mLWe8Xt7dI1PLci4q61w6araBOq3kAKD4ogS9RSPDuLrJl163oppW
3kSevJfJB0mtqMFSx7ijDZwrPCL3yBtSVEVF9mRcyvzUsdodNOn/1yM0y3yt0u5T1itpnacRQrqW
XfAYyJ+T+zSsn2weXeK7XjjxA9j2ckyZDlSoPh88yKXnXFTGGqULQnAPqrekbpAJYbPDfhbFl64M
R5scoBEOMK9jGDD8ymE4JVO5bynyV6hz97ygFYf6vw2zjx9o0fez67czaG/onVY2uNf6RT1MS7wl
bYIEsuHY7/9fq/e9ywLwATD0D87IQacoZpaVAwLq6MtrIuZnhiFJvRdXXPlzNcCH3qg5AnxPhNQF
1jIcG6ad/iThQ4d2Gp9bltmYoL0T6B12Lk3nlErA2w9CvZchWf4Q0OSpsZCrC6Ug3dYV7v1lHGhL
CwmazAJa2xZ1aTyqcLCP76OeiIXqGjW9LX0q7PoYMVr7OSePeYudNowq/mh5vVaVHCGG+xSaNSjF
HrwBMW/7Qt+Yo223icdTudABozf8pgcN8nkixi5TwcjIMo7kHWcJVctkDAHgMbC2GiIeMY1QdgKy
/nOmdv830XNz3YoV3Izo
`protect end_protected

