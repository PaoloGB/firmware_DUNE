

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
ekBAz8yb9axZHH68gkkSszs2QhGyjBigxY+h9lfHkc9ZGDMFNVVfdJP0K2+dUFwgsQlLuetsfkxn
F/qqneBDzxucfoqUBEieomoP9UwSRnK1DcD2zAe0QLL8Rz/TzCU1Rq+v/MxTZUEk54Fwl+TEV8HI
+WZE1hefqpJOgNi113uPD4kdpdVWpkIZ+Bce2V1ZzRFhqGe6AFJdh3J6dvw5uvZ5+e8TxAmIhX72
OIgoVnQepRrcuf5zwawzD/du4nPYUThVW8UT0Z/dmpiByD6oygWEtt9I0VnNEwpLl3y0yuwN7Ojp
nD3DRmGV7c7ZxIX5IzHn6OddoDcm73p6etxabz+BE+GKgzxAE8n+2ZDluMxF+tCYehmTWpJtL9hY
EkxryqKoW3J9+9+W0loNf4ncvGPnnn5Deim97OTwIU3TAeR/KlIsQ9XTMwmBULRwcOj4dh3sYeHO
5kab7QgWsJYYNTcMIkws2mGLXLHjZWZc35UBKiRBji2rPloetPyrR9NdJt6KtCvnycjs8Nd8k+fN
S/NnWd9ms+kjmhSEG1f3bAq8OtFUXMqUoWjGKZN+t+xbbDyaUDq0WMSnuTsMaLaQAApLkI5Ey6Bd
Es1AOLv/s+EX2pGj/1cThzhZF9vS7hMbbE53echtptR6vs4R0RHMm3KM+KrBY/N2JXF74Ym2MpXx
E4OvpNzpBQzJiNvdPLXPY4mwP9nlMyOxGiCrMKa+nUWKlsc2gLmgeIHJ03yv8H2X2ogM5GWZ0gYM
VazB8RPDPHYfTf/iHqhsB/yf89o6uc4w4atzTmIoBcQ9t1obE6F8AnZxIfOIqrkMjwkN6iflImFf
Q3e255BkKAB7g76y7aH7YR6qWYUnyoYJFtEw9S9q+nMyI4CxKFs+LTqRmMC22bVY2E5rWtckL1Vc
GRQ1VtewWuU+XbSgxLmwBeHHpo2i6Tzi/1bzLlklkpDBFdwz+XWbYVkNlQ13QBYgU0Hn0oBFNdW7
Zqjp7hIQTEO3/lCrr2xOb88VudBmLqJDzF1Y+KP5Qq0QQmlJfUFMl/iWRV2IYBqTYe1yIWEDosbs
mHVupwsM/ri3ClzwiT7A0EFzpjrbYqfrKIgflZ4NR9f/JURlz0JY1ZBV1W8HmBWo5neoeJKKLifI
IdEdEYHEYvSYGhj8HqQxmrm2kHDY11puIbJbh2OjWiGsXPeKa697ZtZsUDi77qW0hcnulk2sySLa
hEhFGo9g8keN7yTWz9YCJse9v9r+DH82xkdLzoCOY97+qKISj6FduWXT1p0rZxvOmW7VxEuQYWCW
+oqF24S73A5mZYR5OvjhINWwBSJ/hnusWdQpSR9p3ZQfHlfdYB5JfTNSggagD1e/kBdLoE6PJFeR
AatmljgAt3GCwoEkhQddZcayhRvIoHX2cLu/emH2Aldukm5WtUdogg/ThmDrCOy9gojSm3X9ebI9
usqC6DBo/rbou24ui+XJF5f4Qm2ICRPSS4hwWRPtWJ1kPbyB60fmDrwQij+ytUMTNp8uimTMGwVA
ApUjTzlBbtm7gNRm4e7GBe6CBMN/R+8iR4QYfJLl9QCFZ5WyV2qdti8Ag64MBi+NxOdBpExi6uO9
5aYcPW7ZKu9q9nmT4Le3wS37SK8hN5avrO5QP/YcdTG6rFSI/SQUH1hRFjxC2Zzooh6FPJq19j/P
5UbPKy7If7xeBTu3yepcDlymBrphQuw0xVqwRpj0tW0RScFKejrk7S8mojeJcxjDk7B8TPe8ExJo
SJ3BW4P8IHQb+yRMQCKS9dUUsV/mEbVKu3kbFqH06I95fYjqhawMHDW2viH1F/4CMj5/cyvKzbuW
07xJoaoAFJm6LYCxoJ6E0ODd/Pq3A/U2EKk1pyDwe7wR95TUERXR/8BRW+kyO0mMvP+Fk8oVssl8
48efBWrJJ5I591QD41zwaXODlI5GShrg84TSv92dgoKfrNEra/CGF996YFjw/krc0nFNDhPspztV
HXsScRwp/O22sUdY3m8sIbjmn0yy9++8fvMYv0lU8AQqr45cg4bxrhS3Z/4rbzKY8ZWL5oZ0+gEU
BH2jEX9oFBFt0pYQWyg+sHUgElqy8UyMBoiC1u6DkxCuhAa0ry4c+QdmX4OXqerTsKpYdyQzYWHW
milJajQvaZ/3ho62J2QPVlGr3wQsvtGymvc5wbRwaEEVyZuqIqptJy4TXGZbWzufi1JrATiiwR40
pzI7p7RaZerrTWImg2VQb0t+RmL5YqApPxbM1+eEkXpy4t+SlyRmxxZzExe1K8CIvxtnZLccBJek
6FSM/5HnDbSdHyG0vsdzkorDXVIvp5bBK9qsz7rrH3lwQ298xd6XR6hGKEtHSoUpPG5ls+CntrIk
LBFFFE5zaGBR3AX9rohilikHCP1JRJpfRWoI0E/V3Hq3FCYmGrTSta1OmeYQUHmJBb5v1ERWSNqK
f1KStXAfj+NNeUk8TsIf0ms5qIXSMcyGFcnBRXsODrjePvIXd3v0D9mK/ZPiHD2tjiZQSBZPcNfR
1nFFf8CTeI0zWwTDVT+AWaLTl/wR5n32snOdHlpdBXsL91HnjEqE9Z+T627uY3ISQT4yKEVwU+Fq
YlH7uzj/sLGGN6plQAfgdvuOQKhwVk8CyM0ydJcmFhMThLtKl0jxm/fp6DWGKT1xC0fHf3ojkZ28
VQDYf2LpP4Rz/vlG4hVaqn32BKRHSr2pd9uEZX+JUdMuRDaVOubZv1AeuCl4sEs9UzwjDHxQ3tyK
W413U56k406D7eORjVTyEQgHzS6oxWChRQnf+2S3nTy+GFnm1rIWJj6zsX8JREfGw1TNKqAN50ZX
m1A8TqGiUPNnM5qYGNSOpZkfaUEdPE6l14B306rObpQFChPhxWV3hSIVm9qxwy+eQPOspxVYKisD
4sFq/RSUy9HKwtXrsu2GXpaXunqO1RVBeOI7aqi1DrFaQhHIJYPDvGxC40gSc1dcrXnuLU4Md+zB
jlI2mgz6s715Lr9JTl2CslK9Ob2/SyrV1A/L622uVLEs5axdMKyoSi5MpqZUJpK+zqz3dmUv+oYG
msisDP7sljkGAyNrDqIHDuFdjNNQe2+5Yy0/lLBIJ9nEilzCSBXo/noC4Qmtd2nctu6RCQL1kj72
eAFAOb94S96yZ/nfwL5yLX+Ke1oJu6h6kclhCrkm113q/fM4VDTWbZeY98+C5CBZuuY0/U012+3Q
VWE6y0V1HLhkHdUfPDY6lOHsm1SVzE9nw+j7Zt7LxpwKv8C6/qKYAJ8Yo9wEDphoDxDR1uMuIJfy
UH28y+SEmsAR6BAp2hz7Rjphcvwc5SNks3I57EyqrRPjJXHkEPdr4k99/8lcCJoXRlXeQmGPbG3w
4dWV11cj/e7oO8bI8FRjXdITr/D57JaBzdnFaYqqfswKlhAKxLtTYhFxyH6BWk20HZ4BT0D55bYN
0EZSPgBBu03gSFVrU6Kwru22ba+sb11FjTlP9gB3eU8MlSkE1u/UXCjWeMXcnfxvwAynfDOZFxJn
IjXXBgOKv+kYaB0LJYZqWuUx+abQK/nKzRWWbrO0ak8GzuGcAE/ORRcj4LXCKjCjkH3UeUvpLRd1
euQY18PyRlx3X5JGefsGqPSxmL24NPhG+WY/aBjLFKiijLLMXLlo7cs+AOc4ENrXpLYJBmAn/KBB
0kcdJqLgeH8J0IvHs/z1XgpwQbwJrBqeMfk5jgfaQlCXATQzT7lzH6Le6A+wO2kRjSowKziCLeL6
C0GCJXfdyBouwwV6O3RMRKeaP8p+3YL/uuqsHTfjnFH7xuhcxyiVsOLUocfJlDO0qy2J4yp4TaHJ
2h8df99cEBdAwZ4wexMzWXbREw69dQrlHNzDZTHX9hV6op/AN7nqWsl4N3a5ZY5s/epyY3JzWYDT
6UixNJHnYQLFmUNiaGD/grV7zoooy5HYRq40p9H8dDU5E7Z302a1pW7eOy6WAkHag0tpvkfjcZT0
I2VIIQ7sElGshyp6aJg4OZVrtEobJ1oYI8vSlK//FojipqKMvuSiZVgOVV7MywEOccBldHEUYATP
nGyreEIhqZCRgzNJTvs+ULIlljqhzziFSF/UiqoN37to9oHWMLaDeS+QrH1EQF/6HWCxrBuU79Nu
GI6BQBkq3OM5kogB7t/z0qS56AhUkLhEg6oODV4f5vQsacaKDghozfht/VqH9dW+RmQ9jJM8qQz6
4+JoHuvF7tmQfyDUEYqY4i+Xr7bBsdD22+NAWXkmhHjqWSFskw6ldpoVLRBwmzayLWKTMuop9+B6
wVkFIVcs3U3oCOpFbasDTGbCIaniD+AV11hVuqbedjOP02Noa3zHGKFcI3kkZdXbT/waCZuMJTLf
KHPCljwR7fsdS2NAnK1hTUyRqL2JRWhfMwsiAD6J5aA4SlFz4aTuZoK8n8Q9yZdNjPaqFJ/mMLAB
34IJzNakehnN/vhwPYg+EtA87CyxislwGHenpgpl73gqu/VElG5uQsDsVi8A+fQ7fy7JwbKdLtcI
WRED4sYwNSn+2Gokt9YM8NoCcV0RbXECmHPa6yYkQAJssJmmRLCCY5q4Vq+5Ie3f5ruvERBQU0Hv
PJ8FVxdKE+ZC0l4LhmhpKaSjJw29x4bCNaJMdICNQnaEGRBrQk6XUz2JG17aKUp0VAIIkc7ehAdy
SFmx82/4AnkhpW3kt89cNKt6i7Qf5uPqOzAF3OZnozYHImOzRbXYNJstN+2X0JcK9L8yvUMC5K11
46hylha3ZkRWcYpcwYCGo7PWXpv4f9FevPUTZNkWkbBvkSQ2OFJJFZOEZryUC5WSF77EjlVt9a6M
zKUan5sYaYtQ/xnj7RzzFoC9lI+32r3XaWxHrpBqcBE55xyKSa1Lgw4RxjmmM3iGchyuJxlSHnSt
njiL0AIsC6wL5XtdiVhqS/qEUfeSjdROvozCAB36/6L1QevDm3kSQhvgiPS0d8aZxoprpna1Tg3T
KqKLCuSG/pikxy/bDRrMIReDormkO5MAZ3nYwhK/HDIxgT5YUY9adq/5M4ArNZsNyPYkHihVdSiC
aKirMjXYMGVqb2VsrBN9hAMxdWSB4+0eMwE3y2prop0EcixGRmu2vun4QE0MAIRipOKOh4CZgsZ6
ZScPURn0AYQuJHxZR7QGkpo6M/DnCBUINwWhEhjZI/2+UvFy/8niuZPsc04Gs3+rZ45/DahAyK4p
WqC5n7C/09yVdyOYbmwoy9C8BHxt2ayhrm5opRCr8HNvI3N59RQ/x8NMjf2UiTL8Dubj1UnlHzzf
NEW8DeowKLScxRfAotzocVwFebyj8EUOrN6aufgVHpGW7U3tB2gIWdNqbmr2VVRKYGa+DW0Lkje5
6uuYf0tvjDMjPd65WQiHiCRDhKEL8cJIIgCQbhKWgPZ/BjMBHkMv74RfiRHgCsHkHyLLb9zSLxlL
bLilg1qPdoItJJPM9fIb7ZOldROunZvaxRAh842jfWWOenELmc60r4gm2bkxnzHEqz8GxeGmqXS4
LJbEA9XbUrw8EYLHXFVN57ysRi3DKIVKKpPfrtzEQqGLRxjl5y9Ujn01jtqnZpX+2UVNlwfHQ1nL
MYZ93/K/UbPZ7oVXR6bgZm9NJMY6EY0lD7uN801a9BDDIiGoKHniNFQVjD7Rdc4YEplvf1yht2ji
68RWWPcSOXivqMM1cTAr/dbSTXtFpG20FJhbBTVtTM5r+qBOr0aE++4EtB3EYa9L5RPkox75aY2x
QXiypfpzVkUqPuoXzZAgeGMSHAAhR81sDGPUcNn9nkC0QxitAcgOhNkCzvE+IApxN6K6Q0x7EHl6
55YZ89URreevD/eZKD8BkY8MIaTMrl4K35u2gc4ljpSvaOmLCqkgneUXNe/FUU9hsLNohkyY70E9
23XX0G3uSRQAewQRfmOiTQccflwbQy/3/rCr0TBgY7hYelzCmgF9VEL/dtA6+vDMlT89z68KLyB5
Zv3/U7l2zAbamid5ZYGKxqYUrKTQu6vKkq8z1XAZ+8jiQhJvIKoic4dZzwZWauLLJxzDULjpXPmA
r/+6jMuyc75/HSmmBs6usDo7EJVarY3dRv+SNc/631nEIfiKxxLbwMp3XbByTpbNOLJbuEIRGtTr
mJxGbidYuGwu5nQwIiPCEAaR97gSjJXo7f2b5/V/xHDRYaopLjo3XVi3bQFjK0wQRBxm9aR0m8ap
vmDLr+133HDy4VfQEo7p7mCVrp9NoC3OGHjGO989Q8MQjIYo5wYi1GLQA2xTQhYV4cPsuVJAWGB3
YFEkkD3+BV1XFsvR83DgvITrVhWjhFqn04s00HLXblj14jUSIm5UPmRzjwUGm1LUUkyBuLHK+RBW
MfhejyBKI2DjXdISp8aVLMfca/Ok4nk2LXdLpPm7Mngkw+fArN+6PGAhEtEyqxxT2u6nu4p7GMbS
S5z6gxWK1v2dOjjh0u6SuUiQ+4Z1nWuF/m6ygjxbkXKFCQp9vYnBkeQoIMl41zq4zNrVSieyy+eD
IlUGGFkgrWyfqwP8t73kWPMarkQAJqoU8F+Mu4YjzMwHTlxVbyxnI1/v7TtMbvDM+R7Iz3BaUDCU
DkqNQmApUPaqO+ZluMdpmMAm0K9ncVPPO6yUyGOiZ9e91yt3EajxKUKdzDAB4DO1MmzaFPosPooq
0OgqFiWTClSG4X7VXjIGGr75gzwssGhYD9fIVWdwdtZUsiEKgz3426a5db+UUQYyjlbc7pE2HxT1
umCF5gFg6eWnp6n9gTV5XzyFTwSQRTvDUqkInZU4KknfvxUagoLtAqO2xicggTkc6j/9pId9Ze+3
5/SBtRQCvvKVEFrmGpw3psVpS2FM4M7TvsgKHP9HuGNnXkIUpA5HvdrD9GlkGRwQSvY+/N62+5mx
0FKDKXEGDMDCAIRXUHz5w8lIJHymKYkn7p+6dx6drzzRYiF4UZ/fj/QBheu8tVaQX4eKXHf8IYrq
0DJUmJmrAb4pv69Eu1IfEAVOucwZqlKcZ1FJiN5QbD1yY3iln7MYBApv2wZpjg3oe0vm/yoJe6we
Ynfd9x5s20yg1tpjK7sUO35sPVrMRD4z0RFErfRGyMQKSTTWTOpEXxm7Ee6azsBsH73T+vLOKzqd
4V+Y2mn57hAJm0Endeh+xWCWX3860SZ2DaEuBl6XSGil/K2kjBmVgkx4z+xLi1vz4NVjUU8DXu97
qLRSj0a2XcP4WAbSqiCbZazaYN4X7AcGG4YRUy8aGIGd+4CSPZZ6qCOXklWG2ImDbMbrIP4RDBnF
51APl+1QIRvdl/bTwxGLyeOIIkYSF9DRX9sRuK3qtGgC2UQXHVRJeIduZxvD4yA2BweYC7Y/8aCG
vsp4dSL0kL2yNE2teifBrw1MFt6zopudTxLjpKt27VDPdLQT26hOCVuvTLIpU8Y/Qdz3Ait8Xus8
ftzqz20WYcko2Tt2OuAnqsp3WbqfpWKJ95ru47OthEkH95RFhkruA1RFDOXptZXk3tRFHWojXH0X
GSENnPUgO9hFqfJEsm0lzj6niEsKkTtzo0xwdA9xEaHKOYenTxuAnozj9bb2aoQCqvAQIRpAGrvp
WwiRXCd0CMMtrZjuQHhXQHIgYGypuP2uzAFwRFiKq8GxM2zywfJR9sEoRdG4kidzLMJx3zh5a//p
X4QymOPYRcdWLpEZUozsHH2cMy3IPlC7aEhm7IyFVNk9cDb1UISo8xT0Drjy6G4Wn2tWTiPVQGMR
K8P2PHObU0CxdYRL8liZJXTlraYkU52WM1wSTOGbG5jm6mjHExBiLlMqEQca14GVpTwpofQTtJFn
5EY1qykvuYULROjekPS/rQM4fLz3st2QBeo960lK1EyeO1WlH0AJoFLgr0fNzx0ajA9gEKtdG48O
/1TCADf9siFWvtZ2FCQr5OOCACaxhJHob5EmR0Nv4nwexKdFQ2vc9NhRVcF4pS162bxl7b/tl7kC
+0Y6/T+14EBv6sXR8WDEQTDn0jrRO4SGYlLZ86YSd00qg5BMew1+XEy/Gserr0N+0BuCWNBkVwwC
2hC6rzNYQXREJzje4BRiQ75j9aHnS9IwAVxqQqxpHFITo7+0S229SrvutvhtTmHi0rdI6w98hSNO
dSDbHnZ2Mwc9UbpQN0x9lzNAWHLJKVolfLzcwb+Y4aKBg9J6umctOf9A3Ef5wvvCJ3YqcylWu28Q
K6xC7PquUBmOJ+Ajm7rLgDNANoq6kG5yTwaWmULzhCRCyGFW81/2nvlrEvU6UchWUe7XPScqz2fK
u0I5IJKKHuY2aS+PN2qJdt/3dWp+1otedzOIw60pu3CSNp+RcIQE/HCJtjrtDd7jT+1IPryXeCRq
whPaG/jB7vakgXciyByUyAFu6xeKVFhwRO1+0Fp+ySfmkX8ZfQUIJFkCUOPJkZbDQwNjED7QmRJa
WshSX3ayir8t58T7u4nOKTjUMScB6N2Mq2W+uPkVLNOBKFCL+TlqY1cg7Gvks9sfJvjxTT1Tl+4o
8cGYI4CE5vUk6c0WeX3+RM3dAsWj/9SVzftHCwm+MH0zJT53mm71aKQGZyZX0XW9kWnHcPzuC08E
7/ieHEq+X4LgrjpcrFMoJZSZLi10yvwW2QHDvZik4eJWG/VzmnEvRC15JZjhpLl+NO/XU/Sak5wW
pJrcqfNsYqdlUGpQjH2NXluOqRIXkQ8HD/7teeiGz3ob9fKhKfwOEhKcVFsZUwSw5SxWfp6PHegq
LOTrUP2YBlCQHZBiFerQP2BWBMnoKkweMxX2mQgR6f+s7PRsxyW9rBrN9TxwqdnADYj6F2LylY8u
Y7oTySosG9ItjNrBy2Z9bP4xNmwQDCEVnqjxynF5XvWHRkdeEP3l9aVzb/USEf7RenrcWFsAS6J0
n8DsoASALfUXrLJJEmvr41ZWFBWsjDc4rOFKB4y+EVy3O6e3/svqjQQVwsKcWNlzHsAxWPOU9Wzm
hf1b7him6EkxiNG0638ghgcyIkdNbGmCYiIfxk5IBMYpkVUxNfdqHpHwsoCF7X14dkiwzRUByJTZ
pHm2BLOMzKQpxBulePdIgsq6TJzCly2Zt2uUYjftI/BcsjKT3cgCg2DbvqrlO0ffIwvzkFXcRq/P
l+33SPvrnXDQG8TIDwZ9vaTVLHOtUdiFHu3Sb5fAaBiVexGI49OXlR5T32bT0BNm/iFaPjEnUAXU
xxE3lLZYSN++jcMPf6XE5Bg7+pZDw8zSenoM/hRR3HA7CgtemCwsDtvYa8nbZhIm1jZ9n6cocNoP
5d61RpMgnH02/5Y6L8YFBB1J39wTdwzo5iUwgMuAZgqkOOcFolhbwfmCiA5Fsv0HBC6/bxYetuTb
BE40lfdQmYEQHgGdBcQVCqG9uDQzzaYlHvYckHYsL397srjgqPCbkSgr45w09M2+/PLiGvkM1P23
dvR4oyk27qNul/WargHJiUwHm7KCWUYX4nhOOhFsEK+N67qkW33sL/0qcsMHoo4B2d7s3fcG7SvJ
PLSfUtFTxk01dsQQXKmc4armtn8hFgEcafCSkw5MHtFEn0zH8a/UCBMngL294Qu5USbXvdTK8sJy
k7QafWOENlIY8//fBVVLWt/xRUzxWT4GyiM+0ugQLU2M6r4cKPZKDy3VxM/7vwjqMO4Gn+ZS1KyL
Y/V+C32VvU1KUdL180L1OnBzdzOieU7AhxCdzx5k5nQVx5A0qgTCw55VCFZIbWBaPYYxPzm3AGGX
GOxX9n2asRdgoDRnNWbKXKd7l4kFQlQ99uRBuY/2grQ39vUW2bGmQvF6Jr0P8+GLv8HnXXHgd7Ha
VYVFFPJd3SP3qYDBC4updgwiGSNOfpMWI2Ca1nkDWAZ0VpwFsiCdocCLMceBA5oKF6uWTD2COQX6
SpmEBjzZrs4h8N0Y4a3eMec+llZuRy68A+9cBdmQswXnLxmNNEhYNFxIb10sSUgG6HtNcaY0qMbt
bZ79JuOgZsQnfrWF4Psdy5UYoa0AdNgee5abQJMTCkkP5lesQzTA+Si5FUzSas2/sOG57ncvYJVM
1O5jBUFz/OtI2VJne6Ljvr3XZqBmWdlM9BKRpw5F8ec6ToyRVqzDzL6fWOndN2bHZHdTS9QWRf3X
0C6glW03OoBgCZuGxu3ykitYlTCrgwYfQQ1lx6ht0ZkfwVnsRF7Cq29IifkUFOgQKdjhnhG/6Olj
cWiM6nvGuxxG+w2Bz/8w8rbvcbML7WjaJecZast9Sgg9f+xRZs3RwZet6W6NYNCTNKBz5VgfLmq8
PW9eAKJV+qhwJs1vrAOrYRT0cZFLFJJG02MRzYSZw0fGx7DLGgHIT7zZOTWCIGhOJcxnMtnN1xqz
s+7812dN5apbV4bnlS125Z+zM1eZFHHwpwA40/AymToWtl/FWN2HBrmZ9j0fQ6egi1uzb/Bnsbub
wsJ9fAnABo94LJVVYV4R1+pKZ3YxRxBG1X2l9BGsa/HCPOpvyQhDQmlC/lQrDstxMC28nOE1z/Kd
QNCwgnBqnT+5gC6ylRWI15e5/zmWiE4TyuqovomlpS1WuF8rNT0VcM6f3y1pWGgeQ79reirfLNng
wGYoLWqMucaq/WoNbh1f1O0FGqErDlUj9q8OSKMGHsmQHAlk2ZJh0OJ+FovdGlRGmIBv0d4lC8ht
HtMNy5ormt8DmSENj3sSY/h1uIWurLnctSoFS54RSP7zFhHoKP2v8YmR1Xweu7OtVfo+gu9p3519
Hl/sE/Iwq7JEHfHhTkv6nDs0SuPW9X60I55jX4RExtLN8S79fZ4lO+URt5BUDFSkrdQp/n93jFDg
TnInazcJ/fC/uSSeMND0IWrquo7Leuh8K2Def4N5Z1hC8MmBlrSMfvijW9j38+mJpdsGy171hJNQ
QyjWv7uxEpF7ruxxUzrEMFx8zwDQHSmlaRBibkE1cEqjxnIhMaZLHI8evqElkaebDLWSRw/gtTlv
JeOjDTp7QtmvtT/ZuKLT/FGp/9gFj55xzmq5juhgMyWJYaQJ9NUENAhb1Eg000wvePxUod0cR/FP
rY8/EdKrG1A+tgv4JLNqHSIDXPzNdCIy0ROnAYiZ/FqyIVP74QAiD88SEJnJNkVYskx8K5T9qFSh
HRbwzmud2HTS5urSMoeq/OWo+yy+PrqHMIMAHIIJTVzv76SXgSGKLDduFYWbasSeLhQsio5fZElb
uWsPm+yFzZrdkcZcL6dTHkC4UZfkCREW43RTtmqvXFi33FvQPOdOuHMGbyAYAN39m0DFUZMGXUim
Om8rmK4zgiCfQrddDbY598BX0y1BjvooGwaoJo3gJbMpv2UFsIGjzGHzYNh01PGYG9N8qWfPNZbH
c74vyV30dUSAo+vyOK+AeyVXL0p1j38QFHF1glhTtpLlLEVutIgVoAsvUO4xHqXdj7nOE4XP5oGS
TZ5m4H11f4Edrby1Yox6gUQYtV1v9EH2gi22y8MticlUpvxP9NkC+uURStFQNuhET4SN6cpAyc5L
+OBzcI+ZrmBA01TJoPArmwHdEU0uWn/DbqseLtvfeZjAbhAaPISlwgN4aK8hcXNO5k1kIMPklnQT
J62tp2tmr+/7zkLuIxS3rsN7T0hBpMPN4++DsdBZxunKiSIt1Kyt8fbFEO3vntF0DVrA7JYxK3Lm
bLxP+xmjRf2bVzLCjsCue0WEbyWHGaVDwHcXLy56JMq0BDSLOt84buOuQTG06X6AXyYaDw3dBscl
YYM12SJb40yV1GW09c3AbHJXTrtjICvm6JfvaAZkuL2jcexVZt43Afe+YDBjq3dZd2ZK9DEcR9gP
yuoFS2zOkTkLigt8pzylnSUmStVeGX7spyQiSz1k5qWvx4229arnPj9yIAYN52qHZdHxfffbhHVn
EPiprjtnkMf7IwfsSG2EY73Dv9CKMYnT/iFGQSEePdh6WbveF8aZBQIc0P3JUNyNcX82KaKpN6CD
0qB9hY447Cv+I5mSp1xnV70NdZQDb9eed67F+VpZs4mLYnH80gYwUsVvgfFU6KIsD4cKM7eo3eW/
NHJNI1KZ54KF6pnzluS3qBURbiWcQMkvU329P5E20DD/MUs08MjvaxXRgX5dDSL2AUrS+U5oFEHW
MdkxhSE5VPvywMwfh2IcA3j8ULO5gBcD4OffigZAyrknCQ0HQhYnXHQpaxSnlnnpyK9+HAvnV89+
h0d5QecZLmMX/QTDkuKenWy6XhhlfAg5nyYFqKyxGWSC9mD2bqLoeP+QJ9gjd5tneh0XUav7tqvs
4FNEJnAJeS2zqrolNp6K4+9KflySJ0lb8Ra6oefP6dofp/jfgwsKg6D4Db8RkBgGtThomBnOSo7K
WEaCrcNB7dHXxp+cyUNyqflzjNmJq6IBzJLwH5jUG7d4MLTyYbMRl/I57MwHLmfDcOz6AGcrywke
0Id7GlWO3KgM1cU1cjB6RmOruK10TAkMhzIfQbkiWpRRGkTnxumxfe7QtYyfEHDlK/XDOI/DTwfG
bC1qfvrqj423q9i070AIEz7vlMiCxhWJmJ+nakx7/k1hsji8tWstRsWepAclFxojNrzreewoHfZH
9nOssaQA140KXFgYx5NveO+b5MEbXkyZpzy/WaBDNisUqE39/91yPRudTtSpqVQzJdj78YnOdE1r
Ct9sVEQCTakV3HgDQXtIwfIrA108t4/T6YT1/3SENzU7AC6AbE1gvfG3q5Eha31RKqmqInDV1G/J
nx1GT+eDGhVKlKUfF6fFbewDZ3TqbCXR5fpCNJh8rm3eBoQXk5uloXJSwwGylIS1rEiI2Wr51chM
wkT5hZq2cKZtoCPu7KMlmKE81CzEgnFYWlbEKwwGP+OQ+huX5+wvUBShSp3W+PWNQq1LPkSJlKsx
tHlV4mci9KQMkKIJPd4BeTF+zRkSWtXnhht30QfS8yplnde5Qz/eCRtRH3AenSp9ou3LvORBmao7
EC4LfqR+8owksegEJpL6tCgZO821WRflaTYT0EgO9Yb6CNdJ8wAQDccnqyMUBepu1pPAZ6hQVuqt
2H2wEGs+4iwgTrejjzss9qYFLnRsisJYK2bGhN2HTXELbGjnc91zaR6caBCwKRkRDNBHXZMp7fFI
39wvZ/btukTd0xNsDH6QnoWKMTpKC1nYouMnpjerlx/gqIAxx9hEW2SXUVxjHuSSDeTj5cIL26TE
77OuCZuXSWG8D1MAsojIBB0ubsgwyRe8Ibw1wqlqpYYh+tyK16v5lOyt3/YkV/DeMb1E+H5xy/jG
2YJUDQ27Ya/CYXgxXdpk6Uwt5x3Zu51S7hnmO6P6LapfxaIuEdfnJLYo7fXwHn2JCToaAUowDF4y
pNMXQJpl5eNfvBSmaiul2lHUugv4nE7yo6ysPrr6YE4nzorG4cCT6X8W7Fkl0jh1qwXpZd4Kk22r
j/86nWMgOA7cYiFSmCfe+ZJb2Igyo6f6TJ3RBbiemwYDbFTD7glK1la7G9pXrrFF9ScOoKD+wg3V
/z4Eyp0WNm0b+0c5RKtj3ifQO4qZySJHfk9vFmekGxzlDV1zeCPX+eMJhOmGQFKyZVh1/xtv+GVG
PmvS9xryRkNWvX7/QnMs00nLxUaPZFTqFdYKRbwqWLIIbDkusr45GMKIe/ydgP1tr0ECazBqv9aV
4ATSRkte0jxudWmYEpybrvA+qt0MDJbBOKJuzyp8mSmdihtuG2Hlk18dfCFE8IsFHHhV2AWGkRT1
iz26Kf/HUVzvHwKG+dED54sqihT4o0cT23yDkTQ+i+28JIDSofFiCIzF1VmxsBmn7bamJqEnxSRM
kaIkEhoyQTjBUDS2C+Op/qpgcncTZNGqtN57GCHkPMhAsqndsuRjJFRyXWbArYVgUEUyTZE6UlI0
Vwh+vw2tAyjljswZFCQA8xVK6+eEx9W3GHgRwFeVveu0cnTkLWhWDqhHbuitfyoKmzRgwrtZvwPL
gxS4q09Do5XpsmJIk9Bqm+/wR/eJh/GI2Ors6qEnEFuchp5cYLKL4TK8lPxdURXkE87AStGFExxS
KKF+Xr79XhO6+1glg50xm0Zo8YfZNxqfPYzygy8t3FtbP9WUL3oBoiAEpx+x5B1MI7M720mg9SM1
rivOFMgJhBmh/w/2nyUB24gdBdwRc/dvfGzeQ1hZSn//8yxFZN21XgCweJZEYxtkOOxNFTzyNrbD
cBTxa1zmIopNaXweGA/uOjkg+ulv2d7qLGqQxKjURbl/sdG2nVb8k64W7kHv5MXx/OODJLKluda9
rlY96xUlJ8XW7jA2F0kFDMaMk8jfGw6/V9B4kUWBZU6K12cvKqqQOZqF3sBrbtsyfySTeKgdehet
2j7MgbYulK/W8TGBa0/rnn54lAawAv/JlgnmRFrUk8fyJokiT68sdAfmqWpBNzWRVKKCF3OnCEks
yLb8HbxrtvMaUndB8iHe/8AEciqI5NLZZ1Ep7dOho8w8f6E9jCA0YDGgJRO0yQ8YFQiyCUCSeoHl
k/qQuNoeONpSMTIQ/cDXftSg+BLxkzbU5vlu9rzYeFn0hjiKOsnILLoiAOwBBG+8XyMgvXQ/uP6L
kiXL+5PEszj2C8eUL/MHDnLCO1lAdJK0Uqs/vEC30xUkboYQ0tyLnGH7TmMSi/6XU+5t77YyGq3k
xd3ImMDf2eonOiKPGv5fP66AJQj2Yl/ZFP88OsiKpSFpEtkbGFj7pgffwyLPZpDg9zG74xdpvnd1
VlJEHapqOtND9onCwS8NwPt7DrlmOo2NRE115Tqsmq0IT+UpjHq8u8BC2B3c+/FLqABMEoxk8+yn
ttekEFIInfohRNIWHqWuwwFgBUDd9Ml5MWGqKqh6IQJ96my7V+vwg7z4zBi17/JA3lOOV699679p
B/7EAZlEyleMsRl+xwM3uc9Z9kQ/h6fTRxPm0HhyYuN68b3V50y10waeRNTUxeAcqIPy/d8dHIi8
frIuceuaESyMGEaHva180N4cMlyu8yEJkipGD+UeP0qto1vyp0XAn95utz7MBVVQ7xNNukSMEKrQ
/m4SiKId+PVnMU6qhS+brf1R4AhwX6EkO/hYw4syvZ5VGAIkO0c4LQFWBnr4g+10tkMpOavPnrZW
w2OFbDrYxI+oszZ/7kCynv/99MEatAbc04fR9+69gd2A4pczZdrxW/mU8Im4hpjl5FplqZ2oNohl
kZ+CfZRoWsysoNA6cJbj7m+dfJm63YAnKogA6KzTP9vUBigEuk/O36YLpUXiSjJuUMYOP2y7eEWD
DQvX/Ul0+SCoTiWUN7b+rCaU4WFcpsvivB7Oi/HfoiM9WW3py4lNf0Ifwm3zejrkiX6k5iTpkkl+
hwUYvxIvBqMzO+/CPl1ERagpQou6HRcl2t8OkLye7pux7hL6BL5MGKmCRTcixJ6RIB3W7LuEDT1L
/oKfQHDGsGL43BJPpnwn1H3BEiBVvVsj+GJQ/ftq+fmV9V8dKoLvSwKvQlZb68cz9WQHWQ8HxuBD
kCatzKPk+kodYMuNG2KMU55os5uyBuwY9Ac8KEkFPScKl68WIEpkaqaImYuJTxPmDas0+rzP7PCj
jGPUzc3SRGIddSWjM1gDPBeVKJL5ev2cwkh7n2vnPoqiNeO2vSLDhTf6Ja8+WTUGT90ggDWAZ2qF
UmV1bTNaOyuIEUIfjFS5AkySGKzHilaqRfXSgrFJeusGkfK8goGFzUKbnsTF+W0KvyvSjXDE/3my
t8xVpL4TaOYINreyTG1O5RX7EF1NWYxkLyKD22tHLWaSmHtrk7ODptNU5cUGCr78BwRgPixSop3P
T8HZL7/TMDYdDdQi9JxacyxcOf+C2iGcIjk8JQO8ZoVZ9cA6ZbNVsEO3LMhzRVwTavxwXUleG30c
pWQwz1F/ui8pb5XTsIK15wAmQiXCLeuhZM+1ZVIUSqcw5Fcxm2UoeC1sdofTBufZFm+JEECuJTcu
zkjm9UPSzh1pSe1WwK/9PIlsDKM6o24H4tisGliybUxt7PLLAegcnct15LHkiHNUWM+u+N3iIxMn
qM1NrAnwoMT5L1G6usmOain09KWctCNGaAFV1XwwMQInJdY/zwZrrCHXeWsBdRB1v3IID0xqOvDt
eCNi/iKjDjfCw4m0amXEMCwFyoSFy3mmg2md6UNwkhZpva/tJZSl9WMkxdoo9G5SvZ6STKe5/LMf
kGU9rPnQbP8ordYBGLgSqqVX4GweHRL3NqmaS7X84kirpDidb/pwp9eOY4Nsr78iUCQ9wmxOcFnN
LV6DgmhqUzmemnHIrOmzyS0Thg8Y9wV9q9g8uhqKjnDg3+v2kP7PywK1ZHRZf7bRmYxwHBW9P00f
ZEOC4ZqQ09J9d681etj55ygCXcYcvz510pdhVXG8Du4DEv0kN3TTMZUmspEo6rGeOujRvrXRZRUT
7J1F3txE7XTf6OU1uo8Ao4UOcPXgte2S/ky6dw5Ag5GBC5lOMilQ+xEYwNGgZZkLe1bK5oyHc3i3
W/5B9y6/+UJ/RuOx4mW3FhHFXKwC8KXBT1JSFeT4hThDw9HCRJjlMR13zcdPeKw/KIxZIq6oVLMu
wjlwmTK6uXRLlX68pZoM1T/QzVFW04j8OWFqVj1HhQSQVAnRd9Qxd6bOSAbw7i2dn8uAMdX81Bqm
aDBQrm+BMU9xBsM5gXf2xML4ifdTXozPefZro4udQcMc4FeFd2NS6cacZhxpngSUrvimr2buX0eG
L+Htxng9Ve5kquFJNXRh7axLAlQruFmoYqCKrFhvsbl6yqIqRfLmB5G0SfL+RFuXqr7MavvIM1Cn
69T+sYU81aXRJzjrn4aEHvCQQD+dF+oAAKbwmlbhEUNYNBjE6C1LX6Ljh2kpSFYAKMs/7ddUHovc
3TPS93KMKeXY8frJj6zhHTx2+z3xULFVVkHfbh00bCRKZua6h+H7ajWv9MM9Zz7y39QcN4eBOAlz
O6uAAKueyO2bVRiuVlKyGyAyaYlaXnkiO26K6vEUHDYI+Q8leA4X0A0VtEMw0RY0+v17dDPbQiPZ
Bnwp0H/tMCezr6/54SG2KEiIqQO+iedqfPO0KgcaoR4d1NNgcrd1+KEOsBUyrlrEeLtxw66zSH/K
2YZuTJaanINfCSFqwoj7BvUDxo17mQXgkJ5CiFEo9U9dvu0ytxkQFCQYExoui3sjKtNrIyWXWgTe
+0l1MgP19S/FQiNtmh2POghAeuHWXI3oyMhwSIFLCL029Y0pfZcVD9e6sUgGX5XTHsqY+W0en5wc
DqogrGNVIy1WzXMsQ94Q1kTNClwH/nkXvbhKGtdAaVEQpKw9vVx6kT2uUHxeW39KLBVb0GxlOMfA
VSRww25B59SJckDY9XVHpuGdsUKqcHBx2V6BFi6vdgpClXBm+UbFjWXAYVD7WIdv2Z4f/h+WBoWd
zB97JL+kSXhhb2UbqJDXq33tAY7BTHyYn+J/uqtmErWvNJ3b4WpRXY4A5cZ0oEe/STkB05tnrchN
5lhWZ8Hn8UFLUJFKCFnJxGi3Etq07wmNBGFP6wfLYrAQalUL92eIRA2NYM5EIk8dnUo1k5hnLEHQ
hPsdMPzAm7XBIQOQvjg+mgLoompn301BBDmpa8U1aGp8Uhqyh1lj0cCJmfj3VJc8ffQSmmrrheN+
BzFHcOMIsQpVUoAWdJ1NlHvR5Ygyj1MYtYnWmknbi6TrFScWKlEhc2YQFmckW/sb12h78Y2g6EfM
v6/xq6qxiITtCSDVnzp8MN9TaVuxpdZ1jUcEOsz70ZPyhngjUGbvfIZbQX1EAiRcsnZLDXlg3lbY
7BzrqdGi/WlvRl3ffKIiWK8us3pSaW1kwb3+7kcrKpA3bXf1vetBGGnPerBB7ByrK7gZwGS4N3mk
KIL2TYiqWQeJK2QtQlJ/HHxxpkgpC72Yc2thlS0e9Ms0OpvGFRcH8w08FGtGWL9GItOKaG2vFB24
d4COY6theCdsdMDUukU45NcZcv25jHrBN0v+mPNbWu1ByswBbwLX/eWHDov8ZhsbClCvYlVYNDdi
ZPTzk0Ui7TvBECIpMlRYl9BDZufCXTbIb+FCAGC8FWgef8BX5GYN6cLsjBWl6oxkRq9suZYWxBZ6
MjJvNqlec7Qqnp1/CiaUtAkiuCnviG5XfSCbTfVpwKQYVVG0+BCuCGoPUmolZT2U1CwpEL7m/bJQ
020JW+TbrNFn3/zNvPYxZd8jVuTujuFGVnVadmKlXTcjDB+Mnv6g2YAsKzgnnucEb2f5GVQPl2IC
CTqsOwqGCWmnV6FEYkHYDdEQ/uDrQfoLC+BXVFyjKljf0bqrrjwIObjTNsD7/Igir37jHuAxeOQY
+5a/2mUi8AIFo8cmB0u26E8fnzgbZIe472lpoYqYHMFsq9uPUMaN1PlUZ94VINBYoU/CnHz3CqiB
SayYPprZw1UkpSM0YGU2N70T91KitA87hU5yrWCH8hp8KMzmdPmTVh4dM+uN1tMKWjk/C7pbTx/q
n+4iaVe/VqdzGdrVNGivpNCeJSy7ZmLQcTgN+p03r2HQZcbe2z1cDo01jRu+5y1h3pbS9/NdAQny
NtzKBNH9r2Fh6W0I9rUw8uXITeQGXIvFgsxCR5X1FqlnqFYtHccr6FWOPRAfLBEQIg30PVBtXvNP
qzrTR9C6+9Ea5SaiQ22suFJ63kSic5tDqDPcsIcK+UOtfGYTK6qJ06fshu4KpmX0HI0d4j+sjSWq
kglro8WT08QtkzqGhNbLVx6rmI873MmbS50OcobBUfUR7tSGVEbJZgTxaOZe/REYf8obYdd7ipfI
wfo3j2NZin4VW+jRManVmpz2x+gPWVLcm0xPexOx3w/2uhvi1a/KOTFIe5KQnU2IgI9yGCtGVd/u
WxfFskDaAD6pcN9vt75YYCVvenQjv/zQvxnMSED4wJWACXIsTL2AMbAWfKJfVwg6BiQhr8kXJ7O6
cMA+Oh7GJJeV/xWT9U0eQ3jm/3VU35MYIjLrsXocGK/PbXB1StwmROkb3+uQAtEmOqH6CjYIXJ9b
VrmY1Q1v7FnOmntbHSdF2Mzf9Zgxo3EX4u4kPTB71wGmaB0M/+lOBvlWBan1/BHSBNsjfeEKpt7I
KH1hgSdhE5ybto3up242iWnCAyLIiGxUOkJy2BpGRimyBE9EwUBwejkRXId1wxlQOS5ln1SVsea+
VxKuHnU/5PJevvF8ccB2y3Ik3w8nDLu4qLpe45bNzdznLjULnDQE5A5l3jFY93AQPfPlbG9npvb3
SHA6OK6P/I2RuXOW1RXLE5OW6aaZ1Nah0Egh3WCePIYYx8Rr8/tJjnT2e+K9DwdI5WHRJLrmBG9B
QZhwOyhjh9tw2D7OH9D1nyjMTtPbd4UMGLLKUqJAZDqEAgUyElZv+AyKRm8lzBFSwflXabuNV7I6
W5Com+eqfr8njqK/Vg3duT21mG3Kn7JIMN+4DXEdVUBM/iBebBBpQqJJS9M0GAi+a/p6teOOdrRZ
OaiJDSuDUrT8y4hBqISISJHWUZ35n81nxS9tzcxn4PtaVxXX03nC+WR698RGPIOX3o3M26GGLy20
31co6OK2l5O1YDF0XW6Ls5/FYy9BxzXcDbP0ea4pmP2kTM0cbK+x6Zxsepx3NqwX0Yb1K2TmAFG7
to+Col43drqIs9eByKbOL1YQZ7s2Xc9Y7cocRp1dB2mtfF7mUrrky2uHCzuHYKplNZ2UhFY6bbJ5
/LZdK8lFI4vc/g1YqKKwasMtKI1sgrNDNQCVC1UYO6nW9gBKS1Nz5NLR6Kc1wL5WoA55qNmdIKki
F6KuZyiYKWr92CuMoGnzNmOspTDPYJXpfZIHOVRl6xosp2pkkeha41hG3OVT/CQek6JtlUg+MgC9
8izJgeXJFyTQvAA3NAGSWFK0mCS8kvTlbE5taJHglLHbUA/lbvlTaI+DYCI55lJgCvNYn6MI7H3y
vGy9/nTVT4yvUY/qJv8b/VEzRNH18PTJ5xeek8KOD0hqZN92JMeu1b45Sp6nh7DuG0q54Zp/xcNY
5KpBmQeFqgSd06CXxW4xOE44Oi1Xx+Fc+EslDUvM1uijvqX0oEQ65f54oJRnrky8nQ/yx1HXccrf
5KKRB5hCJXyjXQpI+0B+G6dl8Na8OtWuDzBWthZ5nB58k5H+LAZ28nf5XKGbf4laeJFaJI8nbfJG
+WOhiu3RRGXEl0nw6WSISLuxYitVOG1KuNgoUyKLt+4ouHXMz4dnjdGcv/sWjmCh4S8p7smTOFGw
kbJAiqV7Kw5FCYhG3gJBnX36p1vw4ePp9sWJiURo7AUjvUMw+RavVGDTqhWOXlvv9i5jgSQftQkk
7awejA2gjPvyz1mae3mJcDhy9VUH7XfHYtK615lUu31C00Ecu2lfpkdQuzjv+OK1qDTy+tnpFfMP
rbjI/ntudtKVO7Vrsx6hB3HJ7i+aEHI0oNLH12KQtuAJbN5pFy0mNj0p4mw05CgbxwDwjiAFv57a
dXho0GjjIjtW1YHYw7hO3ltIp7ovMCXdzuA4aMY2CvDrPTzRbrQfu+Jq6aFz1cP76J6WGTmx78aP
XRZNNHmbhDTa39zY0S+N382HP1+3b1qyr/aimx8aQHfYk8yxRZflKHsVv4UtTtIoMcR1cR4Am3V3
34wpSb+Z2ySjDfXxmbowbl+ZPavJ1m8WhuyR4yUV+HVNoPrLKvFw0lb+ijapL5UFuvH3qfglW/fb
gRlR6Q2uyJu24CpXH2dUa1B3jhhRJaUVq1uxTA2OAEyBEMdMxtK6/FtSevl46ynwDAzoUasBAWNg
3X72sUFoDOmS6LtgG/V3MbNpxYZ7jL8tWuslz/Tha2Gpwxo4aV1cY1slaGy+kjCCspW2Y+eXSIsr
GfEYJQxyxdXGPhNiU8wv9BtYaJEdhqsC2Mcucmfp9rJW08U2dtCXuNF0l4sTzzt5/bO/H4o+ic50
FGkVQwA+5hKn+FIA7C+HUg57JO4Yd0LPLF2dtLN4V3s7pYuSRKfESYG/GOnLvb3xyJlUpSLUVK1I
03ftKLuyaeqlPycsVjqMj1jIo39AV0YJ0zViHM4vDficnWoQ9q+opXcyEtmXsxL5xd3EXHDL06CT
vGI7DyFP1HPOHaOS42nrPm+5Zu3AEK7yBk6MnSejU0yWEA9tlh/3qwJTE56tnN22LLzb9FKhkm0g
j5+tEDn/SyfV0R/22AG8E4T8Fr+NB87lh4k1ccuzzg/ZDUxE6Prd9hq0rfd0hW0UgAgheZpio0p8
1feF10qkkv4WaHRjpvErKWn1iEUFyktUiWTZpJmx+p3fNbpNEv/xzMyb9AlOSqsk9euz3N7tQ05j
XH1aWtZ0SP5WMxGRnVYAGuZCzGBpzjTihmeA1T/ndRP9qcFqS7QwhYIKfxNNrqQvM3E5fDlvfBPX
uyIJDqP9l9qdlcrE1eB8bh6L6jf4g6GbjouHAV7DjPs0kH4mX/DRBwAh0OmNjkbvhljSManEzlGk
sZKXaU94pXURlgl/F1Bp8Ur2cYwaAB6aWVCW+iZAG3fK+m+SawcWLNlaknqwr/bin1S92dEt710N
3gPwmbgB0QkPhjoq9MjqnCJBeeAl2sfX2eqGqHq2lk//Rzazfc+SSjBJBOQAI0tabMRdsK5qgaIA
+sngBgPWHdELKF0ARjFDcNFK7C63wxlQfqktuV2ynxKmYY9Lnwy4dUpNgO5O2FYlWy1NlP1zj1hJ
Ob6Jjiax6QIgltffbSnDmsWWU3KI5PBgwEE3I3T2dUWVgijKbVZPEvYLcW0PhmFkVGXKr/ZnRcKs
wLDxAJl7UoCPVnvae/1p6UdHtiESXSZ+crXMTL7HKFhKToBt6y2J8acz+Usn3xackTINt8O20vjK
PkZy7gqeY3SeQZ5h1QBDwW6DhcWSyVkcOABQkebDNnDtLuAn9VDd6JQ8i0Gy/63fT26KYBVmEjig
fCIV0xGuAZO4dXYHFgjweD0s7S9lY5UwPCOAbnSkfVvpp9zbeP77CxTfpGtyD5TZ7Fy7th1/5aIT
DhjFwWT58xqoq0JmIsooRx48KLxTwW58dQPi+HWHvyE6MpO9cFaI/FdDbTNHbaZJgZ9D5AO9YREv
fWiXg0sR+0cO29WeQsPQ7hbipQRbaeXLiI12ohyodQFNOejiTD6yTne3Rz3v/ez2OoO2/gtgb6bW
Op4ftlGlprpF2NFlFKjZRkYVXVjnLPMpg0TS0kNGM8zlF0OoGssxgbg8TZl98vln4Xbgts8uK7Zn
sFKV2HOXMu4LJnWwObm26VhlUn4osWFYZ2i27fqWZh5N6Ic9/R7KobSE7hrDl0ssQgTGyKvfSSCr
HC1UhwzgHFTzqrSTq+FUkDVsYieW2LLhgD9y5LasJC4vOhw7qA6cbSZeR70qctfMjwabL6Ooyzv9
A9TqQ2Uq9KJiCQXSxKQlr4qJWSTb1DxV8jkTgRa+jwhnfhl5JIjdA4Cre9t3u+QpCTThwR0/APMQ
BWttbt3KoEG3uMn8m/tQsqnAM30FL1gnLHxsag3nDzMX9dvyiQ9/SS+X4yd32ylXFO7nQWFHNo1c
8DJUZKA7UUeJfASmC4uhp/CI/kCJaqkrI3cNEMlXIbFBsl7nSw8XI0Ke2z4aSO9tW2y4Ahdx5eox
rPriASz9rUMWQbyBn8If/P/z0bEo9afW6d59UtuduBmwaJt2cBO9xTK5QIer9hE7RrwfaOfp76DJ
orfHLK/4ANbmf2lkWdIByfTNmdec0Uk0h9N7ird/xy4koP+zuXOggOh9gP4pKtsaHEX7Py3s0pXC
ddPnFtDGbwbamFTorjn+VBQmvlwJFePnsjwJkv6IRkEcfTy8Y3S/GZesxFJuisWIz4ZpPhCwjgKi
T1MSfnfUS8ZG9UcbuYb+kmRGsnDgWqQytpwlVgCpnfo/4q2n6kiO/KVxo4/D87+eZGP6nGfmRctC
Rthe3YjneyVw6QhajSKKZE3fnatZ8+XK0bjxZk5wbXezxrml14Q8bvn9Y1IgYoxivw7ax1aabNjc
/Bz2kpsP1OVVWlWsTKOlb2bTRMP/PZGL5e5Ra/hQv4uEtdrvymm/hozSzj9VTc5wqedVwD7760hn
Pxr7qWdoZqWeFD5Y12mkqV+1Of/gq7Yn/SQr4G8A/fv7UWq0UeAmAsddNa5pguCBuyPFf4PdL19U
U/nsbDiO22tW9J/pHyReQ4cmDsIxgJgH6H2jcDx5Dx0+njLds2Q8B01tIy9XZ0NTX1kyUdLKckl6
fnHvfEurm6M96EgJc7HzrAl0WSBO+PsoS7Bn6q+BaGlPtuKePgbSIVjPzLh53HVNKbE/UKXRwpVm
pxZ7eC96tYkx+uV5u8ToJzysIZWa/C5y24VlRycUpXPx5h0QfOLt+tfuFLDxY0+osJ0eYnLsYL+D
pbXmHjUkqf5AVepPPXKx+CWFfT70sSRlIGuQIj3W8ITIpCVwf1uOdDm2ACJYdqaL0uCTG7Rr+uxs
DyGE3GZ7Bz81ccajbdLTFLGkS+cUzyuLN3UYTNgkGyGe6Dgj9MgJlpGkypXstaeDBH777b2eTm07
l0mjn/XtAAuwKrKub6k/QKWmTmXngijOBvhP/YGMuPaIw4fF3wPG7ZNd24TIXQMGqcUM3n3dy4tB
1TfaC/EScPzA2A8pYW2ahZdNyVhjSik6FJz/JqSv9gdsLreNgobn/FJZ+qoHQlkTz2wQSljNPCpC
hTdV4VzKhZ6C/3b0+ppca/qFPdBeWANBuli1CNdyRewdls4pFaHCnlATgxcak2HfLowjxhIdIEw4
+XE/paPDF9Vhl1OmLL0eVXp3sDSFJS1+MTIlh1fmFd9vnaIZ/XBtOs/zuIbKoe8EMu08Oiz2qn/Y
/o/rv0JF55xGfUckv7R80fd7R48beM+J4XA9h0zpoSEtj58XyP9G9gMRZVl0rJvA1yjmTskPBT9u
ABs4KbeWwWcuGcH/HBwBDui5mqR9iWOA6R1DWY5PVGtuOZGPc/w0Emyq42Oia5UI5QdSymY3t2a+
q/hj5+N3fsxdeNP7BAxr0kL23wQTMEE8soTrt+A+czVBaQNN11DVIlJQC2Tnh8ifuhmZGTSEkn63
h91g1sYAoj8Wae1hmI6fwDfQWlbsepke0xcgXmRx/g7mZ0gdGJafcJYxyCdVWvk+bisEDIBFIxgq
Wl81l8sTzV70O/B1jFsFS7wlfJ0jGBVfFvYxMpAszTEledcWEuiOByTN21WpyHwGUCwYEUidw08M
1D6tAWGjk1WhWNg3mQmmgMpGwWQ7wPBDGQJH4SC7t5EQt9FO0wItm+7BqlD7uxod1pOwZ5tHgUIT
1fSMbcW6Im7GImb+unLEw5g6toTwAmUPWfyrYefQOof3ICud7QyA1U2xO16CMp4eamPkwULMkAyR
QxO3/b76kE0MMSvhCH2V5HeLT/3Sv7TbRoSTXWDPlVEvlqvJTbS6UCnl0w07VvaUmDLRoyceuQvX
kq+9jIelk/F2Ma/c2TVt29dAEMUClWllmUh4ifc1KBqumyapSKdcTURnF2lK0M1hmeDZRoScMiMT
reZb72DMpdKA+eG4XOzzx/9nq4ErXvBJN6Apwhas52iiygURpTIgjBS+5ygJsriSX2k6yQlGagSL
z5Muh5Z0eI4LpXvvXmZfqqk4dK4rbRHbarosEhqD4f+KKRARiCsCAQoMPHJGw9P9Q5zqYuCKo2gn
0+bbnRleXMmjHS8v5AdSRLCpswP3x9v06fwXtcy4srRVkq0XVsx5ZzXdh5qey+GJLP+JoD4bt0Vv
I6FZDj70UMU1bBL48i0tmNzcyDyNhFVaVehm3gOqc0kQ5ue66qzYgj/CrokPDZ5iNHugI3cduvbr
cnFZzq+TNWTn2l9Uvh8P5UgdUU7yUaMc+0cV8V+JeximMl/yYTMiT+TAuNXssqVZ9tLDxYl16ZWu
II11NLOHHB3an1p4ozDWFyqzDajM0WRfbu9QsQN1g88Edaz6DVfWBuMLRamID74Xoc2/PE3dtRvD
1cJwefqgUScmn3igAbHHKilyUCfs5TRAyUFdjLHHDzRHGX76MpgUJY9cdbBKbEjGw7CAb0hL/Gfi
OYhQ81xcbqXhQ6anOOqfKqP/tBbqQ0UeyVzvCmPP76SowXWTdcijkWM2q1OR8BlEaIXlueQGf4Bf
xldwaNlMQPZTcjCNOcBj8YjZIKle/hQjNZJUMO78QDZv1o8EehLrWBNgxDSxDZh9DUHK+Wfs/JSm
Pc74G39cQZr9Iz2xgmXY+E3EAgSP6Cz4TPRtteEFWdLLNwNuyEroK9a4fvmKThoc3QKnk4BEjJpe
v4qZ15kf0LWSHZr4CdrDU8MzP/sbGdPYwub1QU8WwfniRG7e/kkkW7IwKb3ZzFJpqdPgcbmRdtW/
UxUfi0Sz9Fx66WWRBdjbjfMGCDbr21hmuxIWYrFFeptAedBo5dkNsOrpY6OYCFUOfckamEpGygO7
aqs2TiKVfhPW98vL29aUPo4k6YmgsiwnYHI7Gtv4YIoUHUc6ekfv8M3KDW3pSPu6PGC+LBVP4vFs
PCEQ4K1XMVCBS5vd77qV6VcjebgbCcMpfLZ22bJ18d1E+stpFMQCAF6PLcrxr8Jmv9Ca11AeGHmd
MFS8I9Dhr6LhQSwQ0lpiUC8JP/FdKj/bvFh1OiTPWG3wNl2S4UNzQMN8q4RbWBMUQeQDZ+/izZMr
a1SXAh7GNH+E1hvcHOiuknIxE8uhBPHtfzEItjQgK1nXJm9HwfDm3Kn/KufENB4ct5ubxT2z7fa6
kowMalWEnY5TpBypwOwCIgHKF0pscwcQYlFMvt7okVXOuxbiUsQQGdQODuSMUFJHYOW6lpeu6XXY
KUvI0wsjzqs5SrEnBzsEepYVD51lPsYom1k/fFyNA367KotLZPp0CQqVH1ClVScbERoWor9+vHa3
8yILN0EyFDBEldjCf1SG5hS6/JoHAZ1louChRhA9PhNisPbU+AGdbUu4g5M9WU4tTsaO2hpZ6rC1
IeummANSbYG6BVpvEVZ3/mRTWYwvjicQpkIK6GcSw+hiiSHuiyTKXjuj2U+BBFDWxAov4kcjfDRl
w0lB18adrOcheO0KloEQEG3KRKBiuCTGWE4/GHqI47HnK3YxKc/HwVX86Mhi1rdRTpHkOoL3Hq+B
HyrwLe+p5tGp6tCEp3sHTRkta3WzO5iDufPg3E+tP/mqcRFoVzNR0ko7Vb5w1PpvMfJz1/UX4kPD
298KSjXbNZOIXn7WBCY40ZOPHhZdMjBYR7k7Rp435gHmwuJvVMg7Eem7LPb4cyf5NHyE1dxMkpA3
BP3nHwPIHoVbR9DvdVE8xmGlRtU3A/6gHF8Rb6XpE4ORha63Or5GV7PShKxKln7/FYkjJupU/cs2
Ih/m7WZwEZwUQulyzlqn/Au3CM1eSXljaaXdc9MCCQo8qUu8JXLoEAwRxqpZdVaC7TECZO1iS6KF
6Ze/cwdyfMQaBjoA8BM/y0QpOE55osJ5dSTN2prhIEx+HiF2ZVFDD3mcqqqIH2wZBMVhNks/1fEn
bPlr5DuhX8mB8AaOtNGq2gMlG3ht4c1ssoba0TngJfd8bha5m06hOK5jiENs4GDL5/PWrZKx0+6c
4SUducAfAJcZUQSiw5LdZdzQ5PrOdTA71+rLqsftUaC0Ho1NeHuZdTwGrjNKVzLLDQ5OaEI7VwqL
LXr+0KTDx1Seom8eb6du4XbthcAwzlLgLtnHSondul3he+Cnbdi1r+911NV1kCfiGSVrXXbf+99t
OuV1SiIEdabR1IZudB5Fi73vxD2aH1K2l0kcrlQ2SikWH012hIeCCYfwxIm4t9Wxyj2aTfci+0iH
Kjlbq8TxY4mN1mAiE+nZd8iGEuKiD3X69hOcuGuhovXih8FtdL/cGLuO8K528yb4LJzNrnaU0cIF
0g5YfHIHBjG1ac7g0LkWqZFDTYAblbJD3LWXXdn6a9+POdtGonHjmP0P1QmR/GkyzVsyXiRLOlji
9Z9wewEF+vhiJLVZp2+XAXDiLD5Ug0bBd5ObSQtxx2PNdylPk8RWLb5++agpq3gIQKpD58Vit3p0
nTwosEU92oMAeDKEuZiMbh1wp7XppMEfjJS5NwR7dQ4ApPU+OTKR47fa0NSZE6pjpG7O3RhAL/dt
gt01zPBgaL8tuG0G7GH+AdwIQVmcWcXGDcNsThamLu+gnmJRjZPmodn3qP2XBOWdK90TKqrCfoCk
ZoThhoMYdmjw8P5B1q3Lru9n+usQEPpikEdIgNPFkFCm1vSlITCTlUIrc6UIM/DUlQBVRJPx6/9J
PQCyBMpDbrjMBS9eEYTN4K4qX+IoFALnf6Q9HyYheZwJBkCHo2/7gdhztYxW/HRc+cO45F6ijVZc
wqd65cwlj0WzN/WlAQOHnTOzKo2hkCZeG7ft3nOSktuhXywzL5aYsW2+75bi/IUqUVAlSVEg7toj
fvN7TWnVp+mvxbYa4uwARf+Pp9+oA2wuVw22RFzLF/5NsZ4S87lwvbKkPa5wmhJzN6LORAMF2Rp6
eIkl6T4C53fNTD1Jb/g7brvZxvS4dUjEKfBbEGDnsWZl0ujxwZ/iS7RynLIe7GcHr5BBKlMyDk/t
G0qUeQrZ2sYRox+92EqmbbmI6L5CVqwvZ1FDlYDTiCqFBbU3Up4wqUwEwuTMujkHg8k9CkrxCbur
3ckVpub+kP2IEmBDGsdSg4b0SwqB4bpdsOlK6ThkJkepZmSLxJ0bx57C7GwhhaesByRM+peWWUdc
I3s2Rqunpwj5PahCadIajSe6ToTHlh0zN74fmBSvdo8mEsCbfusaopQoakqSQBHFylHqSny0qf7w
MbpzJYrXilXFUvc6SDnMfSOwzEOXXc4HxXQLrAbHzz0+wwDxi12DoF0M86J3BsZ1PYEceDgfrmGy
l2EUkp5mb/M/Qa16atigstigm9oxccUP/VxfFDe0b+y9/CN1Xg5Uh1egl13w88BFTSjfOWAKXcNx
LmNx969XRlQTIfw8OxwZajevHy48XWv4ADPFztyMGaSxgdTTHRafTAFqObYu9GW6pwE1KIWXjgdG
Q7JiKa3CWZDtbmG+Lx5sBR/Naq6XCWfOQ9sUEs5f4mSW038HahTaHTGijV+ISocDECdZsNkJF/zK
lXLzuaWA+9b3XXIVyDbeLknBBerQaB71ceKyJ2TXOSgx4Be74wTyPtqRsOHWVUF57ZKOXa34dc6w
m+m2g04NT3OfRmrcLK+CCHqpvw0bJTcLnheI5Db5t8GaTHxd+PZf//i9/hET7NDznV7pwbH5Gt06
xIxYmUlK04MCUJ1IpRESBA3oZvrVlIO/LG9mH4uTG3PAH9dGS2UCWWZ/yv17Hrj39irzJeWhTto9
nWqJjChOIHe2V1XhUyW/ep6KiuRBl8K99u3h2YHN6pJWaflr50Y9OEgAqgSVexSZ4BEz6uHtnqDQ
MK0o1dxm+qpbRQQSJzTWgu09ivKKXKz0aWz/Tej7o4P3gfl9VlJAaiEZQRfJCw5V449sUPPgdIdo
SKBDG4GAnsX6OnvWMYpgoxB/Q7/hsvGV5CV05IEE78fVfdFiHJb12a+Jb+G51toHROC35JNCd2Wa
8yNPDgfpsMbUiVwUhe6x7dFaZ8MSaoZ4ZanKtag85cBfn7EywylBcCMyfQily0edT+Q27xnAsa39
xHPAOjqgaOygHDSwgUZMeRQdUbhpctbvcIafIKEn6z7H2lAcLqF06xe5GodEmZpQiOe6KqvK+xQ1
sGyH47NXc/e17U37rx/pZAZm9VkUMzNYlY+8i16+BHco4RJXEcRgd9bctyKPGZx9espBfud8ZvKj
e0HEV2jEYYiPYxxriiI3f1XJgG5uqPQ8+45Km23D83dQ6a+da+Ol1KR6tTWS8j+d0egYxgiP1L8D
UYlUf38QWNMlwGySGAjKtFX0Y3KxUVCY77ykd5S12bHUQevB0787TM2lzeaHRzCEig22jwghI0UF
mqLt5zM5hdq3aOVerJJQXbqC2POsUlDs0lhyZiAcNtUZlhvzeqeCxeDa4oVPqZTL47dMM1aErDc+
r3fpJaCD0tCCH1NDIYTgkcClrsg4/Ya7xDYcr2s3wiyKjgjXgKqvy7ySIn55+mEVqHbmzzHk07gI
JUL/tDK+KK43kEuVNNbfDJSFVCEFwizowaFg5D+osVlf5haWw3U2fytwciIlc0WE87m/waLu7VNh
GNGtRyvUEDNtTh27km1Q4dKJYyrJIlgyl/WQzGBPApIB60q4Sm8UlKKXVb0NQaP3Oi1VveZHSAOn
NLFeVQzbSmLPW1YE3sTm7BHsZZs8/S30MnKWncdR++0Y7ObMAn01Ix9elHsNsCk+8zJlPx6BY0we
jfkGSLyA2LnE/36K0K89gKmxkHEX91Pat2OBpVr1vx6d2Rgyoe+52MbDKS0ioJNvUZ1qz/cqIToT
x0DEfDMu64sOQzeKp2CREZDmrimCmsz58PyO0jkH+VB/72XelPtxfZSsOwHJzXJWuHYHSu7UULCW
FuhDuhbg96gPJ4HFcmSBukB8p3NTik16DkM8QcAn6PsAOgURP7VML7ruDdgEAFAu7sxaTOsmC3kr
ViK4JcmYttiftKBta/QnnohOay+8NbTDYpWpJ/O1hxs1XZBNQbnd4N43HV+ajY3ksZ0Q45/oa/tw
08seQJ/fnGodNViyoAzgv4MV9ZquLNE3wr02dvRu8W2eYeMtmvmlw3gPw1Pash4DszekzTg9CLrI
aiy2LHm0yKOWm+vTNfiGaZFuPq28Twj6ivVUG+sir1TRtPLeF+c6cWjI6Eh8MUbd6P2GrbqbzmSe
PmX+ZvCkbAZHc+2+MG2gmi90qmh6McMCcbUQFD02Fv0EHVNiVnK3GQyv2uneWQk97zQaYYZ6xawF
KUsWyANRnxmq6vrkHMbkBoBgwl20iHqyQ7bLcZScpQRxfDjXp0nw2Swu/d2PA4RQ/73oqcXbG/W1
gdiNKKmerXcgp9DbKqna0vH47BeqdtLWy2oDOc4f3Ww1eAOMT3grJnHW8ho5SLIhyUzdDAtVswd0
OMFVaXMa0bMORoWsBazBpEfuTUhXX9xmLN1lK3J3y9j3rWgeYioFLz+VPbqpLd8r/96sH8d7wwXh
Y0QE5xiWY/q80LY9/m0Jnos1qdVn+A/pnQhSxHl9A4/tnJMrC35m2UorsKuQ84E1DxyUZJ0zM1ah
sXU9COMUEiN8gy4aaRM178VxTMnrqDDoxWIyp6BvgqMlNMV9HWKQEruliGpcBNl/w59ordsTluh1
5dzboC4cyGW6pGUIXGRs2wrzl3Rlpp7/dkOM6Ht6XhbzK/a1JzVLETebvZ22cw7mEgsto4KmM2Is
ONbUfwP6lvP+tbr/U3/83bMvKw3/Iq6wCU5LzUgUqh1CoZ2LEimV1elO4U0OeWvP5Xz06hvyo+gf
KLeQMHAf2I/zeo8CG6vAnvG8wqcvJPXAUX3XxfYHYgPzFMhkH/pMti/++tbT1OZQNNd/cpA9/09A
yv3h2x355bExyyiweauedRB7+9Xw+YYFeEM3wX7LVS5WRFOxt/8kYT8ws1z1xN/ExcYirD0NEdSH
/PuLZv+QctT5US4+VfDJ/kUqp5wS+aCeTP2z8DuI+Jhd4RhrltYq0zsk24Q1H8/8myK6sETBw+tb
RXTUi3XpaELARKT0esZWe8k/e2l+TAdfbSdThJVZwarHHyAg0cbXK5PGZHsiOizGEwYrEVMf5L4o
GPwcA1jFwMtldx+UQsl3tqSpBs4qm50YwVMmewPkMulcb7ydEuw/+AggBe5K5XmNvkn9u5cN+fAQ
W1jJ8ErjESHCnM6LJR56fikpmBKCFE3GXxQW+Xxo1hTmUbQlKAEoHUHDKMmlUVZ9bd/B7M9MqHNi
KEouJEgVElebRcDHaP0/exKjTtmqjbl5vmZemTOfEnjiRjkiSFaYNoy5DJ8Qamqv3fSaFq2BEpgQ
p7kZ0NK7hhgJ94FBfgyoopW9eOu+7SkmqunsXvInOPaEW3IA4Qs8l7D+qPUGg6rueQN39gxIqeyo
/W7fcKS8DDlluXwhBpdHGVvLy9O4TYNx2lUlcgmDwtxPldAh4OEuZU8apcGrtJ2n5DkkXpJCzqsJ
GgfzdR0XIUVEo/2MhsdwBNuJQ2Gwqu9IT5ZoAR8pKhBxCwSIfZ5cktwHJyh7efh1Lj62djzAGWYm
1j0KOet5ukOETNFw4H8Hu+2xE/Ckt0wB11mI119I+5T21+kDffB657XzQSoN2utBo/7kbh866iTR
DRHRX80rdDih1kEvBUyl8VF7DG1lfHaviobmQJ7+erUdBMykDzrQSWNUvclr6kCqygERphlAH8B3
un9vF0WTscqxcude9xRt0pzb4DMQ2ftxqdSoPqKxst5TGAX/PJydNm2TamDnXlNl7aIMnGJZuHmD
UZK+GXZzNufnK6Qp05HHgMny25FIKrCwsfI7/gQOyGdYY878h59kbTOo7NK1Ei//Efc71BFIgp1B
+ixwEV1X+Lc677i6+CWVZKg0TLLfs90B4BdgKbuuS3SncPgWvI9gvDgJI8KdzpHLxqriuNmzJofB
8zLZoaAW5jCYeqzw+BUJ6KsBwIpEqyjf6aoEG98Mh/EnrTziBIZvksUslHJV+ZuQ5VLQe7mUZzK/
SouiegraKgrmBwe4nKItY0MCyhXnJeMc9O9pXrEPWJmmm90CxXHyNup3JQnqEQKDAk68/Ay3wx9s
C2cAq9xxP6D1FKx1JaWOOFX6rxD8v90YJk+XwY73ui5vGJiUF7x7ITStu7bwFnunwoElakzfv7tT
Kjc1EjFKyYeKKIfwulYcwsC2Z8NoYjOIgygRXFEq+JOGF0wNUxPI3AZAgs+Tfp3NYt2z4zgpisPe
Pprto3a3zGNs0OdO6QnVohbiLRhnfiTz8AYHLsv9y8I8V2TmP13S/Ci7lSLKoZY7jjAAU4WyD7aK
DsYXcGJRv3ZiaKtKvGPd01CQi78igKd7MjlrI6ficNI7SXDusSZ4PsmICBSbKdNRfwdxZ/xMMPyh
QWIIQxA2dc0QTHhdVEo/yXXjImpRxiR0aHEzvINAuWQvvo/moEXRlgGUdxjzA93qQjcBAuvngK0r
qjltZV/7aSKQb/qGwwsVnn0E6NphwaIzSp/oktaIbuOpMyDHZVyhlY1cu3zB19JmIfRoHRQPM3UR
7wEbrcp5Fv7Kd5gvjuqnEmQiaA33zemG0dbSzI9Kpn4gWrDv3oizKdPijUhsLiT2P9AUylnJs+Oo
vfxrITo9hY+k1AH6D3rc7e77qdV4x2lq0Qf8NeC7OFJ7+zstYJaDK4CK59MQvVcpl98VEwRKTExe
wgfZCBLGgmZqEkpbMPBsiY1ND6gftNhoDhnNARt+1CJKemSShltOg08F0DqGtt1ZHTLJ/X9TjrLh
qv1CdcYpAje7Y6+yPlPHjpRzq8isEU4R2gBxc8090MsiQcXcsmjJhYSJvMpJD9ZE/XQcyt9ss9Qp
nij8PcXlvEle1oivw3S98vOUvj5cLJawe5au8vxMTssO1Rl7SSR7an496BhGu9+p2Ux+TrBzED6h
+XTiQkbWIHUbwdYDwRWLxZBHoU0q9u1hgVte2yZ9VIWPt/bL1mnA4zIPQtuYouYoB+SU6IkWMJyz
PU+q0qx3VFiDaF/gPMAuAOt2jtZ0o9WqfePifuwfEHbJMhT9u+8bXomUxJRz6uGJ/hlcPxAjxs9F
BkNxiIWsekGkqamFX9nOVPrUzBnuPhFaAcHa1NgqFFLMktbDBFpl94le9NoFu0wekm5EdQmdIDLL
jurF/fs5tfKAC6MIR4ZN9Qv3U5WZFrm/z7+pFz8RsLB7+O+F1bAr7uxABp+QYGPnXk6nnfmkit+z
I6BOn93gsEkAMNMhXyFND+Av82zRKbml2/ZassENf3U7XFqwYUZ9Ch4E1p2/vnX3C7TESYSRPu9a
Y9wAssKglDDJ0iul+fSaBa891ZS/1fF42dHdQXMSsFadZxQrbBD2H5aHGeL/UHZG1RLhE5o4fRUE
Be+SfoRJEWUorN4An7eghLp7NoEzMdxtnVyd08zSaSTjt1zxPiNkP3jH1l3geuG0cPaU6yr+9IFz
Lwna7LQqK3hzeHWj1l1mP9Xl8FOK2lzuxZxNI5ydclLiBsXuZ+9xqYgmJPZ8IXIo6F5Y/mDwBPiN
Jy0YwUjcSm2Ga40cQWbXEEvObKc+hnI3jjZObBQO8l1WlQ7rO5DXRKFTB/GfSQLfLtm2uKMTHWzW
aj6VKDeUEf8M+T5PEb5nompD5liGws1mYXbMQ3mNCHWjg6bNFoxuN5vET5H7qtKDa+McnRBgewCm
B3N8nEEQtjHSXVtbAa5IM/6iontV9LD+gfcOrrYZfVcRmx3hdEilT47ce5QIagP4DPj1Akb+z3MR
z09l3tyAgW4hjIOb4aG5OrS87WHlA6kAwsR0X0ZlSO5le9FBD6kGCBRMNyshLFGYIrajiosXIloL
U6ZwwTyH5TFzy3SWnTUdTDtrFHT2k/l6oEnYAClr2k212dNw0cU/1SBby9B597vf35fyXku4i3uN
VJN0ZpwvqHOpyzUHzMiCcKOaNu9WeVZPjqpHt7HdcYgjc5Nd8Fz7cHUqe0TvXRFzy7VZmte5nbKt
BtHbYxOdbFprXMkh75/OxKc5m8xro0QpIpnLxH4BIP0wwUBDutOjLdWcKOiwPObEFepLODt/CceS
tl0VDSl3St09g98E/HmGiZAioCDEOANmP3Mdfp9PpUDbQCU2z1mMOWDKry6jkD2n+bdRAtLKtkjN
F5FfyOUe/kdxb6honLM+xAvH/kDH5vMCWdel+gawnLluJSZOz5Cbg7l3BmcdHChnJPkrQ1RL5gJt
o4mYCMTtJYr3Uw21KPxNAJOcU4o2kex39Kz9mRtiARX4MsrE3WBcVFjrkvHsxuGl1y+vbTeR5QI3
9Glu3XXIz7/9HpR+u6SbQIjdQGqSg4239UdN4s7wMA+C/q2DfiZJShPidctQF5K1k80aAOM8qt78
x4kFOJY4o3Afpqkf9dwjSU5+bWyz/89HXk4M2z3O0fT/k38LCZzVpG8F7ddILmZmCd+HMTJxBw+k
ggaIiKzHtH5PZpPtnkO/HdeC1zw4ix6TTaxMiV1Mcf+LRWTqKJ3QjDBfraM9Jc/YfwOCHwsepdE7
tCYS3zDod7K0EWx3BGvBGq5fWyM3dpIXdL6xb69sr5QdVccgeQUDPm/wLNnEjmu4PUX/4yyB/Omx
rMj6y9Zpi6xkVq3uMuzMfvif+V85KlxZo5O5B7+ud0DzbdRsFyFus2HmH3hJVEWz/4l1ubRSGMNh
77RUQtKDYERQjfn//ThuZ3QsGQQ/21GV75K4aeE++Hdq+R2HZlxVCSsMvUdkFYUulp87OMODXd28
iQtIR2IRmg2CBWue+kSH7sZ4sQwCGwCYSvwfByaLJBA5VqW3RDgv1FxdsiGMcBovJgaaUK01jxy/
iE/GwcBaoyJe3GVdlTFKQvMvTqlULG+Zt1evX9II6Of5z0qPjf0BKeBzHG1e75ThLSpwLs5hGqJL
XThrVEsuEd3SRob/CjMfZSfXiVp1nxz+EFo02i9Iea6jaga3bCFGb6xhRfckAfU0ksRaxn6pqw/c
XzjtxWXlGq0f8VIIS5U7mPrkp/XRVg9YXE6f9NxxITYRBfzhIosmaY+YJYxlKiNNE/I3hqpyVr3q
etpUfTBxDTUCRTtimSXk2FIeyUrhwpCsjkLVKRdI5F+AruLyO1vTpYUYhIGyl5lSvMMBMKZjDGKU
/j8LOkTQ23NDrTcF7S42PxzlvisQWQTAK/iiQ3wSsgNRUakkF8OlynLuW0sc/UBKoo5v/tGPshTZ
HVyQ5Img5QJVhmJya4dXa0pHfwh+GqK+RMX70n2OWfam8niFO78cWpZicN7G6lD5BJiii4YXxYGA
0U6cRoJrj4c7BUaH0OUZQIH67uCq1+HtEtUXcJt1ud8pg4Vqzclzw8hIranP1kpj+gg+M0HlZYMn
T/UmWlAUvseLJex+pZmYXl+eA617rmE2l9cBgGd3rQWAkJJIONorYugJ/x0yuU1cfXC/9N411nDG
4McbxJu7a8IY7vGdwCJkZH1cndTn7JlqKBSY9hffy+wiFA1JtPeWPuSEfxiSUJ5SnkmxtrfFWcAs
r0WFKwCu0em7OeGzeohQMwaIpCSf5kGkdTgb1ZKrX+a7nZ3ynz8rR9pIQwmh37cakDarfVOwIDtH
liyYnk0ecl6EIikQEFKD6hwYW3kSJll+JZvDVptTlVWYgdaKY/PLpz3mtc9VDzfpF6E1UUuYL+dJ
SIk8hMw/Nf9MObxrWrWeZJgU7Ou99aW3t5z80u6V/0nFsz7USgdJfY72IltfLTHj6lw6mI9TZl0F
yNZOYfXk3IJrejIgWMby+uEURTARDpp0Blha7Z0LNxY765nbh2yNIThJZa69rUN8RKHMihS9yZo6
Nx900hiaKI1tsyrz1mp5TFBn+stVuOIytunlgVhl+j3KKc+V/zPngRbgoEZYUqV93gvzBZPBV0Bm
DwpIBDoJJakhdFoFPLsdpoxY7rFETOReYr9mZjHo8SWthgqueqKqSz5OSxssSBVuu/iIecomQsgv
QMfeVr1Fi/vc8ifYFSWNKcoy0ahylJOYvT2Xf44ZnHh4HuROi4q6TGT81auJz+6W3aCttNlo+qtE
Mfg8okOSTLIR7GynbNyd5SPe/rkjAbGB4sQVyjAhuA7U8vPuFXwZi4h+yUngV23TPLdc23QGupxs
IuST1DUP/ibiL+O3EvwpKTFRC7QGxcgULM3sauHXyzWu/jhkHWiovdGSsILGRIc052jH0SfDpQIJ
ExGFuq+o4Xft1lgmbQHAbOw8UJ61CJN5Djv4huFVASu3R3TBUPkL7yKXMNvsPukDeWNf8A0u6Dhu
wWHoB99pjg21QmQF6QUtxVK3iFVNfRGMEQdEgMFSBL2U/9fBCGxntIgZ4JSqjLXrNAS4vawPDm4A
hWtAPcbW6fwDWXbIBBXlxSnk4jdoBL7WjN8B8VhJk4KSwHu/NKAGfLR2kka8qicPOfRGizILUPD9
JgbOtlPzdOWqIV98gMWPEeSbIrXpbc3ltkJf2FAr2I1jzgIzkLO/m6ZdvmhCB+BSZ+v3Kw1g5EHB
qi5yZPFvT9BF7GB550MMA5IyQQTF3/BYPPbC+YmK9ZfI1mY1eJT61ADgLIZ+7rqOV1oIIBZ/1Toi
0jj808PvsSzrKGGo4EWHmi+aNBnsLLCASxi2RcnLPhjxTZFgxlZky8I7TcQ1LAUSPt9lLUjyMMiM
Dq2QP3M+kR9xbvNrVQsXTGCbRWATFudT/h9S+wWWEzif1zJ087cnQGGEfJB6XPxEFhvrAAvSUTZw
glQQc2Hg+h9j53xt2uwvmVWytLqV+rmMRuaW5VZvCqRe9zBTjX0EKng5FEdNzzXSi2QRgC1kdcK2
3152NEfiy6LDPLh9Q3uKC4L4JjLJl3UrJBWcBZTiN/P3ql7r/Ka6kjLEFwiF5TwyIm6ZxTIaUZI9
2/6oxh8GVi1ANs16RgfcDgrgu/ujzxh11fdHqL+gDx9wBczNlcyyZAU4qvyEEnOvhwZPmlgp2mpw
hjf2Clx5Qxbyp9rgCz26IZPMvcfrWFK+pUP8iFLga1D4yA5MbmZUg3tnpHfLoGOM4Vc74jF+X4Az
PV5YJ4rL8Cd1pHbmx4a0F/q7ahrakwCsknHrSsWUJqxtQmmFQPeemp17vTZFTHsfClbi5rS9yTjP
QA/pbPXlaZ1235erlNlzNEZf50gvTyqbrWeqRwcLhp6ZYf+OWVPZFfwdCzcE42ukzDH6D+16p1Fs
UhfdjKk5yQsrr3U1LXkHsBUbKTfwcpviW7HP9WRZyaZyTWgwc//sI01XpFhh0+b1MmAifZaAA7D6
F/P/jvmiccgXaYxydDl4fge8V+ByOrPtX5KQyExN/3+otQT1TxO4oGaysKSlrMSzaXjMlDW6kUpv
dSic6LkT+VZOCZGXJ9LyGkW8I0RRin94x/cBnxORjr2+wHEd19JNb2+8iizK4J5Xhy3SyvAtaSLl
+xVdsqIsbF+nwYuPx/0TwbaQF8H9S3iPTA75nWTpe8l+oAh8o0CqoTjnTw2X/384bNmCtu3EMHf1
nFSopl0h9VcJ7YX82d/RYsdIp6x/TSE01u+JSwhmQO6mmgvAvCEUMFCJ7yXe/Wf0L8GQlQr9+/5s
ZS1FtyKb6PR1gpmmDKwUp7ZFJt2A0IW13ZqdCp06UlafWpGFqe7rfz2Ogox2nGymDeqfgJGsQggZ
ypIZUBYZjcbMjDQw1r4nYpN7rmXpGSW7urar5GwWtuc4NFirQ7PP6inSx8DSomuWBp+m3vRe1+ng
DdEkUNhSGXx3AffJBYkGtQiE2EXXXjank3pHhUhhtWqpst9dimlDolCrsrPNiMCjnduAQXvTtrri
dO185G614oFYHfMyaYVIZlr8g+ZDuD6gL1vTIiXbrii1W5DLeRXrOkEu1s4tB59EIrtqkkVyY25K
eLOjbydusxIo1EoosuU5l3EM5n/FjY7A5ZXW36Pr5SQYmfl1GwX9+MpE/Tdoo3N7Tq58nHp2W/Xx
HYr14wjpL7JKxHCTEwqRk+HFSIw1FwyYHSDCV3jPimUojFalNVeuRZpUdhpNxW9kUKI7X9pA3MbK
LHn+CsRCKWNkMAd4gVjylHISExvBl7qValqxyaEchLfy+ALFs+KI6eg2ptRluaR1x4qUr+2M2uOa
I+khOiCutC4MowTDsXWrZIoQiDm9ZQ+WnMpI8qPFnJB8A8vi07UA8W1M+EbBUTI7+f2ZjYOI+7x0
Z4BF82EByNJS+M1b4W5aHITlledpIkGnKPl8yECDD20qTXcUXWHubgDNHMmPK5FX3QCZCLd5Qftt
90uSQX4e2a3oQtx+CJduwMWv9wU9/ZTaYnS31EoI3QTyvc5YolFigvy0KE5t1BC8o7e7Q3dDgnuG
HbcNa7HYFepPUKdydUcNP3eKugEADEsDIWsoNlf/634/w0jI8B3h5o590JfUjDF1XfmRWolTMIs3
lRrgiiYLQI97ts8ie4WDhs0BWSQ2k1cKSc418AgKwvQUS31TOfUow2vhEl09q7hAQ/noRb1mpf8M
txq2tDeMbWUj2qEpqiA1jq5R6mlpd4B2A6aVIMxdHUNx0hN3Lk6zPK54P/BQPwyBR2SPomdB1cDl
9PiYGKJaE9CkUclY+sU5KBTCQKjzbXMyfiJih/xcKrNlA+ZvnPLSluVBoXQ4iBKZQXs2hnlNNevE
ezDtRXSICw9hK66N8BQkgciHif/P7LaqgwLY8JFNVWq42iIiIHDEUx/jGveX+B7IXPVr4ocvKwjS
wuKsqEbQkrVv1O6HqL6KOLKGVMzqx5Dm+fyL07N7okB1rc6lPCAozQ6lu1JpLXJzoqoZBhoZ3BR/
G4QvdFmAmmKT0n/2mFQsAJP6zirYK1n61yxDMTqYwVz2RAQTjUxZxkv3s9xWiudremR3bt8OR4Nj
2NncVNuXkXtP75Era9WHbdj+l/+mkJi0D3pqzpkzrKdU5Qn5O3eFEqJ7BXQWeCYlXzodE4VOWW/i
Hb9qlfHG61REtXTpIApS0Osv5M+1tjxdv7r5ke9DzBkK4mew6UqMESXkD4XYnLmLEdAYWKpnt7Cs
4OmIj8DUmrOHvx3w1w7jhhakbnhYLjVbUTUPL46c0yngKj07wiFTIcrJ5JDwnj7MBMu2eYDl+7vX
Q2NKD6P5TzUTguqwWjUGsc4bH8PlN72Hu6zyvwaZyuJndGsfaL1XndOSqauQtlJaUhPX1Kb86RkA
xVaiCz0vxvUqP6/ZT/undN7ZvT8kbP3iJRPTM/md3cc9c0R437jK8fLg9ZXgPiWuwtAgCl8nCr+/
zBFry7qPezYhQ5qAq/nLhkEhcP4SjyGspPJIum9axHu+eAMclU9RJX50RZq1M3QsAp2jtDc1QajN
wX2mTBGF6S0oV/hflU55Pd4VQJ/0oHTgNnqBUOrM/QyBPyRx81w0lvBO0o6YFm4IQHyw58ueh089
2svVYTKi/dMwEWdmfONLzKg3PbmZ7tOCw5hEahxa1MUdJzFyUYqLZaWY3PuzaqYOGQAil8iAe3Jk
Yjrl5od8g50RkgdgMfk0aMu6fCEkv16nGWiEoEkwTCKpJKH27QEk723qIpX8ftSBjO5qzc101fQ7
beBeyKS9SxIWtUGMfkDB3Q80ufLi/LGxbpYcrcxjT6bWncI4vpz3GxHDZcUcrmYj/M+T5V72nqqt
lhxphPM0LumD7Cd1gsrCj2jWykrTBFc8vRtH4okGFRVFYSHxB2dpPxvWe5U8rLS2hPWBet6Ii780
1bYKBUuog4J4VP1o85PSw/Fn7CFieWgIfChVGDxPtJs+segt20udZK4/NQuzZczsfFbl73ZSrKye
OYY9x6H9f91nXwfxFXprH5OTZ9NcjnbiTKkEhbxtUhz6JbkZ592ik9ye558Tthe+pu96yjVIua5r
JxpHjsVlge/hIoqwS2UOQvQ+PLKs2qbquoHvbUCoCv5k4IRgZ3CayMkwXC74yZ5rFB4Zyj/Vga10
ldX6IE0v20VRRwyZzDamhQidz8TL65PVTFrdFKhRuK4IDg78sLx7rle5sPqi9itjtP380vHloO8o
p4KPkymoEnyLHFLwy45zVNJpG33u2o+09aMAaCGRWPL1TrXZPWgKpTg9aarNaE1M6A9Jqbh5xVpW
BIHLKFYcEI3H2AfMeH+SmqV7YBCs0SQpMv6w8Ri7TcR2fMN4/BXkJk/30T361idYMcRvtLw5Q0LX
60AfSWGkJrPyHc2U0cEDua5duHt98cpbNnLy/FtmlYUCRkyMZq5Ek6gl2PCneLE42l5ZFD3/BxxE
JTjuxF4aqJpb90qK1hPrLc3xIdCPBVSnxytnKl2WHF+RwbaJmv+LCeSoZqhaX0tFFw/7MnOuohsf
IJP/OehSNtWdzb/UVFSJEY9R+GwHfRH3T7SZLvarNcxP2pyAfT5w0w+8BbbvzsX7UEcOgDt6s0iv
H+TbTaU3ZN1r6nUIy2FJktmUtPE2TzZ16/kXGX01tXIS6L0J3GNfuxb6iaX9BWdyd8c+pFOB/yjs
MUiT+XXp1AMS7w5s0rFuGENKv0oDHRA/ZNUSVlM8csAdG7qCm0AWgaazNSCRcPdoI+HcEYFyrvqp
CLRgF+NPgB6OsMQgNrNvO+dc71A5Ys3x4p+AZ1fFrBKNvkKMdbQMmqQ3SFQKQ9nkFD+7TDR3k703
u3jmweDRZMLy2aI9rS6tstcRXP4SCBaV24LXCCCjMcLQIrEp8rOvoBKz/NFEh8ZIgxpM0eAl1wPI
q+/M371jqQFreVwqfOD+mnP2ahMajXUBKXAIN5y3AE+issQL7NFczivXulIZPwO25H6+lDyVvBga
rd98x3DSKTFC7MGajr59zNTsb7mJaQNKEOHg6spdj/eAQDM5Vd/scwej6+ymoaOQvkX+NKYPZQZS
brtgpVYnwn7qVJD8osgojAfU4xiKg+4wV8nEBeigFs/GWysMIPC7Li/9duKiogyNSHhoac+U5zKP
sGnB/JhAvLRw6smvxsJg7hmYjp1CI5o5COXucxt30pvbiLARVru7PLk+9XDmsbjc8Y2O2uKXImu7
o8oIpw9U776hQOEB/QzHZqlIIFZWZMivxUb2wBnX49dUjcXbkN3urg1WIvTbxZMYsjlIRBMq+6Ck
scQu9Qnpd0Dhawia22+zPqhxIGkagFH8tQotmsdE6hNl2kVTmS+KcgPQHsol6CJQZgTId+Etp4Qe
XKq9rphr2nsLZOrCxMS5ECp2W/qBwhfF1MKL+bwnesNXsxpBKX1EAccftZRKGs392Hj1PmkCdhZW
sejEqdZEhd6cxsbvlWZNlPqwOsbx9Br5rADl7k32OkCpbio+YIMqAoTTTBF9d9VH7vR8FmnDjrOw
krlm16LC95XbpD4KoYwp+qU5h3XpKKqidqFwMQJiwMER9s8z8Cp/SU4Kdb1y0ioFB2IHo4reLwmJ
H/3rLU3TPIiJQzX1EzXxYN7eZbwq0ixocl5UtJ7+EdfKNdfjH8wppWjRzayjxDS0pNZeroLLEcR/
/b/H75rbIqVHEsfEK4W2iT0hrx2DYtK7pdJJMGVdpGZF15FhiGQXp26Cvf8DvYHmvvFxgFinHnzt
qgZ0c4Sv3PFLonAElvurowzPGCUXQU+D6LZG2kjq1HQdRBgO73+ia4OCZ2meRvwhOda4j1fiXFVS
BC2xLAmkfXdUivuiI2L2uNxgxyV0XCPSRftZHKKZBG4yxvBsEpEzOVstSCvfe8jYPocuZH3Zf2Bp
fGt7aBBGdnj/aG/7WDgSwve3+ve0w76CNWNrvt/WsacfgnwdwrKW91b28iBxM0OHEnff1PwehsE9
JIkBYW7Ab4wNSUlkZCeV84QuphU2+VXrIgztze/JVHRghjaBPasQ0/mW0HLNR3aCN2z9v/SlfzJv
DDgkphoTUMCmfQnvh+c7JZY/9EJTmxQ4Tks8By9rhVLcnfUfxNJh3UbZCXzrHF2QhvtajfeEVvj5
azBS/SnjBUz+oUm74POBi7SDCEfDYX85Edq1NXYPUE4fdgrD4CtYtCd9NGN5SiQ6KgdkGOokHgHO
Esw3gAJqc7TvMazvd07hEJY6XnR4lLPQ4E08LiqR7w6qT7VvQ9Pg0r3kBoENK3fHrDsPz5FEExCc
RqBnRMzlIjP4U+cGhLqCg1vVN+qfxrhwPYngxJhg3w0HBEpcPm8z9dUE5EExG++sq2/no1CqQXqI
6ZdjwP7DrU54CRtOZ3gj2j+8/aj+wMS9u76+wz8ZHd40ODRlVexweHXmqzBXoh2zoKnuPILWQz7/
Q9bQJ0v68znkEUTb/5ga8LrEs4rqDJC7PDiaJqi6OJR7mgv8LnoB8AA6jemEWQ8zVRLx4v1BOiw5
Swawb+zaglwqdP+4U1Npha81w0a80W6rECNmMZdKPCtG3bxN/p0tgvneiV8ZwCCqgdY0+D9MjobP
QwL8TQNV5fp7RX+Gk993+QU0pPbs0zfQNmaYGjztEPf93KsMce4xO9R4zjfVVdHm3VsoKBkpgcD8
nGaRZ1K++xcOR9uiBhWEGytZ0Z6QKyw5MruYTfdp2EN+kz/A/pwEdhyrgumPdlZDaKjcyd3Mna3u
0xLuF0ei2YvV5wvghAM54I6EWpcBXQ9tKtYEX6kEohP/mDFVOVLzd9LMoCLpfRbit4qcE6Hf5Vl2
5qpais1EEf9U+xg1r1s5yrDFiZgGaZdYIxFcWMt/z4wyDiK1Du5jB2NW2HDAVJtTLAib/7XCWlop
aPq7a4PaibqoQN4mh3n2cdYcL8yEVU7ERR9IVa6GPS+xwLkl3nqY1+5jb1SPd0w56H22HdUoWcDN
KgG+FqK1b4oNbvsqzzJPPyK50a10Q0Vl2GQDJjv28B7nRwqGGIxKvm/O78DWMWMr6UEOZVlxzns8
HSGQwSZ241yEUInMZaiOFXJQE0We6tlYNUW3x4P52Y26AJ7GS4FfaSwn9xu5gqRlJj/HGDyC6pYM
w9ICXfr7XmSvKi8FL3Ob8nBJ17Bwy/wMoXeql7M8/FxWxt+/ysS+w0nTH7WEzxSZ91o5wZ1etnOb
opWLWk4r0azYjnl0gcbMR2swDrmHlXlPVnjrGdzvcG7srrezZv38vkQRecX5OHpc0ytmpyipUXN0
vF+NT683eUQriQ5CD/H8cRnY0ReDMZXwyJi+GYWAn8X6xScK3Wx3Zh+aIr/yWBixY85Zra3ndYXw
mw+YjYOJoxJnAfLrUFCaxYkXu/itued/wDMyb3j6SLengjJJK+369s1sdYXdUGPMEYJ8DpZ8Yt1m
Vq0cGpKZayEhlUlfz7EzAtQam5J9xDtxa8o2RKAlHZCBWLSh5RhfjnUrqLM65tjjfoBQNWHi2BHe
lSwyZ1aIiodc3nM9XLXdEQZ+YddwHF+QT4nxshor0MDOs/B2SE7N5PfpBaIDcugUW9O09e6zNfc/
tMkzLEjMWKxXWceHrlBddHuliSBmQZCiDG0jf6vT3fTzItB9DTFxofgXxu11rQq4hvULNRnJQpcf
u7UYK3W6C9gzNuB/WhRu+sa7j8pCZPUtU0Jqby1Ph+xf/E3XCdjfFjpVyHAjQk/BC3+u8pOEApa2
B9L3e5rbYP+nMbrOhVTSC2lJ4B1Fgqy/4CPx4qw7Ss+DKBQ1OPaR7plTm5zuCderUJyEylcql/9z
XMboP1Chkj9BZZnuSQKkhSIpWaQCYRkS47KRJnD1g1qVSnd3YW6DbMuzFRWf9t0svZATeCii9AjP
GI82hM+ee4v1AETTwBLyeTY31Xw01B90awufyy4ISL++Iucwz+ECq15rA4QQY0vZYgUdSMh7kLSn
k6RJz7UmChZpYRThCRjLbDcaBbGUfEgeX3+uSZVUW5xmEYQUKMC6u2YOGWI98Z9ugfMyAJVeeNOn
n6vX2QW8y48laB6T0i1kYjVbpQxXTr8q+vzTDA07G1P/yhjCu9zNmiUgRzt2z4o9bm3z74RbJtQH
EvJ7lKDtbZtqM1jsncA4xLtxHcLMHT71jymhh1XU53jyNAkR8O0uMivCT0+YjFaIDu3e8ebBHGFh
/gF0+RaO8RxHpwjLoNw13XX+m5EbjzEicl9cEzOl4gWzWJHKeCbJIOP2aPbzJboaHEz3n6orLjaJ
+2nyveVW0RxeHjqBP/+NSc+OvDIboum0ldwV8j+sn10bW15FkLRT3AvzHKy1dC22wo5VWUN4PyyJ
AOK0+FIFU4nsIw7kX0ymj67N1/0lLCNHnvQCq2iKiqnZqMjTGk5q7pN3tx/oUX48E52IJNt/cEtR
4HTav2BNOL/435E/TkDChlcZ4zGzxsv5tDeE6Vii216lUXa5gJAZUggAm9Um//7rCLMvJuQx8JGC
+g+WWB+KjAvZUa2/mwkelRm8HWmfRi+FOpKHQBUSSm9jJwVuZXn6pLTebZ1kAChoTolfIvMC/zyD
WTu5g+Cc5a6li3mJOolD/KXr7lLDqnX+gqqn715dtCAd6gpMpuktrXki6n7PkZdc2nIn+QyKdlhD
1FDniUTAxvtmdnOHusdnvHy9fF6Nq7YeqnRGC+i3HlSIl8gKx7qH+ZryMcpJYNIt1/nh4LZ1dcB4
C7lSYYBAEzXX+umMRrDI+GrVgLfXFbL43iooRO5igrV50gR5tg3IlTlQ1LYUkJrwDpaWKAP/gs+z
UKfXuKQt7akiiz5GEbZgl8ekLYA4k6F5m7Kqp2EC1eejkvbF0Yng/28/RlDvs5WzV+KpoFO6GiFn
3TDgB80e3YuL3E+0OVrtIUXip60YNYdArZDxPkx3CWWBvROe4Q6M2cSeo9hXkkXSzV/EOe/HT+4k
V9n/uVZqbKbvM0xpUbANgnZ1g5nBuoSMFAcKbdO7tLP6uhDZC3pPnZE+PEC7QU2ZDV3+EZIPIr67
L5ZXnEdaAJrhADsQZ/0YdQBFq0N73oE5Mi9b2/tps3wxvtkAIxomgug80wCpP9FFi6XqY9Vi3UYu
IAwNg4gzShKyovKc+G7YND9d73Ga/rWa2sCAploEQqora0bIeKvP0ucpoNEP9hfrMZAguD37YDyD
eNpWfwAmzpQ+D/Alv0urfVcEkMpivf45VI7J2r/cHJtaISryKN57W8CKJgeppLYQ1Zyc0xIbPBlL
0JryLg+2QJSfXMCZh/9fXAP+uaPrlf6tTfNrb2F9WVP8yjyMw6JGJp4N5waHRanxV0qYa4qEtzRr
Tw4J10roMNgKhgl0kKIygyl/aIoJOj0+igjKMvyyUPebd/s5T6ImgyoQAAvc0LVYiyovQPQmbp0l
JwUXRBCw57xKtAKefOb9Te3IlM4bZuJjsBXgqDSxJ/x+crprO/obWrjTIEmxFfok86NoH/giWEgd
vnxk9Jo6tvX6AMk4/AS442k34dgQIxULg+uviNeTOvMTnuZBIm0LsbdNAliFyf0ZzL1O7uda6cvj
dHL0N9MyoeoYduT+HK5Blr+nvOyBRZHECrdsiciKqNxWEa4NtgX+d++oPegv84yzoqQA1EZRDlVc
V/E+4dwT56MZDnba1o9rjTpX1hKQoWOkdmNNcFbAkHRiFPR9fdQykQ0kym/ELgMDPWT5/dD/UuPf
Q6TtqH2YZ/oeGzeUt1bwGeV1ETDZX7CLT0PwlQYWlEASA6nBv0ZiMOimZZgfOIRcehJZzqvAdlF2
96k/x4dBj/RUsaNJdMS/qVApykoubo6x+BpSWd4b0qlWwq9xhO1AK49iSbQq7zf5piTuoU8/4Kgi
MU25ZjjpHmokCc5qA2obsFX6kN4/hEHNkwHRtwhs7QLhfqSIlmS2yX/tFyOXZFhNoHnkmsVm8WCq
FnFsE3Blc90Hxfoc2h/PJ8a41Fff5HpkuYdh4nYKFMPmCV/03QvTwSfyn3Ykd0ZHFDpnM+vh4V8Y
alLF7drrK5BsAl8gVhI/v2S/FH47PXFgyZGJVOC93MZ4pKIhSixJHYrgidLZNepR6R09Nc9ECrfH
YXtc008fZs2Ue7u8YWHchPnYsogmK8gr7MusNnz1UjF8PoEhj7AY+CE3pb5lHZPcClPhlU4SMeXF
eKKINcASnRA5tiyMQBMoIy5GXDO4ZUg8sczCx7Bt1NEuIjPQ8FvyiL0WDoEse5C6nS7MMFYQJQq5
jbzGTfeEau+G8SU3mqnfQTRb2CwJQXs9YkG7VezzKtiu/rBtg30fCVhP1GZljW7bsVjRiMMHAJ+8
HQSuHyI8AEJtRtawo5ad7kTKx74A2pKbnm/dbZ2mSw0U5WFEMNL865Dsid4Ox52mlvz4o8RObQCP
DyTwabocx1/XI9GWzIay6GqFTVr0LG4Yr9dyTi8eQ/iLZ7j0v2pydYOfZZ5Nn5ksHFZZYReykddD
e8PsjWTDolT7+EXIh369MxVhsNfiIH5gpD5lol1BLh4XEtAkbfwfkTZCd7D+vCmKCEa8mM3cAzjN
6E4JnRG9dwC6uTTm1vwRp0sRKsYRezBEbVSkfswPGhfyqxO2Ea8AlWt8LfR1xdT7p4iNjxQRdv+b
5dFTZFdYUjZpjyX8/NCxBS9CCkQ4BCycR67wgb1JzrrlQqvlGlBANtgq8ncDAWXhqscfe6kLHb5V
MyZcKmpK90gv0BGto2t2XYolE6A7Dt9KSICC/AcDoETRuCpxO+R3ps6CXchgrnuvf2xP73IJRxow
mRZqZOdxs4a4W/tVx9qE90xrtrTWYzTW83XJBg5CYDE8zPafFUrkMbXHPT4SytWskedivQxeEinP
DoJU2H0BWtBLXgesDHMDMFSbjtW3Kzo6Vs8S0oygktGTjZhAf9o9y3AN47B9irudahO/kscNLo8K
dDEOpbFPjML7Jv/LmCFB/r36qUeccsg8WUeNb+nErGor1TDT+1rmeXnEi4xBBFGwrLFrjviuM/eI
uBpgXvo6uAUjX3VWsY/zPJg+tQ8IFCzyr+MZxm0/PaLPZ4EFEUUNylzwFz4RwIgBmtZs7MLy1c21
o8477Hey+jgI6bpbF+/hKHmm7N0h+s3YChSIRUQqf/MkvPOJ6CYP7DcKkxv9h9nOorBwcvCyZh3X
+ts9OegL3yVYX79q9ZZLauMA2SvmFthy45aRfUVhqVcc/6Srem+JP+ldzE/gi7W//SVbs8datpiF
51WBelOIPLegYC6v6wlk2JR2dDAW88i/omFcIhjnpw9eucemu0IPh16UzZigWffzbzbsqse8pu8w
a4v8Z6ks1WL+ZB+usFokwGbbDAVHBN2ZR6lOGHepzOJFDn6K+WU5O/9aTCxuCeSwu29jnGDkwD4m
TT6Z/9WbeRpVbcOZG23yXocvVTeBzHuhLc+xful3b4ZI0vs5wna5fgvL5uRCKNPvTzYdhWhTNTS6
2jmotMgrp+UYJys9G6VMYtVqLG3eD3hZ2oBg4zwzuz27lUkjPDfW7EVZneuGwkJzPjJyLeQO5cjd
0EFR2LYp8au8EQhEJy/KoFqx3o8UqZrpdeEaK6YFqKTwoHkqWcVxyIaeBUzoDZfrDY+sx+V6p45H
7Pa0A7RI52ksyLuMCjGjTtgg8SQXIsp8dejCAXSxe1BCfwqL9gcwYSTvwVAVRqSCoRt9VAMzQiGE
S7p/jSPj9Tl1DEy+NeiGnGzWJwwlJevrjU6lMEX8padlRMfN29RkZhsceJkPp6KXBRtHy+tZKOaT
910fwJPvvpfRQ3ysU8fLFQUoumSmEAxl/8nUHBNHmRCam1bJfCdcHjelapXWvpFgmbvTAXQ9aMjI
KoHIloCRIHc1uebVqFqzhJD1LbcP18Rm8R2lu8mXJFYzgpUFgt0ovtS6NRUwzsHcKqT4KPpspgmG
rD/AiXI+S5X4k2p3e+fxSGqy/2mb4PbelZ6Jv63ufD2xK7MbzgkhiIpoBNC0p+Fxh9Jx1s1Q4ZN9
S7wKBKYJdIZ8d5A5EC1cASIvK3wAec1EgwS6ukFxiSkcRgpffk1jdF82UgCFYD2RnxFe+arysC7k
hg8pl+wYqsHB3hmijHYGvz0IDa3RVC0vhI0N32Ny8haXW7Dp4SfkzA8/25TT39KBmran4cQ/QUhT
fQXSoEqBliKKxk5Lf3JQhs6zVrCvtgcDmUPvL9OfX47MlMbwRD4NtHxY2o/SBvEmuYaBnQFjuHbC
cMPShmdbFNfZ/sOMUZv+mggi3YycURW4hVxsyMoB7KiUD3EY92w9GX6c8EjZSEvCdY6YQVbbsf1K
buohuxCccBYiVF1VsjNSqbxAUVC9/uHOwb48M/rfuWf5Qr1ZnaWZOXbAbl+xisRhn1SGNOmHfcdx
xBVDd6Id6611NARLDjTmsqwMgla9YxnfrjvW6prgPRjP5lalPbwMFdsNFjJwitH5dmjvw8/XSBeO
rDcQPJDxqv2/zxB7lpRi5K/ZhXVCirJI+lU/YXiaZqchLxn69kE5Tn08Pf7HInnhExqfEWil47Ho
sTJHDtFiYP6GItn7MTMNHQtzHAKHseN35UMyi3RfTTopLmtWTPdK0UrS2PhoHDwoBq+AKo0OXM20
Ki/TrHPkhLJj86/sa+jmz854htwugluwX/7PQOgfVHbnenL8JmrF3Xjb17LExsmU3cFk6iIMck69
bDzb0JP2Zvo0CLU7GrIOk2ztqbW1IWe/+llc95kLi2y0BlOWOMdlAnxUBxWriZy5sj/9m8QZz8SJ
Tiwiq1J9nq382lyDCql6e5vKyrtwNz3LIUwJx9mk5WIMUIlvQJfUmHrYYWRquRiHDURKKGEEZku2
EsKQxj5oMmEmksgxIW5Y697zH7xYOV9ulTBq4PrwA8808OW5vNNKuR5O+MlTTDQ6XR41eN19upt7
q9sis8lpecBdUD5v5Y2tOoaxkjTQJfFAlGdM1f0b6vmEK+esguJdvQXWak7ci1EvluKvrhEETaTZ
MdTg/uF78YeGa+U2gg54YWWLPxRlrBCZZ8W4Wf17hxVHfV0McTy/XfeAXAf4mPiLMEKtRyIG+TXU
FY8YmQw7DNb/i3C4aLyNvmm4TcjS6wvVUDkBa9zmgI6q7+eHjBoLKhW2CdtmlKSPjZvptxjtvaiu
wr9fFKABg6LO2NwWrvQHeDW7SpleMDEa5y5QkxlA8wluDvD3poGQ8eu2+kx8YTsuwkZ17hYmHcb8
8m+ImsBMjZkZSUWZpwUfPfeoU+C4AglBXrQhqu6e5XrFwXy+QvfZnb6pMUsE+QO0QtIUYEPgXiwW
IqJ8oMQdCpHMSgyPiUppRWnvrV4SJU881ARgmSXGSHOPYlRhofo7pLU5OBgFs/ZkkbPfg0Pgc+NM
GNf75Y1GDYIp18uLhL52zQVvxeUw55nScFgoetq+Ib5DTeQPwkdlUmWO4mzEGPwIlCkyA3hxAgBB
wG1B6kIiX6adgsYulTvjA0Ys7sdRF8HWYNp0lxCKGTw4d32YtkPtSf4YApsdjo5DdJLbs09MVfCn
vzPzp79/nY5/5m9w4UAf4EKQnFBjWgrpFwEpFU1GxmTnJb5PW8JYzLCJzV5DlzALnDCJCDMyaUQs
oeZsUluoMj89lwtgrivdKAm6L2lLXiMRYZitUjA2X+RF5/BjHqpUkunGC0rmWTmCADPy0C0XfUoX
BNw4j3K3NXLvhDq1kDadS6q3MjMZ0g9BHB3Il6ndCvj5T+i4KPezd0UFZsVONFw4iWP/ZvQgB6BC
XfoGpGaF3S4Gf3haGgvT0HTJky2AB42HLkxFqAo/omK4UFp8/EWHGO59jU1BhjTiUzgO19dpKJdb
biGzJlNz2EzufQzmcwe5mtzLvtCo/xRdcUPWALlpVMrWYieYPl1cuTdadq0SPysG+D34guQkhvC5
9FbJAQhSM3QnGRnrwPVxMjXEPNHTjVyYe9TJjLq9Drbu1mlnvRRdC4RsONLXVvC7Tm7aJrxBVRKa
GOgp04EmRsHcWUetZcLg8fKGYIhWhpuSdRjTDqZNyv6oqhEdfrK036SVHAX+DSzJUmKy12H2Jo+K
KEwtkThYHGzNcvNr6qOjewEsN2Z9ZWB0UUDLtxd5CN1TOerjGnNFMLdyoMuDkhRNRA0ZMSqbU4gT
5YULJMSx/dPMpKoYkZEc/WO9wS9gLUzXnZ62dn/uRBIiD2Mgqd8dF5wE6CqZZLgg+WGImYh/HJNp
Y+GXU6ycrheP98s4FFwn/WZWuJhCRTyLrbyT9FhqO4iBhj+d26GXOv504oh8cklI/KGO9+kaKr2S
u9ZyDEdQDWURheDeZa96UDeJueaQnba/le+r9smBkKE0sp3i9u7kIHMLhonxWSoZuiEsske8zqUM
ktENnRxk2eqrTILdGLzx01J/d+ob36fRF73HpxUiPhDhWwh3Mev7iOy9dHJjGQtJmIDChvZDEg0o
TjXBlscKl+Aik6wzATlLngrSRngrQe6m2BSWPP8LlQHPwOeA58LeHUlQRiwIISZ1TRJDk5JJ/BSx
b187jWk3PZ8njmn/W0dNrfqIqeramxDUHBEzp5rYMbQHTRW1oDWYAeSWivROhD06kUK5+GbQ761b
ADaFa5GY8DCwq4wTBadE2AzA/7TgvCKJ8Cfc62FIvs/+VKyHbW9YllqvldrFYjC4HX8gB5iP5xd5
TV/PoXX3QHBQqupgw3iOWuWprsEUj8JxcAmM0s8NehWf0p44G4pFpcUtalIpJ8qQdDBjB/9IbHkj
D/M30AhloFYw7tcX3FI8YiY48WFyQ1pwzb70HNbJbAfajOpZnHhkMYIhjOirBQ7qpODbfuT9uhft
1mZT+6pquudiEGxFJvxyR8S2bQASFWOqp/vv6+dOKNgZmVO9lYJ9iybsGpuJfkxmQYhoB1FTkjEe
6NqfFIlhYhY0rPdVmDs8gcMEKwY1yeyJkLdSCLnpdfnmObtwBcdouKqCH45v6MPOlheBtrrS0KS0
ewBAQW24+RJUfMjHDsJypRa8acscZGKAthBMs4l6T5zIh1R8bv7CGX23Ti930PXZSMse/bRcyGHl
NV7QGSUwz/tTgBmgxswyFMnVo/cIYn6HGE7tmUQ33H5/Tii8NKuHntAVJ6fXl3iqJmoo+MLVRkx3
ltpG8qroe7/bRmRM2VQUnyvBXnrPsUAm40j/j94lQ4inB6JgMUKALOHU+E+s/YGypOvtVjlAQIw2
bcDYd+LA6qAKGvqVVZrA4m15t/zvLT9wH7dBaeCrw6uVyjW+NTXeqVM+SysuwmlbG14mYgzXIGbd
7dCmlyzKiytSz50JmT6dHQE1F+DwJRvQb3cu5XB1kGnItPhj3vg5WonPIyDRCrPFYe3hrkZqlcJX
8eQBzcZZwNbonm/LRxK0mjvCTxX1NAcb7R7dycaJvpufvEYTKvXL0ZL1paiE0yzhkWmSYeDzwfbj
46I4IQkdQnFSvVwgWcEDMoUDfmj/an2qxWOpTt+D4yWL0rEzr7r+ogUNwhJ1L6qMZk6HRy3A1/EG
XWbtcVa9pjYAMtNZuNxhSukiZC1Fr17BSZkOkF5TOAv1i8IkvUv3IdPkoJWuRIV18oBttTCM6N7N
W9zl6pNI+4spQUWo4mSHBmh45U6O+rSp8ri6iqiC3jbvWGCkGw7A7UdEwRetufVDL9Oxi5NKn+oh
aZ59eNCjM+WzQk4JYY8bB8feQD+fjJGWI+IY2eyqMRfqG5PblqqFzB0vAx+pe3eK50zN9dEUGMLS
qTR6Lnfjr3f+TUSuXg4QBq+ZSz75KATVrHrUDaflNeoGNziYnFXGnniZS6r3SHlWD4bOdHAmJ2OO
7jf0lzmHg+bnmBpgwzodjn3WtirW+lK185iMUHyMcEMbO4gl2fb+4CYj01AGLL84/OoxDCJ/TufD
UGOicZNUy+E2SMNIB7KNnkR8U76ego2aabtvkWOa5J4kMLeR+IU1Izmdgw8PB0EZC/K9c9z3feQe
42h8J2A84FJrTVuC6UX2S0DI8NzZufVQQAJsUxYZXqb+TzC8MVi2nmZU1gX3ODAq0smAOziw5SGa
MizLWE6TreX/XvUoSiQBSKzVzb1Cf+/Vk5LZaif8u374qv8OoCuXzHnV9wJf0JRBLfYzhLfQxFZN
4G/pHAzz8ykAzxfE5FLViXzMvK2s8Yv9sak7/LZ6oOaTEV2GjHZZ/qLCtJ+kHiQSNARqd4Rg1GNu
MxNxM5xs2yQrCLUNxPJY/hywDcUCsu0XWHkvLR4znFrVE42Ovz+9bRVLNGwQaLzUgUg7f+3uOXun
YFqmWdSnvUlhr29l4YG3dURu/UaGRowJLcZe2zXV6J0QT0PBKU9a/EU3mLEmWZ0bKX57t8g6or0D
A6kKArJw2eMJeSY1Ir9EU+h5oP+dquSGnrck9hRctmMieqY1YFGq8V+yRCtrdZxkmTuy1fyeLtoC
Gsdt81aW14mdboAmfmuD78ARDHpzwa3QCeD3WcdpW5/6ww+qkd/WIxuh2FoXJH1MsRlP6v5MOqek
ly7DUmW6nAhEojN2dtTzluoyf7coWAdHWZpRCOEBBF+F4Hy1qYnbDJFh8mk/fcHKCcoFxRmIuiWb
OtXC3A0KX/6vQ74Lzema0mnbegEs2grhaVbEnY9AFDQxjfDgoVX8uWGgWYOKIGNB1SH0eHPCbR3i
KuY4z6/gR5+ARicav5eLiWRI8Jx4BhkD1QZLqXu5L8oqujwE0FgoT7HI3PKP02DfOj//N55freH1
BW3JvzEmKj5+xBnSaXGBQaZyjXXWGuThGuCIVOG4Tu1KFgzc6ivdM7ZeWPihrXs1qPYqfRSfVa1b
3rlRRvD46Gl9opjZ6j5ZKgyirW2bJ0J39Igba2q6h54KdzDFfL8tDMdHvv5fdhgSs4bhI4rmorHK
HoxG0gr4ZlL3iOWmfFo2pjvwizWrSx1Z7M9HhqywaQcXFcCpSa2fEtc6Mo834sHWJOSP8M396rio
jK0m3xp/VBcHEWlFbQolcV9P2i3nDAgZgdy6ODdV7oSHCn4SIdXnAtqSuMcfZS7U+S7NPkLHgR1Q
RHyT5QNUrRCHGJSXoCoQqelKL1MFdIBu+++M7n1WYpsw5cpOcHvQZNZ5ZbLfVzE07Ld/v0TXhAes
a54bRfTe5cRNLiH2XRcaG5LSpRr7o7ncFx85tQ1OjepesVPub8HuLsflFRDVqLNt4GlSRbqxVpeZ
45RoHlJhoo6R8OME/Q0WBURjXa8mCQvaEIe+wrrPknBe6piq43o4BhMzcZm2NvjMZ3zM8OCOj5ct
uYtua4g3Bhxtq8UWtiWgZKxkrf7HB5j73cazyFBYvrD5FRO4lCEjzR16mvAz+ZQE2pVz2LASXIuU
RHLWYm9HkipnUTUpuvm47g/4iAJ2th1u1ppxzX+kpN6g0RoHpdtE4R8nA16rm1VP0Zu4vXUf+f8b
x1TGfsp5T6sLQh8hG1UDE7z+3S91ANmaoR2B+1FW5lylGoL3BouFVudC/P0qH+9m7rqS48FxF+9D
lz8JvCQbSW5KPsKezCQIGAuKdNpsG0z06mgoXhuwds43F2XZbYH8eWBQzThrF9ZBuLL2EK0zG39y
/FRNXx6HXpsFw1OKUzwPuV6OPnnP2ood/WPiU/9aW05RAS7Teut3apmw1Wra3xIm8MeNcDgM5ggK
ajbnPw1pjoE8X+7FvwRoVRYDBT/pRTszpiqjEgzvvNnCnOohp+B2HNNLH++Uqlh16srRe+A1PzrY
be6QmzCCyucScatTQPDl6NcDgW1zSwtN06YfRPIZGXqDTLnhsILjhunaM5OfSd1I4sp3hIiXYvbg
2F+evq17oXqYCXeg+cCs1AMsni+KXZId5y1FEaHeqv2u6mFkYXmhOffCXaNHtkHDgGwHBkapxdnq
8EiM50r7frqu0HqqDKKbV+XZOw+Oh3oVeN69SQWiAJ+Zcfxesoyn3bwSmRX4b9X9HiFRRd6OD8rS
NOzBgv3y0UPOQuc6VdvpvJvOOBZNrjfkRO0nOCsZhvRiH19OrA/5xLcHS6UQYSqQ5GdQjVbh8cUW
GNuP3ma5y8r5qwHIWdws3HkEt5P1DX9nxSg23aZUpLRoaxTrWr9yagI7KNgBGBFQuBbIMEQXZ6ko
2/TVSjdqiCGep3aL8YQAsVOE5j9/cm23rmUzgnJqX3zwBqsp5wBjgNzfrMdFenfe9ss4kvzboym3
cMY9+1iLmLjq5SwuKttDb4TBPRSU5Cw13b/7TYJNhX050i5Bgh/MQ6BBGRtq10k/9x1PJ+h6UNWY
z8IKOW9EUG9fVPUMr4iceH9KTNdJ/ZWI9SChpUkxfJMq84hJhWpeO+3WPZf9ji3rvH8WXMRsWMq7
ldK60xLMAdhE1aXILOUtuzZpT58BkTzZISjXkQcl1N4r0n6aXQoUcb3X+BeBJrZa6QHKKLJnre5q
ixN95uek0BgDgL/rB4RjMm1EfbYCGY0DnW+kXXhEICzLawpp+dx0qjo+cni6sZQH71CRUqknn3MA
TJC5xLi6u6sHYhjjixhsK75E0ZfCX+lUd+xFggC3FY21lTOqY45gWuxCwHFoB1zqR7o6uipLXyx/
nhorBwRrKhCoDOJHemNlRtYYCqsvWuTEheS6Vg2cfmhcijCrh2VpeHc1e/zqHQi289BDyKU5J/Ed
jucP/6FE2+KPAcZdcBhV2a1yFFoFvF9dPZlsJZCMlaAJkp0xQgbaAcyV2M272iwQjy9s50P0BYZl
cWc7upwqXdq5/VrKGhNH2eGOlzv4gRKgMzs3WI4GAuvgysLBg7kpFKZQ9RBmXM8qzBMJSJ8QprAx
usVY1B+ts4+92+Y+zClbfs4Nui+whb2/1DDriyKW3KNtZ+15FSMdfaCtEUM+pusQEeFPDjsCVSdO
BYJEFCVAC9L9DaaOPTdz5O5PAPNWk7FbcFScp7CN4bFXxgrkT+FOM14+V3GpZI5Ht3KcRjD39AYG
y2u6mxcMzdFlWfgWgkerQh4gyA8FcbYwuCmEFO+0KiTt7IAPVmnIvl+AfCJVCFO47JZNcXfMvDzB
L5W5ZywOzLhDkADRZCflZKduJTsExm9OdSSJ3zYUqQfxxRj0634Kwzg6cliIj77IIJs8NL54CqxO
ieAX35BfNAgfKCExXV6b4I893NZPpIJGxUMF9v7AkK9DXrfBaYhIzcfYoYOvW3qltXTH/2/e4oxZ
rpsWRoWckKVKaTasCheOG4ej0+t1yyQARuTrtLRQ30A0jvYlSZa/uOtxIyLla185HMrUYhG/aJzm
mdTMwfQGKfxqRoLscAIWU+vLnsRR1hgHZl054MqrpRKBgKljsHyhIL8Ir+Cd5eqHmFoTyLmRxmh/
kfeLJZNehnGgXTt/yvtBNsgZsJFojsjp7saVhfRm7HHHZz4DvN+QneM6Yqsze1F9xt84DLqPffjG
NTBKUsLx3sHhKQKTwl34IN88tLKx0lGZt6oFc15ElVPM5YjNoK3RkKV7O0aht1pByS1lX7wJRBPC
6dnw3p1ZtTviLDwGs19QQ6fI2lG/zAykoK403gg4W2aJ/aDI/CCErhDmu1ix+FsxjxBPNNWxqJfP
h4Lei/n1FfH6qVXoWDM4EsYtn8fLjdeBZ54465fGfo2PaR4ZqgpSqPuF1DIsU7AIggyvlhl0LRS1
mtVCN58j4o2j88Oy8qFd7/cRMeKBJmw7a44sLdsaWLSiH58hHUEclA73rWf6544yTbaNfRRIV2tO
lx3IkqJz5MbZm0Uu18Cp316PRS1TIhmTbK4QspxNj5eA0p8GKS0GCdO16+KSutLErhoKEpwfdYEl
PEQFuRhJ/zqvNUg+lBJfgClepOggjQRE7d19qRMNfI5HnhRIWRADB7OF6AjoYPHmVkbnrachl5Cx
1ZkSDwRiXN5DnhnWY/nKF4nBL7M4ddgBbs54WWFrvgVMOCtShPScXdrR8V6Ikl1gEaieOUdI0m6Y
AcVJV5QvOBOPE9l+rrYaBDPeA8foNlPbHz+s3oSojRZJivty9X2D1Uj3dM1LB26Taq1v+wKNtalf
FNwVTMU8h/GRYkv/IZl7QvT0YAENyVJDfShm+mDh15l5d8bfxwQMAURt99WwL9kaJzqe8EW3Tk0S
qZ2RyJtXcC4hFBdLOPfUBcRHjozi9WM3pz+GwAS9mS8CTL9I3QknV0iHVRIrKHnmJTm16F7EvSXa
8y88UvtMkMad0Y5mAV2+cBujYefVL4jBQs9ZOQFr0TwT3QltZl1C2Nxa630kSVExpc5h3B33axD7
71A39Cp1uYvVge5uT6KugDrTSRk2Z6avpLylKo7vWk4QD6tZI0/O6AUVzQLvRkVtbHy0mroME8hA
IzKOXUpmRqUi6Aaq23S8yHhd46/WbrhzmJ/xUpNPf93d0Y8h3jhoUtPnVNxeOkrHBDCXnV/mLdg/
TA/i9HGmFgBiTsGEjKawVLC2DEFZWwVylprsr/Xn+SRdXReSXtt0U2TxpjyOfv3udf74NBQN8Ckc
ki7v/H8PDW5QC/kyQi8gv9fFiYp23yYVqgiyEkVFEzkThXxeUT90QRIvnqtWsHykCtIHi5lEHhhf
sfpxGgSSSc5D7JxrNg2Zd97Qo10BYc12o3zcj9j24pYBhiUJ3zLkRDoLfZYiyFOjAPxE5hajUDrH
7zP17C5j+GSrzgfanFg8RzxDFzfxsnUYQVYM8vJRai01aWjjmTOx++5ZrxxxtLdJH6XiPyutxrCm
SVF5wYnztvfDkDUPseuMX8VFJg7jfBtcblT/7vSYs8LMaUC2nPHDLu9neWnh9RVWAj4oL15Zw3kX
/xN0U4uAU5y55/QsSIJFm5yA2ssYAv+jOfYSa8USDFPGxjFGzbGQM7GgESZWumUEB8d+pNv7kCsj
djY1c0fO2+AoKz66m/jfUnqD6T+Yjbo78EO3R3ti6cyJC3Ymh/h3CFbl7+hsf9SOfeJk9UEApnXD
jBe4zrC/CZ4A9LkopODg54/YQj62evfifdf3Zg10b1uVnLUzwTtulSV2GA1mfiSrLYLvjO7WGdB+
v0v7t6z2KR/LNenHyrTh6+oDhkcYS+qhQbe0kBsNWilFUR1hNJ1QANrB4s5+X1i+JJifIBoMtiC8
w3aRSQlrSLLzwUPtgaOzKWgPT2iBU0Uh4BTmlcCJpw9pC6gOcrb8F9EAYyPT6yoNsRRFH1V5suAp
X/vlwRleq/mBdLu/o9/BnNwlJJrqnSQvwIc6WQgR1L+WMkTgcfq4OY4uG6GJBko9g6obXgK6qZqt
pUqdfN4E+CHHuDaLvCn+vHezRncpjm/7sTGZKYo7sqrsDPbhArYNP5IbK3u9Ea3HGdTSGwH6VSD1
rmuntxM8xlZlIv8pGT1g6nRSf3Hk78TuxZl08dmBMIUQjBMCm0EqRC93cBgzL1BYfyOTHBe/rVup
l4bOvj++fepU0lzhDH7V4LWjclV2jeNt6CsLi6dtvO5jgPHnKYiOjarqtwNipVOeRuz1/fbQyryV
FV1kuX3Wzgz/diBbzw624LJ7DuDvGqmreZA98rTTI2rqoTo7pG/ipLBhdV+mzdCr3s9wUKbFjF4f
tssMwKUb4dejSgXwEBAhGNPU/JVhhhdpr0QpcZSGrZJtkJv3WlFHOkSDnKpLiyG0KiVJTzpLBIHC
cVP7KSZF/lVSAsVsJqSOXl7y+U+6ulvljHwEIRVkqxDeMm7DC7B28KkMZ8LqZqgRKO+3T8DEenLp
aUeXPwGklNWxpKxyaFHhD83VAnbZu289vRGeoZD0qdCLk8GQdUqJemj7cDo9D/kfI7TLRjsDsZeB
3tXXWjqAS67bG3j6TTgD2KHGuf7kkskIOyNIfKtWu9Ee7oVBNyqub1cS4G3BVrnygv3ZAfBSvtwM
AvV6F1Fjxu/n64fkPwyaiHZ+X4Sa1iX+kWWP4IYMN+sCFlSgXvLlACyx9B4WYuJmcwg1xPp68ytb
kFlCWERxOWiihxEMxMNPJU+0cY1Mpk9W7uJXtWfFlMWQ3vCt1khn0IAj2BtJUQwZaKMC9jWlpSqs
RBg9TNknDoGkdcWc+uHelLJqxxO1zTl1kx7Q0eA1oXCZKqEX7evp9B2We6kHo7pL29UMh9vAsIra
xiia4TJZReQxuj5vrcFVoqx4nhPKu8NPWI7Dd2kTSzXnbk/7sa40DHlGzYmwtE8OO0SewPYXRpC7
gEH+lV7WY251wVVtPg8OdJLoxf84ylGlp2V4XR6tvUQDzB85VlA1Uqj4AmQgM6+Fa2xRF2jx3Akg
tfhVqVTm3XvE5+KmCQ4jxhw/0hs5SvCeVkVspoagN7XkWybNPmV6IOZKXuNm/nWjkXrNgs+xm57/
1FZOuVUsiDlDxHolW67EWVaV8/PZVKBaNaY7k3wDuuVj+PNreY17Yu57a4bvML6VeQ6EdLvg9XNe
lAePnyG7i0SLY3t0jXYJgX0sbRCJQ9XBXBPF60pXc8XJ2pQoja2CUkvTv4QTX1weXh8z/SRZ5ko1
FHiJjYw70MzaoyTc5HLor5A34SCS1nW/wLFBpY/Btf9MtAC9UOeoqZGu/tIvm/ejMVuxRIEtwi77
v8zWN9eR3kMS2c43zi0NPZO61+ZX/USRNNp1wvftcitnDt6AwyYl89qymYyTmJhGu81lV8c+L0J2
E00v1F9DxuA8oSXokDlo8ZgCufW406/9LAt+kPeKdMQdHHl4MmqtOp/sXgEsUazb1plYOwkc7iCe
wixRsEBHjvI8ENo5NQVSgjLPH7RwJTeBFjQOEyLnyc+pVPWzKIPZ8P/VnWH0QJzd5px5IS0iMv7A
g2Vx3gdG2Nyr7OvKzvpviWmdfGfYhnERhQXmWVjYKK/9Pot7lJ2CwsQCl+foGG1z43bUBaHIcULt
Ea94p2ME4u3+x1rAXBm6dOLwmDEdMA+y0bKkLR3QwnQqRfFChZIoq85veK3j2EspXEhNHN8W1dDh
kXvBZYjnfg3bs1bBKJrroeqaUckr1md3TuFLXW78VvqxST9CtJ1o/eE/5LLarHiAgY7ZzP8f+xPH
jYvz9NlH0jM3mogb/SKlQ++dDoLhJN8JBeERIUtpRRZ3f3egsbtK6JDOBsIH3xGNTpZF8WN3lgWb
mnPA67smra3Q+uwL7YTapf16rZuI12BZDSrLfiX1/D7+mVNN5n+NggZNWV+9ONIWHuk0W76GOMSA
1+pchg5E07MxgqIu/cDTRauXPwmVJPeVmiQ0RWNrAjgkDCaQPon3aqmPh7x+lVBx0urT42927qcN
5CeSKqvrH+3gDRMb258YT0D2sH1FPekwX25gJ6knKQnIr6yDju1JrrXWJoNKYbcqOuYQ1E+OU8nh
Y8ti/8Q1ibyVnklZI/rMOS3/SL/pCPe4F4bdMXXZ1SC46Zpdt0WPb49gdGMpI0zZlFqdGoQqS04D
cV+yvMI2DLkI4Qz6qjDXRiVPtvODicE78nmTruTu0trajphelE9cZLVdDFhtNNVjJhHQMge1aEIr
SaiuBRDDjHNKzHrSrrcI/AVj0vKnTE0cPL6rvWd+7jHmK/IdQ5FXuQaj4ACwVDBSnbOVpGUPzFh+
1C68xSXGyThyFb4yQqgrMh1+6hzP+05McfKwswY7f8Jlc+zq7NMtlJbUtLytEACSQDVsm5MmrPj3
p+LuBB0FNLvnkCvkvdMljJzlM76+RSQFyEXpSlcYAsniQ6wN9LJXkkwk492GCO0vW9hIHO65pO57
cAD1ryel1vtG6nEPbgWiTaWmkaet0fbHa/OJioo4m5+QPnIxQajwEaPr5HHY6L/XO08PZbsw09Jv
StqUvQdVxn11Ihixndy5AXjW7xjT9tOrPl73bFcaxaC/4LvyQHScZQ6Y+6tWu7JDsOS8QtCoZzyJ
vXkSetjoEMJDAiXje+JF7GrS9SlrVGCTLoE3b70wRMTw+KTaXguDjQxUYsD0qwjqBRMk4Un+URWN
hmHKdKCxg5mktMm+GanQizy8ak64ZfC1aNUMYV7mxGGrhgOxl0nXH87Dq/UtbQsw6s83zg5GVeGe
uP4t7fwwGH+h86nuw7jPujV8m0yBAdJWleyzmqcbnXpQWw65pAd3Aj+gIk8XiIx6dSiVgaZK/oo6
oah9asqvy095arMSeAvNwRF6uH3ziDKVVT+q+cNd0rHb9+au10JU2mYMUgc8WM8DWmpZCHU8o1AH
WV53nm96mHSTRq6+9etWtKrJEJFZSynuIsceUwgIOscnonz2X8jHwe2uyl4fwv73lcxeaiRenlHo
U2YjFdYaRtSr2esWuAxOUJ8Fzsi402Bm5Ru+/FkZ6dAgS1t/2gzEUxaA31OOTAeQM+o09fAGX7Nj
SPRj8HcU3frwouvJvAf+PqGBrSTgpbV6WcgFzLDrBFWvcKjjtTicH/Qbz8yp+87fXdzyA/V9by9G
G7Pa0GwenTwwGd0/8RPHroosVZwDtN8Re/YbOWV9NTI3veC10xIphO7DQNWUQqAfjG+KYHzorEwz
P0V8YOkq89qgUA/n3pDeYwCVq4VSB6HHsI3yAbhkk/FD5qOdkeAJjNlVvSbvtVS+QqexapTZZuwv
pgY+bomEXN0WniaLS7eO1M6ZVvJmYSMFVnJQIEW5ecO0/cGuNvWqIJ7bppbNDeABZMP4npM7TgF4
/YmDk7ni7QMxelMcYaF9PpqV4PzFgPj3z+w80xYxhaT/Tkc5oPvc9lUVEn0+KZYCDHRFLO0yt3MI
iYNe61fcRUYl1MpCk0/yD+wdFo1Ez753ugjqU8sDlz0unpnVfDmKBnN0pfU3yvF4FKYbxCqNjRhV
St4kkvwX2j1Kio/ETWifFjlvsUFMfORYlgocqm1+/ctluSyZeNBJS9BVLTwGH6PfQ3rtEZjS1XEJ
dErXCHeExNb97vdL+qvrWrvdpl3w64V+sTCsm5Z0Z41TEpe81eX+e1PFQagh1YxXBKgNi+p5KfyD
YnCSQ6EMjtWuf5BsXX9BNNLLDwX3Ak8TJswgxGDuza/LGmjoSfxU5oiUheEYPRoTV9a1JxYwSipS
M1v5/67v3ng8so2XLRWJob8jBxZG2cAiGJNhel05ecnT1DOEDazV3p7nQYMwukJ7ELigxnIu/06s
547gtxWdAkOMEz37MnRJPFgWPGe97zLojxla/QIbK04E7r3gliN+Vd0fW/dMrHVG+OkF/L8vO5zl
TKzPgsOKipSdkkFACUTPQH/XKC5V77y0IY9xtluWN3l5X1qQoIEPDAFcwnPC3aQ3cZERD+0fQYCR
XKOxD3BPx03FI1+klSSpX1K2dDTA+83fvQuUehnBYgc/nFLmB/1EAla/Mz98w3MsbYVqjitBhPHD
CMkLgu/MMcCEe1DR8D2dUKv7B4ySpTa4uS7x4FXcmDOQyFLFc8vQxMqHtqEquE4UTUe7rLdrucc0
WcXINs0SqCUl56o9Id0n/7zyIxdSjuD3EXLU50sivGPwq12fsNG6PJKe1hQGdJ6Z2Hycro3NEaS3
JDihF1I8Lit/xyLkwVgwv+GuTmXJHlhWLNuFAWtFb8KWiSKPb5nm3BI/iTumnAIzzPogbVbymFuy
hwBEjJDX6sX95edwq2b8Ae24VbDlUK0HMy+sviuf3D5y1sA0+cqqFFP5LqVoP3gjJje5d3c1XxQb
WjH6rtq5lRNfZvd84uHJqRV+/9L4jNd4huTDs9P1jmJ4acW4nQYPJE2K2t47TJqyOYZR408oSNGD
v30AnCMPqd3Ywr4oYBRXE/JI9taKj0hiAW/lMrWcrW0E3UwNrnitSESBtT+u0z3n7W4NlS76MDbS
1k9CkBUTdhOuZaG9QQhIQcCyZeg2QmL/i6ZfSpok/3oUMDAzNnt+GuxdkbQWadSqBnxc/Q8Nyjob
CcJCggTYiC49KNNKjSGJ0QkzLXsOVLfauiFIsZ3IqVM6BTFQrEp2octH1zOO0NFcLB7fxHfd+08R
4vygDBq3UgX+IOfIOwLpBdtVNhh+OIlLyCFDpFduz2/CFK/Jhe6ygIwwHvS9ivfWbdIVSnkSU6NO
mUXcDfpI2chLm9biYizOcgJFmUbMpq4chtBJDusztXTZN3/ydlnr7H3ujy5Sh5ClgPN7rXVHeDqA
pJI80DxB0h3B/TAdFU6XAJBSiAo1qxgi/jmtP/m7E3C8UQSfHdQSi+aWt9ifnwYexdExbudtIJ3H
4jVZH1d4CBk6uQciurUzgnxiCLnb/QwotUkowSruTk1mnjYNwNKkQ4UeadhS48OtRjEWcQRSoVl6
JgFmHpEEF2bMWaHySJV9eJW5/kAKqwx6yFo4zXfbE1geuSgbVwIgsfFXNm1uvWaXGLBiVesTbs59
Z4Wk8jZ9xlvbEpPUQMImg9Ow7p6OMJk9+Ihv2dOEMDVtQs+ahqEJzLEgQIxfwd52S37iw+C9Xojb
5+GnanJuQC6oVVrwDzPZx5iflnd8wIWFw7YWFAtM29R7xE4j6np6tPTO8UKZGGmg/1eu6egAzZby
J9fNGxWjc7aLnSb45Y52xO23EDloWnyz5DPKeuPi7w0WnMsrjcDr50hXkKnjLXqfdhw5fDBxj76c
7IhlF9n5EGK0ZmvywABri5eQ5a0vh+5NmsfCVayhY5ZgxNReqss+eUxieBNuve65EpF3ei1qxaf2
FtK9AE0hSwqOxD1V87+xDUSEECygh6pL3yuyIic0wzHaG06kpNPdDbBZp2if8GJJiNEz/P+uA6PD
FWRQB1K8FvpqKPrNegHIrw3a4sLyoDp+dDB5WRQaC8csoKBIS4BVs52Sdj2f1ZOgApLuj8UyVOET
i+CUsmz+0UAHQzNQMvDehhXl7U38T5WlVVk9Bbmd8O5hY06kXZRYbmW6ZxyaumZB9s2yJ1fbEB2H
F4xhX5X0qtUveOUZ8ttxFTLBq9LquZMEIFmjDyBtz5e0wpXrkar2biYWRetfZeNdFQNBTIE2gKJH
GGIQFUC3RAtHf2UmtVmo/ob4mnnekQtH1JtUuXDWvnp5C/QNP3AH8Uk5DcGvHDodgk8/k3ra3TAT
iaKcXy8Dz3pELLmQND/iZ30YBS2VbfOEx9XvbfY1mb6LcmJ4ubLQ3fYkUsz6NfGbJxni4M7/FjVp
74cvnjy8l1vxA9bHVJ2poP9xRl/0iQR12SLQ51kieVCxTsbEHySGMPtnIL5dXf6lappFR7qlqN1C
0rD3xQkAznlR8Fv18fZ0mUnjsYxtJyzyROS9/8zk+6jCQaiIy2W9unZKnOdfc4P6n5LDO/9Cow95
Cc4GCG8sfJ2FpsI4BGP4PhrDlHh6j4Jtqgy2W7gy7DY03mvDorRVOHBv0ciZTw960nPICeK4ii5Y
19pz+KvU2+PFLTx6JVGcHHib6JaJ+nGiWf0yvruhtggyeSZwdOmlmNVYWv0J4JaBi4E4EooUX+Ht
bwwRa2eiiG0SOE0mOBskN0e3aTNuRqVqLY/hiBqAmlWgGmQBFfIAYDDXQejLKlLKwWz0zadFLwYu
HxFw94PdOXl5H3P4emawiGNSNRV/Lso33GUNP1vbXaJiGfRRrIriNdf0zVNPUjdoNXZ/KvAnvkyL
ErbweapC7PwLY+ZDLxyHat+gyM7nfjYiI27ORB+G3LWT/KMaZS3ZRmNyxYNZ3dxBZDUhdduQRUg8
JQaLlYbgbrs122KBipl0OEYo57b1LKh0+ge5QpiNw5e8sHd5WeYzBNP3ZeeyDAWj7cpXzIr4VC+R
RZYih+23jAPKvNt4d0bxHxezsJ+az+LYhytLdsrntuggm+UAT/tNVTLN0WGh2k4AQscojwaqvFVp
E21uQXZNQFEMiYsh662ien3W+Cdy0Gi8WzATUkmvM8Z+SkXAfBahPJEkBPTT77bGaiDXnu+EWhtg
ZjjdfU0zjKB/kJeLmKrkVKdwA/flDTddatbtG+lXYu9P/gl2FUFcrBb28ZKPHScScYM2QjxVQ1zM
aU4jOotKc18bB16ewcFf4+euiViz6tR+IkS5HYT7ZiR+r51zCN851fYQkN1oWYtLnKX8Z5vLIAcL
ucB23yfp5fyIznKt8kX2LfBgY9RcU4WH7YGEHjunyso0Cu0fbmlv20EPzXezUrqxAf0zoOGP56WP
r8OnEFPclZ04aDm9qDsTJ83VxHbhZYx+JobhFXjDYyU8qkexfwkx/A4skSq52GP5iW/5OF4ZBh52
v1X41d43ijaTGXuZSpltdUGaf9EqvuKcVTf/XY/gqzGceyC3tCMSbKWw5AxW1G0PijvcySnHK4se
SWVcsuKWWnGovNdYc4LeHJNch4KCLzAuCmeoO7phsK5ehvo/ElEni5IkKlBOk7699XWa0/DaWPHL
SOovhG6OQHSfftaOeldAjOmrOKGrujRnZ3XvDEIheWs6T4WHsVcTpGtbh0hI+CvTQEy+RRMZuhk3
htHpsrPmjYpKfnr9gEGeMbnkkTzuUJ+M/jZTMbyasjOYnYoBYwI0gQURYH8JfXP0tRQJslPL/U7t
7PptM4xYkfIeBZ8J+Y2hB/kMkjt0mNGTZkfbzMq82KiVYVheQQD49FnkMs8nBg9fi1qRUxJVrKBX
EbrbRfwtzgoJ73Nb3R+kBZiFSXEUME/jCM2RGNYoXQcdkNUB2s4Yet39gihUxExzrQv6J/CQSKB1
e7HUu+m2LyTRDUlirHUJZ8TpihHn4Wu3U+eijIIoUtqfW+2Qhd6XS7U4hDDOaCx23O+35gr5wTRm
25/r/udhqoDHIDQtp9SqcILvz2La2tgk9Txx/BDzPLP7BmITZNtYnbcLfmq48V8L52w9aouRbg1k
OEjP7MTaC7cwvQ9RkqO8anrqTD1j3f79GQ4ZiIY3vwiQv/+heuQ6CGrHYYedC07a+daKDTzZJfOn
2TK++Fyw69Oyx1se5tJQR7a7u7Q9Ul2tNBFlaraJfQXul+5kNWN2GZnVvgj3qwz2I/QgC/knNr5/
7dqtpQBT1SCkH0COZX1Bgk8WHEeO4dop2Lwf9EdI6NSAbdtroxJnXA9zSwLpBg9F/1VQuTJBELxY
LigT8hXBIhDTBxmXjPeLzx63uqbIOOg3ZlH9Ftyq4LA1qI1/AQ+wxSfePtTjRPbRZesh097p6MNg
Lw941xYYZhrsA0E7AORJONyoQzYHiOF9O+t350o9vBJMs2kJQDtJHNu9A87PYlWmNhn7v1NCPsv7
m3ID6JB73+o2m3VVGHR7zbPVyOwFeQ5SJ3Ukw5tdnE/bnMVG6D/xe4TEUi2zgDkpgVuwxAGdAA7M
shZVfJBwqeteDKnYMZVymoqcRTgc86w93GB9gcWXacyyrv47bDXRCaPVuuH/qrknUWKwYT0IEtwu
WOuw8S4BXp8vNM/CHuaIxuJrpiOGhzW4PvkXpDiUEy/YGrMqQU735efc1LnyJMdEeohWwtNOATb1
7Rdjw7ojk79x2RQunJ0yw6Kv/c2/nGUpWLOoduIrO+UFY7VqU647F1QaPBccQ+Ys4OB3IKwL1VPy
WdZQNpb0lK73+efdEn8gN75twG3s0k2RjVcmqQQfr1yNk7ylDHNTpRrygIt4aM6v6vBZT2zDH9Ev
RelzL/mkxcXJGVG2zEO838kHLQj8grjZR7pRoCQBlbO7TnZxNfsMeqSnomCXNMmCekdso7VDEwYE
8hCNxfHhSAACnazwn6vVxILb352gO9LMiM7+NA2GYNeP9MRKYJyy2M5oIeBTsBM03cdSqr8smWhU
WuwhaToqrh4j0t3IHoAUE+GPtIcirA+YxLf1kr7OvHSK8o2ERyA/v2ZoqJiI944stChixfIS0n1E
Ix4KmBH3l564/LcaeTsWZamSxsTXdj1QMuKWa9PzPmV++x8mPkzJCIprX1J0O3B5et6P4U6qNe15
i3GH3ftT9XGYypsPp1ZkVxXyYNx7iHYcKUlTygUPl55qgeArcfLrXmI2E/aNI5CQoybp8MfSbiEv
u40Fs9Zin+Mcd8QWV3ZvuscyVDUszoC1h9mAvd1tcgX/MtlusR6/R66qsbxKlaLfoJ/91iu5RtQo
T82n0w08vP/wFh3LKcg3SnnjGXq+0rCzgn2+GTOIY9uJsuRnB7pldbKG29NsTqONqrh+9AmsKkIj
Lru5DARFdv3pyjkGm5UYS0ttMxARdcccv15AbmihhOk6wlbsTdQwxdUDhk80j4VyL58NEedTH6JJ
sh/pPhTBdz/BaHYyCR3omo8ofzZ7LK3kSRgSQpq6aPUMPQds9BeZv3eJkbGdNWGyeq/q9pwQ66ra
WwYDkr4p0yjKIvTlkmMBsPZmRGnwUU8PuYwC63PPOBiJ+wUy8jQha1B7QYfER3Kq0BpxIo7gjiPv
y+x5mxDWbANOF0MpqOVgRuMNuyb9GhcMJlgN9SOFRhqf1HGnnrYeG/Ljr9AKqdDYbz81nPw6XyRe
xCEluwWRqq4VZDBqwHcW01EHtxqmpnPfHfOd4RbJIhAF7AEDvCqhLWj9zAJ3PlO3nKD533EZdjpy
G/sy77UD6j0DRzUnG2B0EaT3vDJoWQMhC8AbYcLaQFGSSeA2y21cwIVUzUh8nuGHoz9LS8q+FeXj
+IbAItAMRHb+eG6TwN1rBxz7++c6i43G9fHR3mPA7o1BSyDuK2UYk+sjkEjeOpAPqx3SYU5D+jwb
K2ZS4E9deOk+Xrvwz/Nfazg+k4ht5Rt7e7uKncXCLJ7dgANmvS9pM2++H34ieOUMGmGbTqWvrLgw
XxPU0TpUmeuc6+nFUCnsWU7hdmpjDuqvUHkUutndsjxb0d37yp0DKcJs8m4kUu4sOgfItTU+0WAp
bQjoIOpcv3vMF+3tVbhNXOYEqF/NfauigGP7Bq2OuLSvsHyjsfAA7bRJXi4Knep3OhljvNovO8SI
8p5m901kKIM8idD9q0HP3nV3LCpX5T/O1yhbi55Q8+IW8P4qsmc8bWJzYuH5fwl+7xLB6AdPnj6N
+X/6va4dSjKg6FKa1PDBHqL+KziNabiW60oDNXNzKqn5nNPQ1jv3biAeWlFrwddtL13PWsDsEkrP
61qvtR9cmCT/HQiySskIjXi8m7upDEtMIbwVg7+1N88yihBGyKW711ZXS4w7q/QIp2Lt47zESh9L
/PsjbqSxIDFQIzJtHQJ4cky9aSo7akR0HEhY8J9Ug1wflE5IjexDXVBTBWsZfkujmOWI+wV5FpKr
68gksjlXnrXAk76ZtBWLjkugOcAvu4hQvQ4j/cuvNBeat2VQvKsA4omzJYe1Isbou6J6MU43JAua
mkp/Y6tqOfjkd/zRHqlMNQo9ZBcSwAP4DRaYtloZC4bsb/CuMWbC/oZ7KzwUGvKuhuPWbFOAkgg2
fBaJKvlThD82CqWje5aMpTO7BpuRtJdEtfzb2kWflrY2FanKwdplHCLYvwUivDnmzbG+Cv9qohAK
UzKDzRYOGwc3fb7SiUnjopyotcxNZHLTi/A4W9Fi+OarJ7pATjM7zM5arXaTvVbpyNChE36onw1v
Mo04he93GT/yEj43emkVbcydUeH3miYeqiPWVhZ/Rt8tzPx+aSIkLiFRom5+JAP1awZ0Vvd8+dnD
3rf/rbpFeaeW22rech+tzDX2PeUZdNXqG7uc5Ijz/ymm+10M7lZXKG2wiBOPpYAbXiyGH4n4TVWs
pV0YV5TWvaTzJ08/zYLvregAwy6lgq2oEpMuzC6oS8G7CDFCvY3KuQ+vGNVGGw1rh61NN6XjlZpc
G48VlahGk5MYG5ogdAjJABLvB3LDm0CZS5PBzWH5KVRyOciw6IMLIog0CPywJNPJDinUqousQ7LC
yz39vwg/A1F/ojQfdJvzNYQNd4htkP+VTB3hKkiYrIWT0y0ly5OAB9ar9a2SnvyyPBhv90K+w3Ej
LhQw8Cfmk4kDRe3MxqTdv17Q++r5iZ6Hk2P9jcbFN+0gMadknN4ynDBmPx9bospi3DfpMy7H+0oz
oqOM+R3goF0jXIV/Ak01f56Ne7m0Cd9Q13IzWNYS6zVJrb0VBPqOcRSJnsgozrE7vxtOGaF+ENby
2VzrKJRmVYQZFj1ZfMBSoUGKmFvsJueuk5tRM2pevwluI7QWkWwVMw7ir8KLBSCduRBHWUmZ4XZi
ep3yWQzpVE38Dqa4POpvRXTmgFaNQ3GMMsLqE5ri3eCBDlklGZbO5XDxkYGogWQku5AXfkVhIfLD
NCBiv6OaDZqADXqCwF0TKPPqErv2PrHaQ/5qEecMp1KkAMM1w3qegEg83UGm/UVKu8TuTGr9NrzS
90xPfAv48ikp47In4k7/6DoltIKx0v20Jpy9px14w+crwJQyet4Z7ao2SYvv0WsqkE88uFVLcBVb
ymiopPCJjNRqVfZEYuXhskLWe/6dkyDHPdYsCZHBGdQcP2ERAOomExVYSY+OtBebywySxisGbaRK
hasM98Tr3kMmLW0Ulr5fqYBZ9rRKMiD/Vhvzez6pLjFoXWxhjvXfJgCQyTYU0D7ljbTWsH6VV0sd
RgB7bwvpkgoblgYqMAljKLUFnIZ7uZsbe3LTTsjRGaQS6pMFBDK9J7OexDiPI2oNTDuzgUsTbCWF
Tr2SDV4JPgiMBIga0heLfzwMLA9Inhtm6xCBs1S2HIlgXRjlpzcrJK9uFFA1Qvig/rP7tCv7G2xd
SHEj38IfNd725cBpUEKo7KKi76Ck5yhlJGPBJGbQkdo+hWeu/w5fqK3elAowJlxAfOe3+p31YjED
jj070mBpgLt9JwXkETHc4PDpM6q5Zub3/DlHxdzpWaGXR1L6i+8QZUeifqxMwDkt0/q0icnVTiSr
4mPaFLBlH10/9eN4Y10vqmJIAQ2PGNvpPxUnlaiERFWa45o4F+WAdlX2uF9mA02fZht//fZp7HY5
WtFBm76NIi9AKc0h9EMnChDRbyqjTn6mEooKNxLKyhjQJmNPL5cKKLYarQJflkUAdb4eaZTn3LAn
t2HlHJWznRfjZQmFIg39k6huGpCeq0W6kP7L+djrfEshYV/65sWBveDZsz1V8ldv9OM8ty3HPidI
Du/bCIK3IvXxB/FgKlmAUvLfAyAumiE4dF5o1kw7QN70hhGRSgAqY1UaaYO1E5V1vdT/ExfKneSg
In3lwq7H+JAb75fLi0azMJSiw5M0UVpe31yFu9Sg6Z+Wi+5L5dfXC16049X3oupS4qYLNrj3J4gh
MFsT6fK0SRsPAzLMDazAED2ObvsaNbHZjyQZk4Z3/bvKIEZ75tOxkQJqiqaG/wXTsvVAkHU0wfVg
e11wemFeVtrrAW1omOlJoC0rljMYStehggXU4NiH1+vsBB/j/ty6gT8wJRkyLkGwSYxYD2r38at8
ekA+riAWDsf8x4D0zpKz9hnhlufAjPxDEdYFiqQdWz+9YVD2VMYlpk7+xy11ojIemUTNjQAamjpL
RhwUBkjJn5hlhKseAX0bcmYT8pSEtRnKAj+JPq0DyheBmZOqK1t+XHyWfR2bVFDNm1BuzdxL9kod
eacnJxpHshay+jGm0gILSs/+OB+6ds4aLn9soIgF/a7okR9pAi9sHtp/m2Q3FJM5n1chRVOW6jHL
DAEjniealJZ39lvI7DRdyB+Sooql/nZgJGrI6/Xkg4DpZw2oQHn7T4DQVnxz4EGLBj5rs3l/4q+2
15JNzGl1DExWdGE5WQSmdvg0oBeJuTvu62ONy5yQL+RIB8+rG7prfKlZ6EHieNIQbbboshydPbHL
63lywVzw2WNpa77wLbNKUmqt47MuXtYaLGie/1Wc0Leuef8EiooAy78d/qejFzNazQjNxQ51d8rY
l0gjLnetWQonKp32psVzVESMhYGMot1edwn0hTBVMyCaECxdVB4pFc7acsjwMQLCgZ2zWcwM6Wfn
eGGhj6P/XYEyk+rDfypO9MtcJyXrJSTsxjlxLDeCcizeJqnUGpUDXw2ohctWy38vNLI0flgY/Qrp
p8ygr9656D8hZ9I4kzfFS3izdpsSF38gRczsH9KfJoEVxpEO9GIEDBwtrePx4VCNrxA0yEB4mWe1
+95py3wGkPRxAyHE90Ccf7oWdP9E7VlrlweUp+ZEVYHFQWEK4qedn67l8BDndY053PHRmmqOE3gX
5LvsKTLatO3kzwOUFvD1Jtr4udK4ra1aUGANjEqBvMbGzhZOfP68NeXO7/tsPWxy+HznXy3I/gQg
clu5B9q5OqoqDwD0otZi4E+LfpAHLzOKXGdZ8UxhdySsTe67c8BXBZeG9w9Kao84sm3Qxtes9bu6
9X562Izuz80RH+XXLLnejUNiyD6K0n5FtWOPrZ0qohBS5j5V1C3qvO2WDkh1kYcR6FZNguXSpoPF
ND6noM4wOP8tpeNRHAaUmKyXMMSzOEQRKdMRTo96vC4jpVux4dWyJHUG1UeTHqrAtaH+Ipgaoz/n
gCAn8B5iQfTgysez9Irva9zOoQXT2zJNKy3vJuGnnCMBC1Y2oKD8vWrpVIJLliEgIgK7zJhPtlh3
9iAkdUQJQLYC58BKTvuopkzWHRm+yEV9wXpjEqBJeZr4aKzG5jjHYGNWvRlkvmJaZKXngRg/3SPI
9IieL4ezwQX6TJ9M7PJrsiZwSqdb3mMxSgpMFLuB5KiaKCZgnN2fiZ7gHaRrRfGDxa0XrfnbS9hE
0hBD5xOZPnUm9Mu8s9CqlSFufRD0XTCpxMBfKqoFIY775nmjtgBx8l2FLv+wrW2nodgm/k8JhGLG
2/+lukH5Q+4xWqnPBWRxZ6JeUZdp7it1277KxRymCxy68caKwVP2lErwDmxZkUrcvCQNZxL4uUVr
qeo//o+/vQJ+GzhLDB8zLU3+AMGIHu7mL0nXQOkCNRIHF7E2342H3T3zYF6BNmgje30E5l9LCWV5
u0OrG60EGZxOYSgKNc/z5wkebgChZS9B1jDbcJ7e1uZj9yEbNGK14gk6aq2RY/zdrXvzpPsXLOFT
McGW2a+foF3i3CuGlLGzAQUmvumWtAtZaOuKWQnIFp571G87T7edSUP/6lC7890BXQgfAQ9uaSkL
puhLa0Hf1OxVvoItWHAB2n2lxtwEw25t0Od3hq4uKo7RzvMoKNExpi4bOCRVo/hOrX23mksHoEfN
QLfcT0ofCZKYunzPruM/iuCJf3rVpCusEgcPStNcaYpBGZX/LDjN8iZ8mQ2nP8laZK04Z71xaUPY
N7QyLMdM6GVA+VhN8/t1v5i5GJIWTIY38kAYpjyxCBKjEfV2EiKTu8rTiZub0nsxk0+NdfGn20dl
EY+19ElUF17e0MH2imbIPJPWxnGUA+vbu34R6Pi46Ulr3gPJVMl0n8PfSp1P+U9p45+Qxn1rR0ZO
D6KnKtndHY8kixQIx7dO3u2pi8yNufV3rfd5VG08hXWcr4sZZR9ucS8bfnXsBMOkq/8F+HJE9dPw
AhvHbzkRHs5X/gp0E9rURcNFoW3/BU84yjLHlDiJ1uif+WhPtznnGcveWesKC8jYeMriugvC3ka6
bHsrWvBUZz/7u3aJc38gRlkVUbloXXJSdMVtTjwxybAUdMpm39KKsl0HaARe/e57Nz59OmJbytlx
o0sA3AlbGBareMqWv5XVe64ZyhqoyUbtgEPLiCc13JW3y0dD/UtqeqGXzupxMHx3QyhzJWfMeiBy
zr8cd1DwNqrSppZGFjURuU/kgGIYIAyvxyF9/sVb2sl6X/8sygPFfC2yJ8i6bA21ImAeDKi8PgQT
a+IM7bRh9gzezH9LIKfF/E5UqxUNzBLEDA+88Vi5o2a9YCA53UMKE38DfddBTeS81Se//zYKbqLS
pX/jtozxF+/ZsnyPBbgpxE1Q3/78V8bgeUzVA1t3khycoolNCNg1HemIrwsEBRuN7lBXrCNGSMfY
Dgk2F6MtSFhgO4xceRAzqlD7zB5eYQ4HMgJ11m/4Byt147t2MpI7nLXUg7ShdzycGP3vZfietGLL
XjfM//ULYoLLdYDExitwT6vNw7DTEhYy9fCntdfO06pNhEx2pI98HgWr5JopOtToT/wOSD7ostnf
YVJPui3E3NOoZIf9Q/P/2xCmgMsgKyyIGIPs6QCy3YeSTEs/1/bHTR8SmEQSSCQBolewHpI51ix9
CQB4z+eXyQzVOF+/2pI4NNNkdcezSkLtOkvcTjRt+cfXoTuAw1GT6x/1u6bUAgsLsdui109JlSaC
5rkX0JM32gj9whD8r1993dzt3A+ON92lLg5xp0AhX9dqto9l276xAjS9/r8aEMru+6boxJ2TzNHM
Ydzvxua/rCr9iWAUchxni+XoWLJat3r0yEBmrFltk/17Ix9ZzS7QTa5NLfP/k6VhMPprBMNN4eMd
s7HqR9c04reay5hU/fmpGYPJa+0+ZkpBWy6sDqR4BAtG2JFWQoF+Z+xjKuJZtqB2avS7WnAHZ/2j
J4D2I+fCTkspL8ix9AQFiF//CZ46Yd2UWBtqgjIJb+45ioupVFsTjDliH3KolCB6idJVLG1NNYOT
J/Z4vAPSl+113OV520jbRx3Nm4zrdntsFIDe74rNRB18el10cA8yK/XyeI1b098ZDWPRubnmgoTb
le94MuSMLw/l+kP6a/Ws/mRLVDL7bHyoHm/fLKEXsVtL41AV+9pYPrgOLUWc2w2ST6bDp/Fx81Jm
P7hEPcpUGmayisGNGlqGVTCT9zMek8Nu0dO0dMl+AYQD4NGN7y1Yu7cc9Nt8AdZgYI02HTtkpMA8
Ro3bKGse+XsGXjdVKg4Cx87WkbBXun/gdBzHwkxcQEI0+LJBgx4Xhkb1mnNzCmXdfIKP9neT/TxJ
eM7+REVIwpmqiuNJgo+MXDATEBjIG/L9X+J2CWRbljg4hx/ArlDL9EpOfmBMK775rQIq69RM51Z1
/jrkIu+rA0GQ72RErnw3TVVY/WTo0eN5qQZk5W2QFRHlMY6tPpfWBsy5ojmAtASD9SD7B+Xqt581
gAIzc0msAPThfcN1W+ylP/3v8v306sKlvJRxsj6KBIfamcPDCVC0rjPul7b0eBLyeh8kR082wopA
3iN7IgJgU6e/MdCYEBfAcJ+Z1z0HbuCzk9C+1PCsanskp8Pv9Kce1k1d+HmckGM16z/LDFs8JJ8l
ezkPy6xo8pJHhW6YyAKlhtKwCy68WOChkQpnPhG41ofsiAdPt2V0M7BalQyTpA69g2GsWC9QY1Ms
bckAinpxY3VqesF8CkWJ10SxWcFo7fFnNAnSljt7Boe6i7k3/H3qzAMCTjQStjN4rONsynCVREMN
WcCRBd4Gq0JVac+LqH1LYo64MeuVK3MLulWJDaUYG6LR89+6+ypp5UdfEyHKurW4tRkmO2oBMHL3
MFFFURiEB3pl7At0e9arpBYfGFUHtwk4KxYm91TxVrAoWAhtzqfGiUB+1xq7/e5H9bYu9yhCljQ0
XsGkm1Hy7UHWixfuWUNxpk5l/TDaQ9+3AbPYOMFXiUdYqsUbxDk1bQyVz6NuXkGcoIC2aLv33NDZ
MKwQHMvkLcHXVG6gf6qKqfYS0POKtCGyh838EHaev72C3i+BU3F+XVzRhTzCogHsGXqs3C97vggl
nQIv8CZxL8toPi4mU4+Me7KDZ8taOmlewt1neAHAKf0FFpgmDfwJeO8IENcphJNUcje/3K/3VWPa
U8ArBcSavZlBZGOYsMCus2qbMsH0lyGaf/3Qfa7XwNO87CGzP2/jXsB3o/mVMe4yldjrwp5nwtS3
0Ua8cMqN7wLsxtLkj8maUBlMNGr5EjB0+BZ7w9Q3y9R3SRi9ONHgl3KTqiSZ+1i/UIDMhtzFEONa
9+0Hkib6HvR+bKrmm7mkGv37kyNTti970SbsOgBYOvpwP00fbEuVc7BGbYimZAyZkduC4/gYGeJd
YhzHKmJI3JYq8McXnxUbbEid/Axitp3tl7D81C0tfXqoEcEiSrtSOVvFzlm3uszNSIp4iU6CnpXI
EWi57HzP+4HwoX2leYCH0hmJuiBeBEwHFd1zhbHr4VdjJ5VQ50o+Fg5f17ysWlRWNgLLxhixbiSG
05wAR8qsczFik81WCB/IFUmHw4mH80gwI+aBwYpXP8HDyvauIDn5olD7HSPrXcdZJ/UKOkKWQLwT
1Sinj6uX1heg1NCm3u58jldO5zlezCVbzAYQunVi/to4SLymL473gdVaJ5wAX1GmIdsADssfGUMo
lKKl4TuP61ZFRcVwL/lCI0No0a6HtPSKJtDvc8uy6HUfI5nK2sru174/yuoiap03vII2hkx0WSeY
Fv/zkC/t7ox/PSqbG2AM1kvJLvB2ooRp91w1FY9djiiZoTzoyJGe+1FlVfjt4Zv9CYC3YmFS1eUT
FFYkfVcPyR/e9yA0VHgGwsnu3ZMOvbG+4q5JLB4jLZnB4J4yBSiR1doE+RReY0Dy8UMiGMx1N0IL
xWCtynwjl3jDzaE1Wo569xs5D9e+LC5TZqtatLqsucgZxAFJGBAb7WZUoplMYw2JcRG4diwYQHx2
Qsqmk1q/ZMenwblJHQ01HCiNgibspJ/maJ4JVD2kzaP7JfiSzi/zLRlG2IouXX2e6Gu59zoOoWgP
y++bkOt0cySiuQJx//VoT/nI/JPGFsj1u8Gvs+wFjFQkJ0KfBSLMZhzvRHvaxCVMMLRhaimC8Yxg
zkXgz0Vs9femxM6+HEynxvyXs9aqGiYsIgwlgQH+wlE5ltJcH+gTo86QkR/aL45IffVf055uPVT/
obwXjbcdcfx3of1CXACYlXX3pYZT2ONmlttBH4NFW0gJeqmjlGUOOa15q0ML1nPLMIa1u7IIKBo+
GHgdUGMKJsC5bjWaVhjyD5rz15y2XSWoS9Vf1Huyr4KYYDXQf/tJnEquAehaGsx4JQAZea+YePKC
95j77gjRs1YJ1cOkBh5oI03dwIceA96P0JElsYZx6E4ocoYIKjEXuF8WeucxFpdmrNCxufsEzi8t
4PW+LpNFnWP6giRueAGmecpvW+9c2finznqoAt/vAoPIA0XtZkECSGJvoHi00uiS6JZoJ1TeVkpt
KNpXPb8/Vy4L1UsDKn6GyTS9/thuAL/tK08B7QmO0ouSsbWzxlEn9Zy2Gz4oKEdxUlKvjouqH1pQ
Wy8weit6tVRv/iXDfAlGOQ6v2i9v03HhFZMilWmIeumixF+hb9HFick9c2CmwTdrnbwgUoHN/kql
PWH0kukZnnLUSiCY6S3nOlo1mxcLfZg8JkUr7tYwJzMgc7tCfUznjayYmPvRaM458unDCrrGIpDn
SqvAChGDpNass9RhmTJQruLeI8npTLsxOZaNXVmR3oj40wJFJdgCj/ABWbNIcLPFeIpq7dapKs8Y
zg7Y5HrRKwniWKp3JtyUVGAy4lIDAFkT3mT+/LO2ks0vcMyT2xberZuvbSl+HAWcq8KHZbNou7y/
OhDnG7k/J3a2ySbz7+DVMNeCWinvQtAP/6lFedYOZxRVxsP0vPoHSxhKL568doDMldXF7t3XZC2/
PAR56ggskFnLDy/tQs1qOib4D+GF7sqRJY/sDOx/ZfgNb9HEyQHTbpTabezUxFGJncVfTNNclbgd
nbYI6Gucd+vp4pr2JC+/HVbeJTZishEonXkcvMIZoBnAbKLlf0aI73NPFKGMPL1VffFe77U7qLns
cGF/gU/amo59tOGSPRnelRVEiMBKM17rLvt2lhhlYJN0FVkkqY5i6QwmT9S/YdR5gAEVcWFH/lSm
Kp8sNdgs3cDOmcAJIRN6cvMWfCt8uPGYl4SD5Kae16ODYUm3RWZ9jP1Tx+ckWpREB/EfmobDWin8
dEjmd8LQTwX7HvFJj4BdCMEFrxUwEqub+X9o3RG1ojssUmDYES7Dw3WKQyX4qvs4DqjoHU9xbXcW
ZtQqDeHrcklSC0I+INTvd68NqSsGBLRWpGfb1ckfUdaDIk9hTkcBt6yIa5JVhQA1zM9IMBTSXSE4
myxBNjtkNaR7oE/efv2NI3zy4xW15Q9uaxA/a41K9wfNIU6tpEdaA//vinrqtGgoQj03eLPNP5ID
VCxUsy6vROdB1ElVvPJBUlKtmHRSNKlAe0Yp5MTKIbuhmmJPjdvH3nBG9Vwf6cUrZgafhoKOwC6u
3/57R3dA+BeZBQr2i5NmSo6j8VMTprKlkdL2walFRDcwQFoN37aRMVBTbj8VVxavdo0TZ3XIEUz0
4DcZHxud00nGADezMgaltz9O1OW6NfskEN0zGj1nbTI/iye67CslfBDWuHK2nAjvOFucu4c2TIyH
N2VtLls1PoAkB+vqh/MkDiXM6Vm1mGgQQpqxd5FFX84tpoooeEeJCHau/1k1aOM+V6flI15Yc8C+
ptOq+D827bYA/JZg/yUf/rZtzGR28KLeiBt11AEGqr5Uu5gnSPTouUFbb6r2SJBEncmAE+n3YDg9
cK70KL5L+Hpr2IiXvdoTMWmzpLmXdJcYycRH7ikFeJrgw1xy78dWQEeuSZWqOelMwQWK8Ns6jFaP
t98jYuK0TfEPVtlruhNHDX4PkKr/WKCnuHuKCbSA7hDJBARheQ9Tjw0xDs3ncvnHi909KsdnHRzt
hGkUnigkp3RnJwkPnk6IOz1UXYSVqPFm8dOb6XAZZWMCX981wqBcg4QBMAdfaQkfQLehL/ZJlLPd
VfC99YiJucb66hFYAIs26uLXYpakTOM/GixjVuelDQvGRxyEW5CRvjQwSIvz499lTsuJqzAwkmzY
KpHYu4P9WFbAGQPjkosA+4ZiDbu6lT3riNFnJnTK9NDxtxo+qGkeA0/Dnm24WjmtsvW5YF8mNrnT
Aj+yZHZTNh68cXbH2O/2V5m0fh+8IOagUKO35dVyN2GDg5HIz7EPc9LqRBV3YtEmJ34H08iAAgaZ
2nmJOb6ctNU61uc4ic/qGCEZenGbtYDttgBfUTxjHUY7aJZB4h6hh+S/ADdUuPU4H+tWlaFhPZNq
tgEpo/99dJUNZn+Y5k5OgG9bAcIm43ghU4W5sAkPhEc74qzJm5RUBlhx3w0Qq0q4EC/RqWhsSHXS
v2I0PJhjcKUCmPVgNEtuhPo0UmszwszwYYmaPMwd56QGCepEvCFglOfwW/C5XU1eN/N2mzK4YCTA
ml9xHDArM5h1CXm6Xjbes9u/OWkkaVUdCzj86/iGpTDTjvmKqmVVnMjWF9315y2cVtwcEN1vH8hu
kuRK8zyCFCPT3Ki2dYBuWPZ3yqhOCnZS3bljZ/+LgPUjk9H47n1zQruFwGeS63xnXK6NzFE/MqXw
qQxOegMq/5IQumJ31WYOUMeQEHHaKPhP1PSqjF0XR/Zbp1eIknuvtB2K2tB4a92mEV0T3wlbRV6Q
6eTj11IRdje1npf+6IE7XSnoOS1ryim/vnYALkhu1ze0Xl1rgQOMfJRrM/q2bPANsTukx7CCaV47
KiVSUBHmXCjDd04iP6ZBioORLafv/Z7aEL2RJ6DDLLJODARDj3S2kfTG9Qah8OyQF1ofAO1Pr/60
EewIbNngKwfipB+mdoenVgG7EX15FA2kaW2yUdzO6Nzt7pY4VrWC9seT3x4Su+qZda8nzi6mspxh
twDKaAH/AHQJbmctYLZEuJSH1s9LylCb8dPRFgbZaF5Azh7cNB67FZWCdGDDif4gp0dH3vfDpEtY
1/MEqICjmGLC3zL9V3meH3hsAhunvsHESuKW4nsOI3VOdLRY1/70k7lXQkPbeAJ1H+LGs4NzQ6nU
Qho80AWRuMBrUGM2P3f9bzf9RS/Wk+wgc3qlwKDvGmPa/oSjZa97+/EHMbFxNJ1ta8hyyAprPtXj
VwxTasdkeHUvASJ6PKdJ3s/gG0TSXfi836oNrBsJ92N/R3zxCV6uWKzyOj+anPnkq6MQC1ZOgR7/
nQ8ugfO8HcKZYFF1N+vccmeDgA7dJK7iHIoB0a3jg9KYCy6a6N4acFEERcGcjNv25EzUGooNgex5
RKXYkpM2RJABormZ57Ojh+Osq58B2JS8IA9khcCNQtiahxnqphgEudybW35UsiZPDVxlKwNObEAK
WrE2tYRtQJXWKfB7Qju2r8a90Sj4fYZ1iOxefFp4kwZrhOE8q467BYj+vljYCMTFmsyUhwt7dbWJ
nM71bhhiA3RvVEOoZ1d/FA2Sn7aF1HXu4itXb6CPr9PpUfmfXdD/6VSbQwfnId8PtceJsws76Snv
mKWBHbZeDfcavwzeZgsF/JOkZNaGkrzQZveOI/L6qcTrp7ierALnkm3iV5Z7CFQYQVfOqU87wK62
70YN1xjaW44wWGWTDOQvlhsjnca6b/6pkRNt91JZXhVIbuJzr5c9d7CVpYaEMMF7z53oYXf0boXz
jNLnrEXpeWkKUVk287kwQqQ9JAmWdnatrKLzmQ2MhZ45CalxgC4BtXmPWzcbPcNSNMgkQGetkG0W
nTjpMl0SRxK0pW7LuR0IIT/9tT9uzo72ifpjGwZFGllauL8fk535FVzWF8zd5mvxFfUsyuxOpbxk
FKvuXD82B7BQwrZe0lr37ldPxWGGToEZgCJvnhrBMY+VFU3zmHBCpnTkW4lwI+rS+YQspO7Bqc90
Ag4LMRGl86Q6nGo3pdur9EbKJdOkQrJuzDhDHL3MUpkIwtdMC9E/d+7TVETdW9ydeN3EYMuR212R
tsMc6KRMi6ZenYe+69DCP95vu0pRZaexPy1YNKJa10zMTVCiz3kU9AKFjn/YYRtajk6JuHR8XBwE
XTMWAYNTC5JmIvMK6nrvBZCG59+Ay+mobBRTkLsR32sqysZiRG1cop+YCj3D32bTugGC1/NDMCJf
QEFi56YupuoJWZ3Yd7Xh9vmE8qXCkPPDgKxocV4lVAzfEwMNIbNFVNlOiL0NkuDliyzUL4Ez7jSI
O+ro5QlLatPpz+F1UIftJHyBilxmRNSH0o+nM76uIsG36RaP2mabIL7lSzLusWrzeO2XIkgXXwkq
8jHpBD2ywkXwpIGzqKNhTZb8RbI5x6d5oF31v57Gc5uQUfYR5mJqQVFm0HF7sqZPRO6brT8m5cpP
yPjlI7pQm3zjzJWmAt3veTJNOvDzNLrXNp2sY5TKRw3S29iQV1Gsuv26Vz/Q1qJKFmtSW+r8+z3l
U3PVYtPGbbsmw2E9E1ZPSeXq04h3L6Yjnw9KPWwPezn7nFz9QRiBcgwKZL+w5e1U6YWhPJ6XPpgt
FRrm0eSQCQC5QbAkYS610+QQUHA3x1DA4b6g3EgaSG3YjFdLBUFoVUq47R5Q6dSJy2l/9GdIourz
kBpC/V2qsn4ykzq4kbfU7pJCzsc7xtDpXv66bEXr6IKpOspILO3idC1isbtrx3NhauNM9V4ovji/
hONRYGWNt5J2M/LoPgBGWnr5mU5eTYvZPTKJ9HCfXZt81CBi8/wZKKZnqmd4ET3YHzGR78Jt3CK8
iwWeYmKs852CFfKB0mpB7ayQ2CUbmSCeB+Rq5Oj8oEG3zzzvm8kQD9pIonAHXgzdyujiORk7dCEP
9hxnVXYpBhf6A9DX9sHavHYHDHLhB0b0n+US0qLv4YOaVoqFmZU0Mw7HwhuKOjTJw9s81iOONtCF
pvyy72rW/d90Yd0AkYwF6iHfOayP2mrZFG0dNGTJRu15+kN07eHzoOkEPMzt1sPPYpP0MSpZvhGp
dchNYOg43sgejeW4n6C5BNIvehJ7uwxk1U7d4pLLxEiSUbxibgSFHqZzvDrR9w9R1HI02KyRhWT9
xkn14cGT/WeS5QFuENNrbgPii5W/FWylo4/DfOCDvXkJGTgj8xekAQ3MoIlTL/dG8OrhL3cJMbdH
5KOL7HVQlPaSneLiY4EKF7dtx1jtYTaPYD6E3kcsr3KYM5GZy4rRQIFRyIW+RbBZWjhea7+Qf+zy
1dtPcdBeASxZVGjALWsQkBtDubWgaf/rIrlnwp7oWPFSg/CmiY/8rlgpRMBFTUJJW8HkDkJDGFuJ
88HpdplKVjKD7dBMOq4jKhOb7MloTOERTGMA7AZDYn5jJ/RXtU+ewJFwx4s4txQed5263r3NU89l
zXL50Cyp0Uz7zIh85Yove7AdHuYY+829dElvBQi2wbomxAoSVby5NjD7Db+RsiD0mQ/UWO82SKl3
OPPfhims1MdXuPfrk6agKMzGljRs8sOYebkOQpF4R70KgqppKhVI3sGOCmU5c2IMtEgtqUDyqSGj
PlKqYHPpT0U0uucDIL4wN4xOEbKIZgmDyrGSLJmQRhzXqzBf6eEPLCUlNQKTTaPbMqRVMcSVWY9b
pjQcQkvMu7Q9QU8vJj8W+JeinrH/vb1M+hnn3QmTYVYwKswnpGRAjrgqDPbu3fR40WSe2U+3Mx4j
wE1OanSArhFilHSeX7C4Fnu6/BAgSGarQ56PhEIO5qUXbjfLp6kDq9M+qzsyfOwCXeaLzKPDJalG
5jZOYiO3xM4e7x6zBKu5Mgox1DQNb+siE3CwlgBvQn1NRklIJqUMKxR0NPf6kHNVVx7NfJuCQf/L
pfJ3CGJJ8PasiSMWsUerBRO3MdCZPLwwlQopYfmZagnMTEoA8dLl0IxsF4mtZvn9DBcXQJx9t5lc
jQr3yjyBtu7Umo0essZcARjjLfbaTMXb8qTn4UaX+q7koqyoWNtgTQKrDjr+ESJGGTglqw1wmyCC
bEKhICKBVBxB5On+0uf4AI41YrmCDWYR+wzix2F+DmJTyT32Bi7kbWnrVoCMVwWNS1UXI+XJmDRA
pT+myiaPju6Ru1fGJLt71iABmIjb3QXWNvKs3BAz+WvOIr4pOjLGvNUJmGKlwu/xkCFbyN/rr+RJ
UWkH1m7l2G15OWTS8/H561XBHZTQ8ZBVlEQZDwtFmc2awaqPZLdmVGJHozyRPnUh+hvZcmsGVvz9
14IwvR8Hz0/73mol2R7Fa7I3gomhfL9clc8dMQiLYwG5YQ0vsqamoMpfgaYkv7Lylw02RSXrOx6D
NGIi5YY90RBILDJtG7pl2LA2+2wVNEcQHwoginU5ax89O0KwrYJcxV0GYVHrmm6G5YrvZRAkY+Ob
Dje4tRzC4z3V0oL8RL+THqkviVmFyhEgrTRjbT6V5fCBK0Y8TMOfmzCyhBPeAy7bSobBGFMt6GGM
wAGGf0qzirs9gNnyPkcZxRm7G3ud6XDdfsMuwGIC8jSQdZFtUzD3UCmUceC2QY+tgGIyTHJjjgaF
nOWPFJ/yUOAPc5zfC76Ir5AMzVL0/JB0dYHcavxyV1abROiQvr2zIMS8GxS4jJ4UQgKbLkxdWsCE
YGTvapUJzmWn7ldbAcTf6hjw5I/eYDPb+wvw65TitFMCbh2NJ6WVhTV42zpm0LZnjxYFP7cRvp72
CRn0hiGw+PvLjiX/X9ffVtbdDm6tngaf869pfybmg6RxWBqtbUsHHaqaI5d6Wf0OSiVY4+MbGnaJ
AGL9gUsaVLs8vkFjafkfh5LtJlMnYb/x0vGQFf7KO7m4NRqH2I3XbrZ9mVO9zyj5Kmd1f2g4ZzQ9
0IE2nhRDWZe+rddgJudIUubkOzf0E2RhIfPpnXHUZIM4b14RXxBydxW43/zMvNghX+zXRNCtKcE/
nk4E2WvX1ksegF9fdO/k9glIYu/tmS1zqhqMZDyx+dXpa+bQVqb7s3gSA1n9V0ohUD9L1SrHF9/G
JGo2b0FMet06sEWT1rh0WBzIjqfHI98xJGFMv80pBUXKn2lknp2GROAk594LEOrIokJGbyPnVsRO
M3sNXBV76M0jJ5munAUkYzDiI0PnOHJ3uyXQG0RiA1DA/sE2R32rxcJsNu39yjcbvDpZWYeX4Xss
v0Kskvlvm2BCNhGAJqOJTP6Tyq5c60B7uEpNFN5gG7qUQB/AGGbP/RZEg76UAm5Gmv0XmfSIeA9L
uHTbU4RdwYs9BrgBAGKG4S7/p4wdrCMy/3Nln9GZZ6GeNjs4yAkGYYHblPyY9bpa9zA8h6wtDzh4
+XV3lLZn9ckc4kmzgV5EBPTrYpkYsGUMbjLb4pTRTU2YS8j4RUQZZma4u60ds7cJhINOjO38a6ol
YpRpU95hJVja+T21cHSekOZpLK8it8XdEOvMnDMgTyTgtXJMxUHrItQhQQafYp3RVcdS5tKIzIUY
1fnvYob+V545YdNJtnO3hd0HZO8bNtlWTRCoyJuwAyto3g+ULt4pU5Mf6Em1F5Chvdp6OO1k8fTv
Hu8Zb7r8p8UDTIBP9X3gkytaNthgQPXGxWIVd84GWpXWFQ9YNudUH2qsrbFlx+EbAOFZm8FjssdP
JihEADjnZVQaereSEJP8W3dJAdNzlVGrfHwExK2HUZpCpMJufSiL6EUYfzqbopt1T7qPsuLquamK
SSlmn0pTqUfZAJk0Z6BSM0XtUYM0AkimLSO30eFwvWAKX2OIbwIvyr/wYf7p4PNa5zJDZqyCk2n+
n0rF4s11v5P4ex8szZVH5FBrOPUwinq9Kz7nvsb5m3Bk5sQx2whKngC6vqVlVJdb+ZUA3hJcDGch
e2J7BAerS3Hrb1qUjkDG77l2hM/cx0yN4B2hfHjkxt/YttRglwVrrFcO9fQ1PT8qfzkyFbPcmgEi
w3aD+FA/lf2ywRu917TwKKzf97RKQZ1PRJTm6jd5nk7ppHwEripqj/xfLzoAC3pRc6ZGF81R9m7x
BO1g4mq7qE1oD85WC1x+5zuAds7VTj3iJB5x2genOlLQWT2j2e1GYvGkVincnIRrQ3Jn5Rt3AocG
X7twqaD4+tRE/S/lltwwlFsQCsMOvqWycejo68Z+v5m3iZSImL8tdT5Zl5bCQVYZM3wn778y1m7H
wn9EST6gUosifHh3XIRoLJts8qmuww40bQtum2V5nEFU4gEa/woydeL8hSmJ2oG2jgq6ITiGTKb1
fue5uE1Zny6i1M4lHJMFmgAz6lJ8Zaa1RF8agBa5qx0TSMwggJaVeoD7Yry6NWFLsxnkF/3IDkd7
WhsFc8esyj9NA/YfW30cHhxYALYCmHDVPPyBlD6ILfTFLwgbAAgHN1ojChZuZPZXde/4gbTSFSRr
bdNtWYPRk35JSHUbPWcPKUA0jFeOSiwyCFmNQ+xmziRTTicGMFQV40JFrJEmuSr/CfIJiX0TMq0t
/BjrVFyzYZV+38mOi6fpdwLIykyjSzSuPySyL4xwC020yINHRMF3ECXl35IuJTJVqPlJGbvTOpjK
Fc8jngsn0rKeB+VHJmpH/S+yPFS5ly1CVoVD1uFgvMB23CX8qKXzGuYMFn5KvCrp3amGSrpDqokm
ExLJ8L/NkKEz1l3c4ddcluI4lCHFhfGkn03gdJKsJeJM7s2QVYDbaW3sK6BCwtGZUeXRBEchHmsX
cWveYEjA7Sr3AEiXZvOVQxVW0J+d1DxS1Yeh/WWz5TNQZ0PIRp6KhYsKhvRt9D6brodEVNayyfK5
tJnL9mpGzztWHg1owpOwoFJtI/Og2Tx/wObJKCwav6e4Nb89iosgosrGCYI656CIlJkhBe9tUQai
2zEpT7QCfkxc9/fttdxU+qr4kyiUmB0EaEsIBOkywlwkAbWjfeQyuK5SV6UHFBEloYHfwr44JcyS
xn3RPcSOELBttoi2Te7dcfYh72yZym6F+fgzWrxrpzwKCE6WMae9bbF+T+w6MlR08mBIWqvMiazL
6ekwN1IaIYL0vwtiYKT0/hehP/pmkJa/rQ1qYrLfI4iJ+hKSFmqDvYw6P/SvF/eT8oAbWwtr50nT
KmvL28akIQtlnHZ4RqHdDay4/Qg91vIbhs0hpG6MbFLnJixj/5BjlCo60RCz4mQIVhrmYGzEFLfO
BNqSEypNQK2Gpvgi3abgvc/OvKwvweWOM+P1weK3SHP0MzOusfd6YUuyCTjDTqK09STDpLEczw/s
gOs4XopzDXV3fnNyOglAEt4BcGZmlap2YA1o8ql1gHjPPVmfj5s8zqs4sQ/WXgJuhLSqsy2NODLY
UmpNCTuKx9qyad7poEVWTanQDq4idsR2XSniiZw6ZJ7SB3sefbKv1ivP39xcObMgJtJLsrGjZdaY
T8E4WpvAYFonRIFpov2MCmdgCmLaJJmZR8FsuIyXBunyOauCxxvFK7TDLndZVfcuFi1NzIWFqLlh
5ZSj5mR2EFZJvlHCIKwAZGslFUNZNUt+xSuNOA8CrNfAaH0S+Fm9Ql+Ssza+YsU5GtKFvCl3JPy0
xDXUlz6oLlq8K0NgkFLirkp9IA6k2nf25dcv4gKSFKAhDb34/UeKf+l5f/wdPwWWz9OA1n/nyiHd
dN6lIl1XBqfGqx3KMVsnU9ulOdn4l2ssCMWMg8WELuZivkeeMXsqdFDhg6LWXndFZrlhXVdHs1wz
kB6X+K6ZIn9vI7+2LJ88pARMzdPA+La2kvlIWvv1vzRynhRLLxGjy3Nz6XfZKlPw9+9R4inwfG2M
UjnRduiRWMNbAX2K7Zl74liSUWjqLFfaQ4bXKkok+UyPmrM0MZj2iES13p76r+EjTqw0en01/pzZ
opmC5HcbiclWyf1CHy8hLbp5EmdB0+ISjSzNLXSvSX08OUyt+1a+S1/glSj2duIj+u1a3vPmP8wl
ZDr9x6GUdxoTX28U24LL5FUXGF3uPsaayKkI0S3QOavj8CRSB0X15srzjoF4sg7hNFDXtIKtp/3C
sVczUm1sqNJqxI+q2yCGFfgoceasKuwBjLctaKK4AwRBLRgqxR5/9Pt89k4+FwXBAt/FijGISFCO
bMqCLwlV8cmKRaOTy99BQ7bN+QwWjWrRvWamyZqefVWrMcT7bcd8wWwTv/Xcuv/E0CgfCS43cLcZ
JQ/MfX7SX2iw/aOib5eXElbRIpdq1VdaTyPYOyr6ogwRMTRntMifMpi6O8scI/Ck0OjSedkXauuR
HoZFj6mD2flpEhoMi4wwwoXAnOvKDF2tofmJ32yNOPNf+UqD63hXOeylHBXPECgBUa1/XAfrrPNr
H4ty4kfKP4/Ra6NGZNhWZ5CrSqy2A6AWifnIyWovsx4BuV/77Rn1JoN6AVqLfdewLXveodSXOaB2
fSs58LT1hLXlzZQEC72oUq1yzLtFlF+0r6px5vOPycl2eOCtDtdOLwcsf3QvmvKeIQQjin4KxUWx
Dp8okNn18Xux6szb2Il6CW3ZXLNbDVrSSCixOcHIAjRXOo1R7Hn5gVmR0hgwf8lZi81GirF0KPb7
QYLrnWMtHAANQL+4qrp7pHaMJIp6M8DcbBZvrLDWTKm/gn3papLdl0K6yTOp8lNHppHSgYrRNZ53
4aDKcQNh5XpAuYaOnqeu66Tf3e39YY5fnQ3xwPbRVTvW6G0sZKia8idO3sCTm/PNOgUUDi5zyC+S
e3NrjNZbxqvibPq6QyWzWyNWR3XtqX5QYW5ftt83Wj5aV8LCRRPZBKgkYkbMaolmO9IdjHsb8G6H
Iv5Ej0X1/GFD+dzlH0N6FU7G9E+kLcHZvnkWwtac8l20K+ZhJzm+xU6l1s1Mu4hj1Ron8RJY8pjW
Vz1DANrLfcfz+Ivh5oxLcShbYe8mCP4Lwgz83nDwxT53sNWfar1CXviykwbk6t1DcqhtPwrlKAOP
GXEWtcZ0nE+Eoo/TiWfifoWzenOOBaHxw7SVmHPpUWQ6ujsHKDnT+Rfd3YBX9QuM2cGrDYuxFd70
3tmrYejfQTy/7VX14XNOyNIR+nJ0vqVca/nakZI1mB9yJqkZq91X/xbWRQ8tertXB/z7t5hdNwFA
cTZNNXurRC16CVHGok9TdFWbI9robzeAlsZsA1dLE2LmNik7xTQ+WIEDdRudWOtcrSRaubhSvEoK
RV6zUd9ocTGLipBo/YNGz68LTVNdtm4ZyqQquasmByM1VyQoctic+b7flPlN1mq45DXtS6DSmo4y
xstyCF1A3+xdhCtH0pKdW7uxtim+1lQynJSKF74l/+QDoBVjl6zSXoJUfg1stMRhmIP7xoxsMupW
ocDCqDucwO1ZYJTz0ttCNyo/TwK816Fh95LFqr/QhZeBUHXOvhoCQf0ec/AYJxZLTo0TtuAfU+65
JyZUi6xqP1bcGkUKU8QMWCB18LkrZPreuyPgQXVeS7igDapBiSUKgsscAcwZr4rccmgsrCXVh8CV
Gxd7pF7zCt0An4r3zsAM3OA/79F5R5FmO/bRWsVoEzxglK8ZXBz+cjVGCIQ7qeE9bFBdZJNjXfxq
/+7yiUJUbTsJMvVbsoLVkcu/4kcgyAIIxg+7PXqg/XHeETJIzR4/6h/cO0DuTYBhmq8qtAT6wtlm
jiwfSybu7oUBHm8tr23fZRNma4NQbMjRw6lNI9H1Zu2G7px2pSEJo7/RtEWQ3rC+NrW3yVwxtSSy
mJkCDLP1zx27bFSOwjNRrLcjIx9rfooOcJZnXn8qFBVl+HodTyxNn0X3rvSgaxpp5IzN+3HoRHK+
D6pi8fjIoFQK70/njqQVouZbwLXcyNd0hWVLaQ29S1Y8UEIWOyZZ5YWsPRgkUfh+hZtTUK5NfrCq
WvwN8C40lzF5QBHb0/rbAyAkQ9YkVdOCezTap0PAyFA1qT6kBXt3nQCll0hLKQhFokyJaWqFI9NR
J/0WKxjuBRewgJqywPZBJjg+DlwLhU3Y583fd/rhAO2zKjv4Y74AkX2ZkNwvoe6U0B0iW+CvYeJC
m63J2wfyi2jrqAVKtiBRz3VOxll0SKNZJFN2VZn4daHYiOR5kpR4rTBptzC/ljtGQTJtz1AXSG2Q
6HkckWZsRmVvlnL/lgEjhN1j7mkUnhEibZ0ZEllKvsbCdF65ZJ7Ft8HDqZinBy9kKTqDzujJi4Zl
EIFLV1V1xEP9TWpntWJHJnCsf0RLi3qA/iOuu9tyJLqiFE/pZmnuK9h4D0V9ZfcoII72Q5MVT8u0
B4TltRJp/wR5sNas4JK5bK56mwNmELPKy7tXXaco1XIS6hq1Y6Vie5Pp/3BhdCgyNDQXSUPztXj6
tW0asPjok8Iae21V1eS0zcXJrKWrVOCRa6P+zsbKVcC1Q79AAxvGnecoiqgdQnBDlcNdggfVY5QF
3A60dHZIrI+OZQ/eYlTd4vUHp2Use6ParQkrV6UFyyQ/aH/HYkzPO1l9e5rl3oqerg5JLpmt44Kw
5nKokcCGKdhK9L4PPax9vE3CqO17fUfRdXhzjRoVxbtLEhewiIqdJlsShjgt7DXgq+y31+Nl+N2k
+lvc0j/ZwBIEEjClG7wo97ASiVFJ5tWvIaJ0fEvskLpOrQUfS5W42HmbBBtqKTd9WQN1r2KXvNP7
AQAp664R9epwWiJ0VxmAOSo30zk+xM4aAUA7+1Y5Ni/rB3h5GcIHgNN57DGkPo89jKMvxD8SRyaZ
fNEXhAEBycn4wBqWc14SuiYh18SXCGS+wDVs3PSfHDeX4tf4HJaj03xCDtjvK23StfHuaZiL9BCb
163NsoIuFOdFfPKQEQaT+fMVbZ6eucsZ0MjTBr+4cuOtubiVothi2czDyPbufx88Kza/R8fSoq6F
j9evEUNehoLolPUF3PKIfPzb2QunfL9vWoLHXKOBCG9HqtyeFJEsBT+shkzgMRJ0YD5BIJoRPqFv
i1Mkku2dbiyqB+A4f5luJlhGLxk0Ol8JBESpw+D4P9zE+UCjXtzOxSWDrTf2GPlyotnFE/PXHGsb
KUc+IKqAb5s+divwzDs/xpTZrIj36NpXn9etxNlkkbogVR+y9GPeqMJs/1oyDTY7YtoWqiei5974
KW25ZHUEav4cgmoaPtrm/BmYaPrFggMBIWsBGkFYTRF198GZF7r5EJJ3a3xfGVxzBRUul1+PMVi7
UEu8yb0wgnze3HcU/UGyL0DfmAFytJMPOLy59g1lwnQwRCBz0JH4mtKdL30/e1R5y/7dF4zhz7+C
+BrnEZxZwWeecXmXWaaXov4B5uP82JyOunNqsJ7AIMlPO3w+l5cQkwVT4HWEZQcO0eQeGYmIex39
agr3xBKllTc0nIKcFTrzUJoDfeo1fwotONTAXrLNdGRaQT9BqonG7cFecuulFDub30kiYtrEEEqI
Ea2JbNUCT4tIfu0TcTwKuncr27cOuw1oc6s3OTwfUb+6IL+4xGXnFDaeg9nd8onQhWgt9OphBAAv
+qk0GAdgAO4yt7rIUOfvTQJk+hu71XrWlILHlqeRk46eg7a8ND5RIj+UKrcdCkcOjEbbD0aGDx8G
uoGTWR8IC5T73+ws72fKyuIsV8A6QfAqYRhd401jwrfHkrqmnQHvvYvCrDTbgNtmSwGS3f4hMUUP
jXCrO0rXjhuRBrpw0l6jjZbw+G2cAvCNWtMb4EbengOmPnO29uPDxCMKHE9680PBCtFYAmOAyk8D
MGNWarxcTJO7gnRNLzHZFbZ0BTjnP2o0nvy7Jkj/cuXvEgdfdzsrOYKZXALu2JzAGqAOiTf+q763
iHkj1JFZGUbLDSSfFg2N0sqAhe1lSRNlg4TZeQjJHbwNdbwEg4Yw03moMPrVFhJxnWjEuBOZvEId
Y5goUfGIDClOJKAzblHLoyohctT6S4VsCA2g2BaHJSX72OmHQqatd29f9St6au0v52uhm0cyblby
GX4xkUeADfRFO7ftXlQ97f+SbQcTNjM4b2at0BlRzu+P0d+g8+e0sTMbF7gQNVLThpacZITv51ZS
OXTs+jBroTcmDaTIF6iL/OGkPvC8zH+Kz1Js/W2zv+cEuSyOuTS2a7klshgJ5oyWrKHR1cchN0LW
DtqxcyAriafC+4hevdOs1AwjOlbnwyjQwDcG51jFGQUu3tHnLRmtCP8ENhdGai3xrgkbiEhCwNiI
XLFUnRYA+gswx98tkoVBmuTEDFQpKDaLwO5Gc/o+iK7dqzX2fuC8Q+hAC4Ck5E1fA8hLSK+VKI+E
GFZ2KIoBMEx9XdzPtyiTml7nUomNF8Q3j1gXh/pkFN09w+Br8iY0979IaEiWf9WVzP9hmjNG8Oaw
q7sj6vQzFrhSwbVYVb6hVjO6Px6C58Z6/8N51Tyy6xW0WTilzBpGFyF+Y3bg1AIRuHapaM41WQPT
MlDplV0doGmqSSaJroNR2xQ9KCrrMiAEFW5eK1XO70iOfW1ZHjswcaVs6zmAV243tvQrfRgMiXN+
UlReDR790NCPVpJtEnYETTePG0Bj05Q90GLESX4pFxOndvFvfxeB8EDGdLwNK5mb96EqWZW2aYy9
fe0fEwsjxDZySys/n2AdiSfNrO0fDbsVvPJxtglUGesiQhc2n/au1pQoXGQWndf5B15NidXJaE7c
/KkFFivZUsKr8gt9co2KmRCgXC2S3nIaALy5H5Bo1j6gO7GB+cTJ8wbhzuy29M24ItcdoJbgGJyo
L8tK1kxGZ9k90RwvAzBm8jZa7s9WWgMNHYTkUhV/9N26ysOQJE5MG8t9s10MedKDsjsOT7e1afyL
PYrCqcPifqTE8RuyKe6Nn1VolRKP6omR5RoNngD6ZqALVwUbfv20UaoRbtvO6rZm7qmKgfW/xnvL
ZG0ZQ1z2fsQbCEK0fTskAqi4QBLfVOf13ACdz+ql2wpx/7XonLcYgJDAeFk5GNGbeduWHXB1gZlA
0QZ0bH7/oVdUmIZnXINtDd0xaHice+NJdj9TdPW7byTuNOry3HIkEdZ0eGSLXjbJq8ORJTM0Cs73
R5tguQ6nrhZ93R+toYUAxT0yqBuioSy2z8cX65oPP9DXMH1ChWgOUal+cv1EuGsh327HGfSQExrG
/cp0dEHRSVGE4/UlhvL1gh7hkCTATYBhUomjKUPMQQKMoH3PbNlVAd+Yg7chc+skxWGyV7fKDjdM
zChCJgu9X8QI+hgXq5ZRZUREv77zLoK2qJDzbJVIzSTSTOTNcWw4MrpN2BS7D8vwLH4i+OOe85zD
VxaA2YZ9kT8hFGTdPDGiU3NjjXJYQwpXlwPn2EyDWNGMd2rZkm1cX1W/IKvzg0p5x4nOWrfMVz8q
27q6NUUle50yXv2ZBPuv1LMZpJqzBadhT+1DDWTs+i52rqGIg8kTEGta0vuJ2yQByOSON59BgaCu
4RhyD0J/a7CUiGNXi8Nc9Z0/1UqgUk4TyJTpBGCCiFzBzYMvUvat5v6IlqWN9DsSJo3FPoUr7OXD
ZAkDKINciUJn+hwnGscRedxNU/UYRIFGvK8Ih3WBSa4KCWY8OlA0HN/+b55QDjlwPdygjSkyHY6e
86nW5riT9EwOTFS8v/lo6nQtUvwvj/s/wxAGOLfinxLvrWEe87lxzutkS0JbmuqISkUrOE+QQxDZ
FaUvB7NleV7YW9T2Ajpp56BawN4M1GMuo0lUrkEpGftIRjhdIZOc3215DTqwD1myMTHYT8gZebt7
3M1sLyefRcfJUqaprY/IB+IiUkgHWmw4PvBSFe4NYtxq2ioOVgRCeaKZ+jue0iVwhJ6RLv8hb/mt
GianXem0g1EsNVTBvzXycG+05pQI1jJmjdyrrRuNYzdwV7UORi5WVF86B0YJRDuYEgV3O8ZzsQ2L
+pfe/eS4nkyRycG7RaGjw92rbf1hAglnHmhXDWnjmM+6/6U6jHdbTyLBLMtZR0sH4vgre9knJbDr
UQCTj4KrPgoSCIUvzsgiHGvxgni+eFKjXg/4G8+CAIfZ/krQRkuqcQ+nZ78NVk2mjV+NGQaIOITA
zbEJd/pjUWgF4VIql7iGnStwPM/YZsO9/8Vtle+kROMc0n1/RcmKzJ3PVyn+2CI0EDU+PzT6fk2r
Dq2X4obepEOMR8C+G1As2D98wkSZFZPUP+5ajJmqSrIzyPnPBpT7Crc4vz4sQi2Jd4vA4Bt7b2x+
YkmhSh6tZUnYZqPwZ47j/7xeeMtmYmt+FcVgFIoGWX+uOBpzifSgGL+E49dD4b4yc7G5qxBeK2p7
LZx5P3pxRkdZpPrXsRL8BDBDbRKj66ip1huyIno672Bbq24TXuh4DXa03wEFrsks3U+wKXJgdDkD
YpjCME9MgeYXnGPiQpCRlcis14WN6h6T42bF8pyFoyVBjuWzlsBrCflF60PFGNXP33w1bObjBBO6
oTjJjdf/dg07R6SeNQiV9Vsxa6FA6bQqi0d/iFMhkk4Q1aHv3yJhejGDBgafWtiq+jJ7FX+ac675
Oao56FDkmq97CEbbYBe3GTUmoVD+o0ZxLBnuG7eY3WVDMUm50ir9oTMvMndy+toKcwm/Jtq2u84a
yX1Avy9V5mS0fo9M9djhNGaWTzHiWxm9zDjtfoy2a4TADscNFmnHjtb4HSdbfp8LARK1S0HSdp2S
LLZeDDIZQcNM7yDiHi5j7mYRXhO4UJZ9n41gh/gwO0cNSvIw+v/3DfAJgutEuLiMiav9MeqqSHnt
+0HKYAZGup25cWZd2tn3zqgynH9/3CBagmhe6UD6RaUZUqTz9AyhperS4p3la4t6Aoaf4mbE9WWe
4iSS1GOIL0dC43XsfE9GinPJDJBHu0ZSuW0CxobqdnlFz2iNLL+YZX/qeUcrq8Ad0GZlPO1bQh0s
NyFwsMJrpoclQu5abNzYA64koCSL6YmQzjZuWDRXUx7pCnyY4b+JrqTxgP+LY1FF4JOifre71d0g
pyoAj0XaPbQgIqhnqiaXJcfDacbnSPaZqzQM3X6770Hj2rnSAja8LhV6MnwtKk3znLnmODsZ7OWN
pA64IUX4oW6tjimA0I96YXC3+/Yn9XovDXh46Ee2I6r/YR4LsmFAa3zl3aLJ5lSWQ3+kl0+iJm54
PzHco3Doxh/gOoa4MwbVKocFfsJYjINFnQXBIVKBZXC+ftt5woEleOzt4Wd9WLis9GS3DthniIYE
WScH0HTI+ohG3E4oFk0/YWdcDVr/K27M1BrJ0s8M0hap0CHRCxiIyjIilYBDuB+6mY5UuY0W1czI
7MP50J07B2B9+GHFPW01BtdLyO9dxbfFC0OrIdUFN/RHvbCybbtS5YaymY+KgQ9KM5mHTMY2gh+Z
2o+df3kJbaTt8BuRGFyRuJ6iLhXFjuM7+K//DBGwPV2zOBjPh6jPlIvsX8sccFl0b0UPtT7L/CL8
tT8xbpiMma1l0L46TE19LDzT7tLykRlkbvTkxworYV/tbCeC+TB+u0kUYp4NnbzkcF6whR9GGEcl
ZSjUFuMDNI5nhhowmqjIA3rFl706WLgJA5xwnigPg9l5M+xtPVZlXDaQOwwO5/v9NUpKvkPdnSNF
peGrbVdMO8kwvl+Ft13CTptuVthNXlKi2f09zYiIadgGk6DOoWrAILJxSoXakNrb8n84OzGyHa1y
rqZ8iuu1GQvWqDBEPNlR0cN+OL+nhtKVvVYblsuHbntrVr1A8tHTQ2x/wnr6jodUEqbnri3I7209
12iSvI8t97CDs6eTQnnrIoaw9Tg4t8jUFv7uRahoUd2joJC3v0Epw7kgPsaRSv9K+Xtdj9V52xT0
n2AJcK1TKmWaY4VzBvjqOy7h07wWbiJ0tl4S+NF5tw3SVd9SqAeYl8Dh3s2hrfUU4Rz7l11rIl6R
9goCyn7TZhrdALPL0ZEQPu+rv30MeL3MlPjK/n4TL8jqbr2TC3LFqXmtSCS2Bj7ne0WNsGwhM2xn
erhPngRXyU41Jp88SDpVhXhCBXOW00rpvZ5Qik7JCHjNnw6IORx6ZNbEyRP2TVZcXGM6oIx31fVr
D4qag/ClFI4v/pqBSnPY8Qk191MCdvjQaaxC6eU5Uf4/WWkDqLYvwxOv35T7mctNfq3sa4rL+6i7
AX7ZiOBsOzAilHAiKUe0G0CP54DaFN/aSa2k8BzCcdoqZmRT1fkLGkEtIVVNFF9Of7Mv8y2DQ690
UcoS6bngy4NXFqH2nmfnDHYINvMbRwRC8N8XbUL2CafZ3hFIhLAD+2p2iZIhIyXohJmj7OMJgjyZ
Xk+qCFzyeFsFvLZd/U3BVXsJH8K+y1E8QwZBM2IdUQHvddFIO5fxyNpren9adyH9HUFh5oWgTG6S
D3HXM/KCRrEZ+7N2RtR8k7L82Ol3ugWheMzDNKs/hwim4MA5k04RFdeLv6glmtRD8IIE2vrezsq3
0qtqtJXLLU6ZcjCkcjN7GET3NeyeJT9hfqLE2xjZ7GhEDF/ZB57iq21zVKuK8+nKqMGZG7agwysu
ojg9+mlWduJdAdVopeShcTScEB8pfiZ07OMUxgr+JwdL1avZwL83BxUoKARjotFmRRDXn8UA8ZDA
+k0Quor0sdi2fGS7/EIiTxv2kMq4VjxrZiBWqw66+Tpeu5j44kXFOTjZWuwBvihyUFVvViJc9pLp
4qLbMUkBT6yK4v3hwh7XrAAmesjUKJTZZHgtMQih8ey3vn/JPjpiLCksJSgWFiwLqSE2BMuaQwSL
al0ASHo5CGyq/x0lTwLcPo/Y0Puw7DFZU/6y+CtzyA5b2XUPSI+8Hj4zLzsr5YeRROxLNGjdY+d6
RtvgJe2KFbVX398KI05f4F8uv2V7bFh6491t8z9hCvHaSsNa6vWBBHoyjwtiqy2/DcxzVXVaPWe8
uBL+Ic4NJcy36BSj4OwUszKZt/WgYTVIL1kEq6K8hP9pJD98GpDNOGZwDe4UbmfK1lWCl2gsyb9O
1GidhxspoG6DzNPnRtsCTu077OoObACu5cxd0J+E3Gd5FC92j5SDdU1TKrFxuBYSBj8XQSykLmQc
wTUa9s1kt6ZO7s8+sUgguY40g2W5QIRy7q7cl+E3mWljz8G4wHBjBOP3QaN6poKWz9DqsrLGXUhK
gHZz9QoJvuUrEgaAynv7HzWZ1iI7qiQwx4g7ED546nLUGOGTQBSQ2KIiVaP0bciXfeyjNwTmU/KV
wV96h3B2zEbut+p0XxKDAkJ/qLxtZRwyoJmKoHg0AnkK6sUMnXfWDqvGbgeUunQh5woU0/AHNslW
jjhEn7bbiNQTBo9qd3xxbryrlzYCuIzkfYECnJXKLp4qo0tzosaqYQ5fzAfpTo4WXVjyTZhobzLv
RhT32M8vt4bsVsSmuIZTwlpm32v+xQbzbxSaDRYuVvaRXaTEMU6PXpQZMVv0IqgdpRrdQeEXnZ1o
LT0YQrxqwq3Bq7U2tKhPxnFdf2CJykbGY+RB5cbrv/xYoLkeZ5Q+r0LGyaA4I6oy7MWvEUlnhYEJ
BM5spB4/9boStJgPAnZcDoEMwxbQYC2I707bgGOs0tltcvLmtQw+aAyXDD84GxBENF06rxda/w+6
Nwte+QoDxt/BjM6N4Eo8sDgPhh8rGTd7ZAeGd0InEdlTrRK5qQw81qihcfJlYIFh3D64OldAdvSy
XARfDPkvwpFYaWMJP7BrvHaxLZwVMXJXopy3/5ubRP8umJKr2kvl2LKSy8hrk6TUJuuBxlM0VGZs
wecpLsbgfZAcWwzC9v2VtxmtM6qsecPLg7r5Y8b+wu5hQxhYDuY3VCFUMTgmAnODfo3Bo7SuV2G0
Uv7SFShNoC0uUi2GKsm9Bbt7lLi3xuvYehiWRctilRaht5uwFUiS6VJqEPI13qxAqFDrhK0L4SR+
6Ka+6TqNUbDw3aygHDfSeRazcyxpJ4pMyPGvKRuJPWRECJhKHpvHeYzdRpYWDCnmNCIvx2u2t1qa
g/7jtFHZZcr7it4VKsfjLeM52Ra2UooIBYwFdmdJFIrEGuEvxKqniXoPwDHguw5eHzZtPUHpCzp0
ZAe33m+4mQTUGsXvEpLPyZ0mkGdyGxxEmiinf02gwHn+ySXKqjrkK59yLsORMmR5JOP83miTzZfz
0i7bSUsIDG/cgZb+m5K7FZhm1fvnOeQZ4v+yCZvN2Wlx9fQXmnG9439E16nI71z+P7H6M0ajOrNp
8rDSvAMo1JqwkCE8lYDaRUfracPuxKutN+q58XH42xNRDLC/XCXw46R3FZxCZzGkP6LbO16uBFdq
hc45LtlQHrCGZWwut8ZKw7Q6F7l92aUfZmzxCPbze8Tn2s9E82x6Moy++wryrbFWpQX7Sftb8llR
NOQ4JiliY0Vg0jmz+2Rngi6JvFKm9tGh35efTA29FIYtgx6al+mkTdcIUOeSBjMBrEuJwtO9EclU
e0ivOimngH2klUCimQJuSYXGAF09LCzPx16PLecacrOblQcdhX77p1tSJL/2Ua8xPVtJvrUjVqUV
I1mHYxrwktzm6vaTStdDAqvr+AcwPwTBTKSEmAZ1JSD8f6kutDvoYa2zluGNvqBYWVORdBcwwoCB
XiBuM3mLSeLStLFB04iBMQvDfb8Aj83JQF0WMcOywzayAaHD5+o2cPcUwpSmrUJAj+fymRnwYZnK
M4f0sgsksY6KGveYDfZUriThT5+Th8Pl6WbOErqUcq5DrxWQU8GARohWfCCOc2ysve2H4mqIHcxT
xyRIwNSKIya8wz7pYxpcqSxWtyNlQPiRmag0p35z06pQrr8FEldXMrEe2JcnTgNz8SxCscs1TLsp
0G5ptjvVimsRuKV915WJUkosJanA9XI+eCnpOc5Js4LlHRUgHDB81VjO5eVOkO0LrpdKFTo7Rmcm
IOH+PTgvy95gZnDgL4wz1RqjhoBrAjmWQ+rf1vwdjkDAAvBIKY5veRY9qdeg8P2yglP022wyCqFT
vNujbq5wMBV4BsetxqPhjL3SdEn5gP3zghy5XIzTNU5OPbVrph8cbtdBd/TUyw1KxIJscis+cfn9
4jUI6F7KZH70auC4QqgMSSaWUiI13nyj2X0hmhQeHeZlaE3k7F2qpt1u0bpsv8LV7jsCQjlBE47+
PIrOSCAik3t/CEQ9fVthzgkGT3+GEi2OratYGtYuhCINPxrmwW0JHm+MRuNkkir49XnKHLBBQU6O
X9rS8gQyGPEMI11aVzER3fU7FWID30+q08aqWDsfTqEPu5CdBVme0Lb8NZ/uX9qAyrVaSQMxvM6F
5p7rEJ/B0DpHJ03S6MIinFCdAxnkfJ2PpxUE2YNvveyhdodC3dTnd63JQljyFBvyEDvq+X36a43C
KIeyduAdKcUyCOUqGGXBJ7P6S3xk8grOQO7bqspQm7lGIGSvveBX1KtQIkd0LReL3P1XP8EJoQeW
QSXXYU/h+GTYTiZuIxikq2uCea8cpkWgbAPY6VH3uUS817nYAjGwGovo8wCchXOLXh2KQtVkU/rQ
uD7a7gDcT2tFg2aoo30zc2wspa7YJ8bxGjj1f8U5KPhXskw7ndjAsQnVKtfVlawUxgcSgG+rkNmY
v9XuRN4OE+dUziyGhp6P3Yf2YlBlzvI4oBeZT+nKBXeiBVJAJwFDrdYJpZFo1URfbAqqNzy/RsD1
g9G3SGXzrSwn/KtKVwo98oSJDDdre3MtcDYj83bu4/03bfb+2QmDy4Gwq5NeCcurL64PrMzQSQsZ
4PGxS6h3YAuTCjMxnvAn+na+5arSc+p9qN5oYwBdCccpPT4i2E/GHv5vgOubEXb1FJoyoNjOZEw1
Rg1/oJLZ2QwCBhAz7CnG962BlYjpBb5Mxr9q2w+of3Dq9F4dJcpkn+wciJRVkQ6HQwrR//A4Nj8J
B3JfoLv9xkZhAbiOXv7d3qNP6WVHlcAedddl/8i4kikINs4qZBR+htaeDPtFMnq0Ahct5UncQwiW
1aFX0wUQSpONAaIqd3GEsTgimzyxMo4aAAF1WBKAQMd3Eb0UpGL2466BqM3bY0LzUdibRPFYZym/
c1yrlzk43wISoc6wnV1gqyI54G7+jx7cIZ01fv7MZip+d2lHi9CGHjTVTBBoUrltJXmerhv3xqoO
qgQzRMhTWxf/Z5kehXeGbnx/6IrLhGOHZFTynqIGU+1ic+IbYLDgW9nr/0YDOngF1oJttfFK4HOX
rL13c9Ipb9aRBTREiHqAwDVfeguiALQA//EH/cb7Z5Usn2uUvAHTwpyc6EdcHIimiC9/DLd0ii2c
3AMgs/glS+FlNyac4BgCJ/kFiMiKxFlX2v9Q/svMRGKSD2zggryZ8wWrH3huvvek0n3wHcmZHV1x
KvzXkI2cUr3oXtdg2NHOCDyz6IyLhwS+zQRscgwmiVjkNqZz8+XVVWcm7nkUOTgpJVFfh7IBhbm2
DwMflfAx4ZBTrel/JII4Jk/qwZgDGRvNLj90H9ckMGq2YVd9YZRTboTgm4UWXDBx6qG7xVr9VMCV
CXUEWoNo8gsVIyJCvMHrAbiue4xQ7btlb27EHB/qyENzrxEm4Ghr1BbWNIU/QcF2TtL+XZu3DzOu
IDc7mk4fVs/B+OYhvAztRiK7v+Ag5G3/lFja0Y+Lvz9BW495DMnpL5QmRLanlbFpWaQdklN03o5f
Qix0i7iEq5pp3+iMzkmNm7bILZe2+SwrfYoI6rvaf5bFJqxykEM4ZC179klV5JATw7b5fAx5Syro
uo/Jto2BKYTXPj/YiAz3RY0JWv6zmYtutNKOB2HWDX0M3dEWuRxe3JI39uERkzRpCqXZ/21Fwgfa
BhN6ldjLY5aY+Oi9rxoErp5ayUw/8fVlOZRhQUJp+nH0US6IeHey8TvfEozoD38scofje8PcOMIQ
/V2FNnEZ8EpZg7Fg73Vi24E4OTqMe4+ra9fPM2oSrAjHAAdCv7uck0my+zzuglcCM5xZk0BJEbtz
9vd+gIrkx5PrA34foP5xqf9T4OG7CGdA9eKf3RrxDNHFm/N2F5cbPHNiciFWDDe4Sn8bLUBCasHd
tWjWoUuOKqqZt5NB4b8C4XyZgnQdLbM53rOizWdHfWDy+cYi3+vOTqwA0CFlKKGxJF3vvApywL/N
Zwtx6KpXenAT6ObL/VTSHUbmMTARAvg1lpQogRCu2v8RD5dfiXaupxlQrStpM6sL5SjfU2GosBwy
Nbxtv07bBnzME8jVtiGoYVGRuabSIE8dB7ZPEWcQx7Gs9MR3AdqSDeVqfW0179OEKpgFvJh7pNDr
3nYbXmdqc/adWCTF9Yq0asAJLBkjXfMj8h88SM84/X/rw1GOT1KDQa8qlLIX0isKLXUlddyj1CPw
7DkQ6gZ8Ka8zUd/ttsTRo7iqgc3gV7VGRgRKP4VeB8xakBNJ32yMNkzAVvA/p7eqSHgIX0b53RIm
OUuRHz4ZphuDqM7jJ5Hmc/0AOFIO3doi19f0ak5YtDgIu6EOVgbz/pD2NOO04bCqCZ/vOg7nWbcv
p9Yoc8Jkt+eeoh7UgTlb9EFgac/1mcrSTYhn88zzHoThA/5P/3KpcR8jgovJhrlx4U+EoQ3RHRWA
cFEFdc16VtyG4D+RVOKPw9WH8aWAOj2W9EeOcYTYPI5lXjiXwCrpKbQuhxLiS7TApEa6i2usAnP+
Hz/sPWEQXGm4Jk/oJ/UHWC2Q0ThTyZuV54rgMhHZsV+xhQSmbbSZZL4X7NCjt1NOeHYhMrL1znv4
suptfaVCrswaLLASlVysBYkCrNbuM3QQ4IFC3ES9+GXCsMwz0YdDfz83lVwywJeNfsQZz/VaozK8
5fs00VixM1/hWWnfqxrJcebqFtH9Lb95F+wMy4+xDQRQNMkBZOtU6OfwQv6xxrIxHZh48Xya5ka+
XoczVkOob9fdyz2A+0ud0GMcyPe+dcgULHBUgkf61STNf0raDTGqwfR9HRmIoLte9Pj4CVg+WB/J
Svx/TtRi8/6G2Du5q/eY1Mz40cLNG8nrJarUlf8LsPJVdvWkd4EuS9+gSi/cPlfKMuPbBp9EXxsg
5J61ySpdwQkzCjpUfRkZDpN3km5i9qgyCzGdn6zQbgFZbON5QnnCMNd/engJ6BRRWDULySKunVPu
0UF5mUPrNt+zyYYxnFiYtW2sH3gKs2MLpz+RobGPdpVQuizcsTHhnw9xmos0kof8HaiXSHrp+uNr
jYA9BPMT/cooOR4OF+IH4ho9SHHq4f7EH5oDIXugt9hfetMOei3lB44sFwx8x5HKKzJpDBJTidJF
HhoLT1tpq5y2bDtl0oMzF3QGvjBoOoxw0JAFendFBYwpVzxhCcjCTvbSePONcapnY4AZZGX5wzBw
Ms2ogmHRNJoTFOlzk8KH+Wr6saGtmTMvpUrICFKZ5mQig//YirZUcWa1BjHJM3RTxhrNDWItdJq0
WfeRdcr6rDPWGYnUP1MOEJEHH/XI3J5uhSomFpg7lzP70yQnsb7SbeOoq18sOAHrK+JDfVD0JWYM
J1CvzFpSsof6quY5g7IL0w/CbeCsG7eAqcxQ5UxffhQc9iiEdF2nvxXlUp6XNkFBUSafOzNXbJKg
QSpqi92JueKXH7LmBRATvK8CNGvlqQFccKIDozfnwNg6eeCBGfrwammOL59jenFR9pYqQj0JD2Mn
0g1Baaw+h7v95/od9ekRGW4ZUMHn1P1D3BLeWBgeni8VHJWyABBhailwShRXbGQgZP44eKY3msnX
2Q0xsXNj6PaurDnjrEocjG4TmmO2QSfsfBwvWGmy3MzYllo0YKw3707hyzOpqM2NlH19/r4AzaYo
Vh6zNN/Woat8c2ExWvcTw4nxymfXjf92CkiGQAfOtr+klUaI6N4mZGG9lR9tSWHncY1l3SaVHKbH
djz1Tj3ucDpK10/sYzmh163pIuLt8a4t2sMNpgAoyb88tZYN2wGNN0tbMzWrLfVK9nv7tZSw946L
PpRzzlZXl7hV1alAq8JlXITtazLAr+7LlAV32zdP6XwK0D/y0xQJAJelgjWNwQExZ+sZvjdgsVSp
h8xLzyfGm5NT/N3Q67Qcd6TvV0Je8YpWSV+8br0wBzZmfzAhEmDKhR2jQlxrlQJ7Lvv3HPxMP4aT
oCTQ2vNTgUeWVQsf9N34S9ZFjYtbFKHw6gndzBC3i/I4SA7R30lyY0eFIotxKjijRqbOueWxKvL7
OKZqEY/V6/5maQd2+y0EycOfMi57TPL8MQjaON5uJ620qmJjsmc6KShEeAwhKc3MwiyL5HRnvqW0
4iTZi/0gOh4PrOJAb959N4QeyBWEN42hIZFxN8j84Mn55+HZiJ4P13+/bjxay/Mun1z8NMDwiZHY
/GV8BQh1nhCiKmVvwDhQA8z/0xrjzQILUmeITgLnE7ww6ByDUNzzZzRyIgrIBIzYVvgnw5VMw/sj
Z/UMHF7Yoc1yCUWd8M3ox0TO8KLY6nEh8HPrHP6zPdBTpnBnBWFAhPayZ8ZhYDkYmkRNWCLc40/H
W0Yfd/2uyN5K2spSCGxkhFcWGkNaVGNqDGino/9GuIIb14lIh3LqSrcS9kkFHA/3cuEKEJPol8JH
znSJeglaYDVzGfr4UdVQoW6H/zy3U7klw7SLRJ/bvvo1uzsdNtsej5FaPp+5Ai36uvQTX6L4CbWL
E5O3uLeoAPCRk1Yv8Hv3OJHcuuKHw0MO+YVIrg/Cv8akx1dVI1E8iUcJ2U1gk/nNkaivB6YWcf8/
b/MakbHw6cL4Z7pz+oVkDDdfO5fbz1AcPN8k4dCvna2GHJvtvhGfOEWI2BUNxBjI3NUNeflmQZMe
caPTf3LhxPdqMkeKodA/CyXNEwzdxsYZC7WGOQorNZgXcUTdOI20IYGTIjCa8IjIaB0eM2Jx6Mfy
2sIiwEmlki8AVhlJ0nTmLOkuwy88qNWqbeXmlzkBZFmOtPM9fNfdcixcI7HzG3RVyeaxzHgIVQNC
aV4OdrXrNhmlHVrNKJRcfLbu0ioit/v/sGFuwiMC+OxJPXgbl6ufz/fWMEdFSXrGgxpOqFhYGTNA
LqyRU/ysucHqJ0W2g4XR/x7A4vI05GEP14ndcmYqjvXQUFAK6NfqoEyXfKzZIDbQoBN22vdQ7Qhj
se4EZdroFcYKxHN++sqV2/iTi2YVlNETs3wqVS1bpE9Kr8RMKSwhhk0RV/tskOdTuW+27+Q9JL7S
ESndI7xLIuGoIWOAzYSZwxR6sKOdFJGRqu6Co9Nd9ZAh9aawDRKLHWeBhojtCBJRRk366SHIazjX
QqN6G/GKVY1hFzZdZgozlpn4PIIRI2wv3J2nl4Q61A1N3HWprr0YuRRQVIM/N9aYsgHX5bAhvY/a
awtQIW8zhQ7nJyQQrDlUhPPD6juw9lKyYiAbITzE2nubJrPPqWMFxvEuOh/XztlZlrMSSKHjEHyG
eSivxAi0ajthH91b/ij0vtC+fglTmlbFkPOpjNIMjABWxlLOKCS0CdtAG6L5sobW8ANxNs/KbIae
Btk/tM9DrUdQsNo7UzRe98EaviyF7nVoTMyp9H6guyvaJ7QTnLcV8UWPOU4NVkQA4jKhjpI3L0pU
lHT7KTW5wXzQFgpdC4wmnDdF1hh5L1+HLIAo3ekO8hAGJFXWdqrP6zQTRqDLVSNnkC3py6YOO/a6
xGsaDS/BJRbUfQtTR+Ie7Ql8CJoZSldU9AVI6IQdWkttlYqsdqdC8qMjh9NRklrW5KLw6fADA/Ee
x+hPjpQb6rs0KHAv3vZlq/OiJSs0ANcSzamoLUbDdaSlEt4QsKJ8gIR9TRNSw+KNPjkl6HcH2Ca/
52oRZVnKN6HW+l9lPEKRY1nwml/Yx/1VZo3S9FunC6TCimGmP+CntV1NJn5e3L3Z0yfMoje73/gX
ZPIMRRxMaak3PuoGm0/0pVj/L3wN+bWXWrB7YfzTH15CUyxmBOJJymDUU1DIGbfTCUUQYF1qRFPJ
uWEPUooMPuoRGOe3GWGxkvgow3ExVEN8NU4byWzimyBhb148Xn+iZfwswfTO5rTWf6cP4z+24ZpM
ndQIgPAmspVe9/WvBvQmYmgPkl3Nc+Vao7XEPKiFKzQpaeVHG9ANlc5FWZ5eaPyZ3ac6PT9Iet1S
w9oPmDCL3BU3QS0u0eMUlgjLGKnkrKFFQFwfm/GRq21PmheZCQWhCRHx0qxc3jKtzADfdRABiJKF
KzYkWvshqvxq7M6privSrFVMtGxTeCjRuZZnTelKxLdKGLbIBb2+h0YaPDAJFpKqQgUWCZudrrw5
+W6hP26ernDAC3mMPiIYhO6u/nhdulyKR4ReOiygLh+DlDA+PeGLSL847nJjBQE/U84nAZGbQOKu
PK1yTjzU/C4k4+FZeEXhcZH6FFtnfZKc3WiDwdMVv3d5Xhe+TcD5reoT5jyHziqRJDDr8vP128mE
gNM+UsoR+QxqCr6+NAhNM5C0Jftznl24hBXKUkVYAOT1KjsZZ4pU76cUDDBfEzjDmH0YgWfaF69E
DRubmPJs+EhYAUGvLBDnGozPVOqjHs2Tggp6le8du0fwj80oiZcl3180Llm/FfduhrS9IDOIcgO8
qaI/tCIE6cwJcRNufm5EQteYGHGEQV53CIRtfYN7ByIudldoNlKwRxu4Q9geSEEC3uETqIBm+Bx2
NYP5osZvwjpDzIriFR/DCZykXv4XFbyKq3YlGU07zHFL/Cj4eVXcpTPaj9xYXaZhzmUecDvtOQ9e
jcR9RBHZW6E7iBqcA3D3COCljxgnaPgUkmOKDpDTXuK8Jj3XoRlEEe3yr7bbouWcAA/ObeXf4XJ7
+Sb9KSg3I3umnv884thLxB8anyxIteawvlceOKefjKkDFSLBW6AJYoBq4PMcMf57jNd7CnvlYNAZ
uWoohMIwsZ2C7rqUNBtRHdnj4Gr10qy96kviHCwr0RQsOt9YmXqslDifZ2RAllnXHot3eZKEXihU
s+alD47n+b4i9Xpp8OiAHq79bIvQugDzTrg3gWzeamOiN1zTEcdzbo1QEG7fOEKLAmOoQfryJabe
r/Hc83nZGAu6E9voCYXzV0cwYrevAnHERr7jPpE6+2FmaQ7gTPIUIoGxFt0DratoHH49LcSqEz4C
nN6sigWXyFUKCOofKNzAkw25p6m5tX28Ch36jSTOp39wzGqxxTuYLjpeVo9ijnMejOulhTH1BHMJ
MTFV5iP0eXTkGCwu4fYR2YIe/trJIc5MjLfQwo30ZL2nqxNiZXWA7nyiFccOV7QR/tTdLHpbKdlk
hYsnCMo7KoOAGS3d0/8yTl/Y4f6Bj8d5FJIkOdl9R4amfQmSo3BR9uKLGPm09OanDhPZ041MaM3W
naOzIqgg8KLvj35wJk5wLAquMnOSPm/E5ZmPQMzyao1OOzC9lVXoBIthgTXNds7p8WFjLtoTPR1Q
0vEj9KnLBkAXG8xCh5aJliWkUVmsqRZ/grl2uvQaLMeVDAjpxtRVcKDSlHmqeTEUkh2wz2EZ27wx
bxShBHSbHsLAo7gvmpwSky7WHn9QABOhrrmZT1SL+/3tLoqd6o9y+ULvyqwsoiwhLpj35yTj5Nbc
6IxU0UUwYZr2t1sy9X3Ly+WpEZrapEY5kWDiTpE0KmcPAsZcGcRJUrMQKDV5VatKmSPWhC9HOt3V
wX9xo4NDUALwldF18eBmfDd1JQQ9pdbU6mf+DesS6+bWfyo2SFON5xOUkSLcKKiVxmsiZ2NKFTOy
l4QM7pMfbB7+VVNM2C1o/KUtY6Qx2wGXc2MrpZgt7gs5TU1MjMTTgLk7EzvVOnW30CoRfiTJ2gPM
NDpo4JXSGYtf4T7tqhDPinyj/FJpF0kD3PShNKM0xHt4WJuJ4vKGRs43/iwmRu3+JecfEcBlnPis
ucVhQIivZRNd98sjGaZN8HsXz5/ERBPoa/oSD3iFCcnruEq/MzMlp3YLN5UNcuGSbDvkxs9rZxjc
2o6nevh0I+fVQKo2Ueah5E4dQaH7Nu4gWSkQsd1p26WsUPcA1U0DRdw114TgorV/MBqW5nCnAg0J
ZPGBDD5DOIVKgXGg3P3uKWMCKe3EzwENTTNMZFMsI3l1ndiuJERldLOBpThj+HBUfWpoupdN9Qqf
NYktKKsJiSsPrgKeiSqEP1LbPREM5zDIDD9zPDvvVWd5TSw9rg/iKLhqwOBuANls6b0XWMLFyoqa
56KaSgAgYWy5D9L8TVWzflhooF3VvLHIfT5h47eeVj6MPywawxgUyMW4Xa1Hw7Z06Y3XSo9H2Pcf
1nlnWZXWNSW8GKr/T14+yfCLjt9tOl74y5ZkM1r46cdrqF0xKpOsWn+LcMYk9ohN6re4pwkcmSw+
cgZHA2BjwdcNvSPKC9R/qTlhjfc1IMOafqnVKIbs6fXuTnYSoQY4/zA5jiidy/1/EcxIRLn4XkzJ
otLPlKRasvo/SWJaAi26vHpWrgiVHBNRqa8OLY0BuSa3w5upOlgYzP4K2ajFS/7p00B0pyrnpKF8
bagg6t1dGm/NBeI/QI0qC19LmI+G1K0I3EJDRNzIKtO7U2IS4w94u6I1zzGK5tJmB8LyzymisGlX
p4QAXE6inFajagqlOBXL63RxeltSHYCdCk9KpY82RrkNIpxRfXA7LnVTZc4bNzlYhqsQaUIwN6SN
zfqXDKxDPE40+VcRlEvp2yW75L2tYaKmBY1vSQirLOi0QGK0qG/MbN8SfKy7/wb6r6ibOWcD5wM4
PVSe0MaJzunWGHemsbLKZ4kvH/5Ujq4irrm4HupUom1auLkZ9xqxckFDt+FhLmOD2ofy3slwpfJF
2iCcbB6Py2zO588HDtz6ao3sgUAdiCFz72YRNCGG9uCDcWhh7slKCUqpUkLkbKI5DvoqkgpILjSE
OLtY3NjA5sDvfDexon82a71ubO52PooLR30QyEEZrddfkZe1oHD2e37uhFM1H2dqAenKO7j/4d6J
etFvLAdSTWpwJNHrq4bW8vghsbaC0KgeLgNT7dFRI4DDshEHZZmKLNaeMA+oIwrgZsZ+IcAP6yRE
oOm4Cf0jUEqMGYCfAzExzHzi6H7v2QTMC64fZVJ8TMVQIdN936+W8FN4GsP66K/bZeg7jZxCrhdw
7M0TCBz7+ogjNDLVnh6Oc/UACr5Hu5tL48KhEa4Ee8tVXv6v0QGNZsIJl1VG2rf7DjsDG2Ibe01J
ymuaycBOZW0Hcfvd2LdvWa2DSIr5H59KKbHQjMO92LwNcn8sqoPlMzBZMvy2wGxJ0AUK0K4tr2xh
EcOJ7mdv4EJLEB4rVp1LOReaL2fC4drIOT1bmuUJ46pKaVQzQ2s8C/Qercd2tYOqzr1g5ymU7ipa
phHmlt5+qYEwNTvVOBY3L/Un7GOseFw27m8gIJRJ95ae9yBitztXZiOZkyaSQSrxwY80M/U1IreG
p6O42kmX8egVVk2j8iNdL4W6Omz8yV0BSvHAJSJOPV/uNTYaaJSwwo1TATecD6RzpVJcpvwRYmWE
OLhD9Fk8L1wGhtCCZHomNZtlvLO8vENGjs0qEgLd3MKneEosTmI6jZw09eVEkFBSs4ubuOW8XWEH
3VnmH9Oc+8RFov4XoTYmShiYQBUsoWKZJGs+8bP90H2TTTHLLuFGAa6EoGT8hGNk5rvHe/XSyfKw
Nr0gCniBudG7G9/qOi1EScEr6+yWY74xQ0AqcBra/tAnoYVKheF3qBX/JGCMIIrGbbSrKqV0uld4
7g8/s62MJ+q7BjygKmBXA3a0GGO8+87oov3kWg2SUPR2CZrfqMTmuTXOsvgFZyohPwMSGuIejanT
ZvQbAnuj7rJ0DXxIE9PKg53zNXJAaNixXHL7TyLOki+BrRR7i6E+b0N2gZjY9SYcYdfQ7uey0SD3
VfeXvV6ASlzF5jR0IMrqN/60+z/mlIIXqvMgGWZqPuh3IHql7CX367AL2RX9cLGKZaS8LPNS6SXw
KVVjUnQXHeZFSjqi4HL9ssUXviLOj5Fo3gxJLtx9QKPT/YJvybanREVLlf17cL6mdjYRUtzsuMpd
snJzB5Yj2hFy2P7Ei+2EEgyK/JFFUsRWasOgc9WYURzBLmcND0x0w3HZ5HC4RokkhqT3B7/PKehx
NGsNKDlAdCn9t1N87kNRqKp9xZJGMG7JZSguK2FG9SNuCV9Zrl6Zt6yBzHnm3JDmzCKB5oPLU9iE
WlR9dMlz+n0anfx3Ykv95L1hXvL+R7U/8G7J18n8ELMGhPID+qf3UhtFbCLJ6lPCqzwdi1AWAmsF
0CxAb1U0DLJI7lR32yjNnnQb4g2BOpH8GF7l06/tY7JSM7BkO+LvapPK+GDgblXnmydQWY8Iub2p
3v0mdKbsEexijQdnjOd9v0EoJIyjYDxq8s+PMsp0fX3dHPFPJ1KFe5wTy+9+hLeD39fcghVgUkGp
Qjlw7Ird0mXtsWv0TGdrWCX91h6ftn8pOObCT9rfJJO65jhz0GhSsK48TM3AiBmVoiDNkYFexAli
lz2mnjHm7NZfDB+sJ1yZKhhRYDIFVKtuDVrkoMAWeY4FHKjxRZVo17f3iqDBI4RjB1ngxwJHw0hx
GV4+Hneq+bRA0ozOVXgJ8Qr0duLsICyoG03kPxId6qOGAzYxs1aaoX3wOFpNavTAu+euWN1NAhjR
QR5tRrbXYysm8TJMliagAt6lL6C4Myw4H+INGCHTYpNNlHIZDg0GdmPK6sfKT+oRxOgIFTY4b74/
q3uJp7RfOxhNPK+ft/2undNADNzChhhdw2mkDGSi9lyiik5dt0K1PtPhj9A/H1LbtpzjqfcYNq8i
RxfSOm8yEunaQWTfpXZJJc+Dhwjr6OycGVF0RnaXNsmyewOFwjaFBBFxfohCFo252fhPZSSiB5xP
6SMkn3HtxFqsL+kShu06o3kfiHHI89IdK65ceGX13MQrlymdIWGZwUxvgQAf7WJOZ94NFt1YnKIn
MM1qYGWC83G7ERoxdAyhkdhLQt2VKD6+2uF1/4RvuyToBQnW580jssJiQwQ2pjspH20fw2Z1hSjD
M8OtKKZHr7qWGTrlHlakgcIQMkoZwYUiKwy67+s4G5K5SdwqRbQSMb4usT/bbC3+ZLaRokB33F/s
YyLETcdSKXFvYt+UYPAiaaaoBPB5/OVIj0UY6zOXZW3SCXozyCdOzWOoIc0UGA+/LyUfCOo1ao14
Uja6Nv9obFCHuiUTpwDClKbP07+8FxgDOLq+yWimLAf3xIyzNyBj3mhjFmWZcw1LeU8DTaMyvhrc
MsCK6udGACS+W8syusZYExqZe1hpUHuSyhz154GSC/kIqGz9me4XKYIOsqeIoZi0/c/ri2dHP1q9
MJbsyM5RhjHMKWBlnbzB5t0/w+KMn/olS+IYOqRfXfHbB2LNa11MiHz7HUy9MDKdLW9uGvyJJ1Co
LV3D9rnEOgPBh4xUM1lRQsZcKJ060yW4xBX7yF5lH9LzsFHFlCUKeyDRpWTLs34IYCYBiZAGhjET
Nn3S8zNRY3j5fa0yo3OKa5uxR9Q5pM8ulhz0LVEw3+bBjMab1qt89LcugDQgUJ8/kVNLUCV5DFGf
or/LGCJkASU4SERhyvb78jLUl/4eMvJseIAaxffN2SRkzW0vjIwPL8eHxqiSr2ZlJoRNgLDb2Kbq
qcSQaWU/adNqrtsaPsrcPYZyOUuF15m5x1gU1FCw9YkjrVc7yCerDmgZMljiFvut+u05eLWyQTUl
HZDSfvxGDaRrAGEojMQMFcdMkBgBu8jet/jwr/zw3q2srszJyyqkJ3Hr6e1IZr0XJ3hz68cUCsIn
lePOlb3KxIWQ9zIKhutZ0r0OmZoW+vsqqEJ1VlWFeOFnC6Zjh1vpH4M2jLOmX0/DEsVuAuIiCxqF
KTU4/m7Le4/bNsAfTri9L6/ylFW3wmjGdpZysJ++ci+/rA91LWyFjcJBvpD02B/aF8MmPCoXMtmR
7naObGVhfGq0hTeqGKbfZVdV4a2GGa/UXyL+m2XFd8vI/END/SBqwYR1zgl42bTw/gs2d/tNM5T0
7spXPSzoI3xEi9tB/WoSAnxLL1seS2ZE4JMCyXR6kisW+u6uxsrO7D8OBRyh2fJmr8zYtKiXuMh5
sQWR8cAHzi9vqYIDb8Ls9rjIiQb2K/Wv37Qa0Skhz3JF0ZQ0nOfbiT3j3AXybYmHUhatPe7pjFTw
MwsAPy/XG6nfxobU+hnqH6piU3RljzauzgadiuX7UmLMqw4B7DcOE/mrM0F8bpoXsj5iU4Vdmauq
wfotecVA0QBuxKO3d66lYxYGQJUKoKEfUVjmAm5EKi1z3y7u3xPlPMkbKjtTo5bz9owSlPjmB0o9
wadEXVDwQwhdtEAdC3/zqMIOmwWgA7bRNMfskubKRY7FjwnZTwpPAqNScLuPSEJ9WLExsVSLmk+n
VNBPowb9v5YbJp9Si9If3ABZbdgwAy+vqYW4K6/n0QnPjbmaX15ge/oYqqZSn5r9tNZz+9bw5aoL
4hPPM9tPWL3X9xGgeLf3MyoXzIXrvn5e8lVboW7zXHmX3viKlLU5pn5UmQZJKz8Kk0K2ysn+Q2vJ
KUZtj2lnayE4v6sKZbVP0wDTbrRwEnhPtW1hJgM/Js1Ho3Vurotd+nEGJC1OEokIa399W0D7dT2y
lkB7MSM/8+uzUzg43OClLVVfrzJfvQAFmjWzn6zFzLWDlH2ZCaJhVVN9dvZ8C7dU89BVjY0+AjU8
2XZq8CGIncMHZVo13lNBuNkByEXBopwySrEb8p/lHY9zjJHkRx2sPxNIDyX54YMY2LmQBQYEDVze
cRhzb27XvhstVW+uWOasW/OUojH7gnL5g303wGlf5DzPx9TlwP1kW/yzBTCoN0Oqh9jItDMNo7Tg
GK1NyQ2RRz1FuKFYOKxAaCqzryQFgGTm9iaVx4/N0mxuZ1LkCT0Ra016oo20m1tzqvFJCU9KV8ns
6tHH1HvD6144AUfUMnwTrTFou68RePT+GzeZ/um0bulDWwF/RCaKbzjXsmHpeYzVj4lY6HnxHPT8
FbW9TxwFRj23jBugqCMGt8AGlkG1XXJ3MxE3cjfio7lDuuqU+UPuHJbKsxHZIh/eoOcA9uOJbxOC
aPEgI5da4e0WBFcM4/2ZMvG20NDxfLz1xNga2h/DXxwfV/tGXs9EOwwXzF3pMtP6VHSGXZ8KJhjZ
tNgK7S8lfkuQF0c7wUJklb7JQhtnwgZ2HDGILS/86jHfJkBZjR/6TOlRMsTDG5h4lAFR7J9vyvTd
uezLeaMNrFPg4EWBTdgo9L8R6e1RPNF9Kcr9SaPQsB5tM3LBOAFlcufrOnLHgpUNNr81MvwzmFxj
TgyqtMyBS3Ky5Hxql1gk4M6zzoCjrg/kV3EqGPzM2e+LkVKZ772NuU28U9BnXopBWee9oqH4dOHm
/A84O0Xu4SOESFL6Z6BicxqtEdVXVqoLdtG5nWqpHBft51B+BhcrX53r3D9d02Wl+uJMhyWTJHfQ
TGYXYWM0io0WT6ZR/oXMX+yQ+tdAhJPOrhJYO/qgcrOyp7CGA8a4IqH6s2YH1Y47o+A3zWquu6uw
Q6vfrGPV1RmFUCM1wbEEOGrNO8d1ujYsCO7HKYH5lbiWSg/LPYW7ia8iZWrSy/1g+GeifP56jT9v
h3h8l7PQm+/3ONyegAbck4/VdRR1ZIN9bsq2N77SqSVgCU+9s6W83BFumoakLCpMNCOJFi1zYJTa
BINNzKqwhAPAx3M4rtthkzR/BM93wpDKRuzoJ8LMKlqSYhjY7B9+YzuipEnNC5T5fVtVC6PUdzti
JwiCuUwkpI2F9FvoVzYTGf8OQ+D1CwhkXSwIn2RVwjftoC0SSo1Np1/NQsXBQsE4v9uQMyCd4tMR
NoWXo8PxeFwLEU60UKiSFV4xtnz1jfu9WXK1AOk9HHBsvIBuH6cnNElLAzx5vMfP0+kLwt8+QFDu
SAth1ebEhQeXWUprfZy4OKCs8AU8DVjQqQnMLvIB8IEdOyHw3o7CwOavifyCxYxU0yzGtferSFsV
1qHDDbdbpphUzHQndggE4Qdfu7FQrUYC3uPLhsDiqOjRiSVho3ro1xZHFbgCD0AYOnly5OiCFBXW
q8waHGP6HBSNhOPUTlBsHglU94+ggfPJIaE/YeWFAMD1hfbby9FG+UY47iQpxUcD0FepwOMuGzXr
W96zvrkLJ1dTi06U7wrIre3zwzqdiBl/OpYR+DpVzuhsB/tQHwceimqAvGUwpXR2HFhFvptvgzh3
Joy0LWsuwHzNhwD7MeukPVWG7on8wKeiGdtPrDXPxyn3dmIn4CoqL3MCRD1RQa7TZjgbG07AxkGK
kfMmdkgmZRdxk7SN2Xx/KswEjYUcYG8s/fxhxK9aG2Oc6RyiSEOWVR7ueS1ZXuDurfZSHVAILAl8
Barw0gyKxwTKOqSKUjvLS14zZB2Lmo+C3tY8RbKS7Y5NSMJnPda5kz70a5A4hI7LsVRvVdrbGkvI
HYe7aCegLvqjrEWER7Qgzh2bOF8CFuV+2r57Fgl7WHRSWfK7AsC8OqiJSv1PFJCPefttrpiKnoBl
fXoEYVNm3Bo74W4fe5TPze+6677DLJTjGYeYrlqTGlDY8rIgZ7NbgHds8m8XbInLZmWDQ111CrFH
Yvz9mNX8laL23bucAk3uYgSDOa6AvcLrrICsr2lZ1hMFW4Ej6Dz+SG1nl7TKIzSb/Z01kNq0d84n
rSFGIzF5RASSudgNO3dPg96eDdQAQIGyQALJE8V/7lq8vdiP7p1FiPYQkbBDtosKtIGV3r7yMDKS
lGHXyry/TRphTkeFW3xyVDQGIBYl4lUNDRqIRe8fgbXUoPe8ByYRSDZqeaBnTbOZfb1KiTc1mVfr
YS8ngv4/995hm+04IboaeVtSiR7hgGqY1D7LRYpNhR+4Kr6/LwygWGtE3fFgFyPg0RoNBSqUeDrW
CuzJIz4IwAZ9ugr8MsUDNKm+u1oIz+3qjaBnQD5UyIFKHFLKamRCb/hJk87qULYgMpGIkFXN9AUd
bmJwpFscBbBnQ0gma0d1lwf8SreNUu3YrFrdggCe3WfL/zSUB8hYkbGPXcxYtq2gm0zR9rabo/Cz
mjbo5x6m/ujbO+toEPDd/lh03DyOuSdgrCb5GvUKH3nISmg0u/+MINsZdxa5a6sVFJhIuNE3L5w9
o73QmmQAgntUl02hES12C3F0WklJzJiszDYffDvxA0B2ic7M4YWM6cdE0k+JZ3MI8UN9pCC/AwfE
vCoVny+d5fem9wS8OTMoC9hkSXf4zeAVgDjnhGTPnp0kJ1pk6mx/7wUf/OwQjZHbaS9VmeP7z7zB
LNWZI0WgpefvbIGpk1QEj2l55Y8gi1a8Hv2Nt0b5v+Pem0l1+uFJ2sR4md4HCQ4K3qWgXt/AU7Ij
kIp/LQUkWSWbcFssf7D6s0gKnqOvjd9K7CH61heAFg9Sz4t6Ga9WJAT8lvl+hlC1FrRzp8ovKCbx
JIzsWDLbJyzVyYJiNX5wpImaEYthKHvCGLSzhUMMk/+KrJE90vVq0LZJz7Lo+KgK0qIwRs7VcbAg
fgEANcfmy7xhI/6RSK/eJ/EnTtCCnkrP0JykSeo5MHxrohwfPUCShCOcn/PQ0jbhPITKS3Gb0vYV
PQEABqAzK0fAk0Ix64DKfzdP6hXwZzGR7nIVX2LsdZumAGksFNqq4kWUIdGcIXDlOdNHeI+3p9Oz
G8uvIwDqxtuHXAUdcm9KgJ/xFTnMBHA0RZcaBpNU5kvbqLS/O7M6jux7kIFCvOxqhumIJvUHifT0
HizAtwCHg5eQgVHQdHBR9vS+HO9b7ZCUaB6GR8vWz9TRa5nLzXIFzW4omBqQh7e6t+t+8GtOOfLk
XPD1/27aVt5u3M8kXwLa2E3gEaoZXMA94VI9wKA/RSOz8bS2uYiuVQp/GJfk4vQ3oVEb1h8ZLUTw
/jfZbO25cyCQykmXfFcmDknIPyJ5cXXOM4jMngJqwYqHvNdCoLBpnWR+X+rJg/17s1q50htGOZB4
f+GCfoKiwh47a9oCA9ujbe+JtwVNipxJlk7Xo/tfPMmCV4x34oNJVipoGG4SEVWWfwY3F6cb74ef
duXk48gd4ceX6x/3wkGPClYIDzmdAg2X9UqQDPvJxaKgRurwzI69LunbI+o/f+A0+dTHXudbx8i0
jLr8x5sH9UiAp5EwVz49PhDZBK6NshZGVadcOr/GUGCzR48XBpukyIKwn/hCturaj6j+OM6ySU3l
RDwqHMoPgSafREH+CNU1mZI0Wz22IonRFcZzHYicxiSPN/rFvGzwudY95j73WW5Fm6xKbAZRvnN4
jJYLy+htIUXETTuzy7e9C0ISOLTiajSa6ATJyEp3yajZwfdXZpBN8qyMvEnUKhWDsbXAhJspTfRS
GDv+JMhHqhhVr0PFxCXIqI7UpRCO7/odVHLNLSO/Vqu0JgFSuMRxxJfia82b/kVT66WKt15ucKQT
vpjS/wdNZYfBo+Dpek7ZSvAC2t270pVz86r4VAPRev5+6CxW1O4d5uHVoX1TRXdotUWkodtW0qIz
RQlMJqzSSMXa/+vW6diaNPyNwESzUekyZcaOb9a41TAdhbVKmxtLzGAj/H9q+q6xfCPiJrhGfXXj
itOa95acoglGkVu9lf/dYJkCP0JNdig4r7XGFguPZc6Z9WWVdHNZZSkYCNiVGO3qpLPx7dpNVZL0
/28HdN4c5xPIHXoJvBK2MQDZU0uJxNcs2ifNz8htCOjiwU4+QA17rT9PvV+pFTqSmUdZY+fuukN7
UD5PRR+xfdksrm3uTMuUYniGUXEl+9sGs2H6WfhYFBDU6aHyaXRpkqIsh7AfJpZr7Qo/o6J4Ybb4
nZKDWtCFnxXO95ZR7EaFy6VPwP5jT+q3A+K3xv5bJuWe6ltyBhfOuCbSiUWKOdWR5Crt937UNY5C
igSfAEsJLLpUvXBiFuBLdQ453MPTtbztNUw0ZwjhVhj1VYfj5hnobokRbPx8oHWK+DpjibZlATRL
cbjWwyXoAHlOoQWp45ZUvMomC1WHI7Xpeakf6VFOSE3CrvOsi19C5iXaK8ILbarRCVPXdHJXyUtw
6pGNxfSKg5oSwjR9SqbkpbeOiYBK4jopkA8/kso0MG83S/O3qfAFXMIMjQXXQHtJaoEYMILh0mpB
bruFrJd+xLp1xzAUx1YI2OnG1vxaR7hJ2OHh6svyHeC+OjaVYKQk7x1cPs8G1rgRPtnNe3AATVw+
+T5El03D7SNkVbLY2s/z3WZGPwLLJTCP0VmHCl1TS0by5KuvRroHcGbiZH6JT+AW6FS2SZE1PVqw
uwH+6WQLfvLaBs7Orjn64jGKSnTAj7pnHq25u319D2xqONzzvWqd5qKQdNhqhiGPVT5YJh5aaB2i
+tPQgzdAFYW21hSdAwZvod1bHm2VFR4iZo9xpB96K2f8SuHx1sMspxHWJPlcCi5WFIBOgbqjd9my
537gVwLq9LCYWAwYb5WNq+x31vsrZbp4jeruNnJHU3J1flDmSGc15m3VVuqKaFIjTrVB2YJzcPM0
U3aflqZ0bjjO/pbAC15kTNy3GGn/FmS4ZF7mkWxihLthZHYvTLDpJ43QDP3BtzBDn5eNDfwbSgDt
EoHQBdvfR3Fa9eU/8Uk9wG3jlw9+kCd3KFRhiaTZaikF+MwrrOMNPLbOZfC3sQAZ5Nwndo1FnlCK
f+anUixugPVLJacdir4edGWZYc2dxhXIj3OBkDpUc9GxVEAN6XrMZ3nJWCK9/qejCufmUVy3lZuu
/o29wjhcbSs6qvoLtpvsOR1PCdejMlMm7j/4nFjmr40ndGzgfu+Hb/es677HoA1ELft0YvkVfEzr
4q7bHvLzKh1lEoiODM9R2Ti2N1FYp8PcREV7C0w7gAlbPpsg3JgxYmMxNAAegumEkkYgpNhRcJui
Gj7YEQVAmbZr5Q075CzIX8iZUuW8Oymf5g9GUlRYHtkPrnAOYiwL3FAkO6Z4p2MOU6XcZBic4C9/
ITZ6ICeKvf0R/+OXLrq3noCzILcB3YUwbQuaLPkf7AojH0dh5TzPs67xBFTb7M2xSdhSbRnnVriD
yhyovXMLO+mO/mEHDZUNsxSE+uSejQd8uUzSxd4LQspl3pDsoirdZgxoRb7OnRDYKZt2QA9TlkBl
zZSfB/JzRAzNHSHbWG09WK1AKLJVJk8LImN0m6f21AmJNMtzLPzhwyk8xLpA913BPzZW+UWupdJO
LulLCawIDgaoaoEPx79uBOQtAjX3asz9158iTwQkotx8+a27NJkLpUYDFGFbKVB90/+1jakgr4Kx
Ocjul6M+7iLCFVazIGGMzgFkmwtfhSsjnvKRs1XBs3KaV+Q5CVnS/ldcoU2jQ/DHBV347oYRk1Jk
J/raAH7sd5hVfAd7tu2v5D9SDWJoOEhXhTTeqDLQl4ZGRYrdTwd6M4XXCIbhQZZ7sTPf0niAlayr
l0hpH8v9MS5nETOqi1uDiqfSKxoHlqS/THiutEjh7QsjvOQP5oLxjJFRZmtVe7MHE59ACZN8FV1S
yaQC7kb3aCIrkW0kDFZKtC6w0mdFWpNywsLDJ1lx7oRsgv/ERcQmtFHd/B0q8mcOitLlezjnnZcV
DPBIQfEUlmz0i7smWt9fLj4kypT3faTBR234JR6P9sc1KwVqc1trig+CWDC6P2guxOV4kOvSToyI
F66BQ612xPFpTRl6oiuj5Md/tgKLgNohNgTeZtLaCuzghg4FmtTtbqw4vwfk+BVxAkgZfw+vX+Cm
PJB0zlU2DMt3ZIMzaD9zNymFc2nrD2ksBinvbOmcY3woGhoIN0/FUm7EZQpk3AzQ/SsvCpe+TsHC
kqTZk6/SBdeUOP2usW28MuMgekDjP9S9T+3hvSP146IYQpfOD9TEKVcG4LQ37dZCCX0xEY9RcH7C
0h8b8lMQ/o6OJhNk0hl0nRedhLyGt6zOgdikpvNVMxjSmKEWHGXrGszxBaQcrH/GAc6LuXCepIFe
f4LE/TYg9hmbZZgIzuGiORKy8krz2Zt4tePtKza/qwVvrxr8j5rdkcZjcAZ7kaOWga3o1GOGMZul
uUkt1rKfAVzfzITkyxal7obiyrGbgWPsyBNr2fdE5xlqBL4uCz0FRsLn91nT/XT/dkUbNAthNtvA
R8qYiw6H5Zm3V2leCnQyOypNCTR9lSmVzz1mi+w53hzeR0DUAPlDGVHfQ08mA96bteYrUqHpWCzf
3cC9g5j2BGrxdo/UDOacZ6/WHGUsRurdPpVvdWLUZ9DJgTDFGGxHAjfmQKb/8ogsNdBawozZ9ROQ
qyhImqyXcHqsZ4KGQlJuVM3RT6MSTBYncMNr2oiug/t3/y3oy0pkOADazp/9zks0V2J2tPXkg0QH
mAExn78b4ePvXgrouHbqqyeYharFAc0H/IXxjvNnb8tyskobpvA/npeWKK48TgeFc7fXkTmq5e9G
oOqBrnk/pL33CjEkRKmXc+LuutKrgbZKGleKUTCsS61BQWe+/Cv8QhWcAfE/BqLG2g/NXH/V3cVK
RHI7Nq30FDcHE/YcVnuAEya5hsbyKW2YtoZDNEvmF8l0Rxk1W72NtARu+ZTNWHJfa5lXVn+p14FS
EMazlh8EbbKgyWcaaCySwi/ieR+Rbnm7ctLJHA1KST7Wfbh2NjO1UZfv2aVsApNcvnw8xZpaJdR1
b/vsrJXzEIcG0479iPkEYXMDMucurexcTdgjti8ZRYNuaJjUxXVDSy2xamh6yQ5V5KphcvGaK5a6
r1D1v37TFynKl/DLhe/hCHPM2d8dEPmIDjGQOH3RGdKRG8H5riUrpBbUBY/IBWEuQfAAlCRN6OvQ
2wpZhHkmS4TU+pkQ1XQIupMbUFEvCOI6AoR0n8AS/FtKYLLrLPvJsmdzfySeQodMIrJNCLxVFmBd
HaNwwcYJHajvbRfJdgGIZuqRIcizgoSBvu79woY5Arl+OEStcu3PluA89tcImHacypYc2AB+dju6
79K8dB06T2JB7JoFY1esq0QF30Aa31MxDDMu63HL8z04q9eWOjCPUwmc2mNzrpnu53/5YF6OUQRE
b+2lVt8tIS7+BNIyPGeg660BEcIVwJdVX2HmyTrMoY0GJlae54iJ2zYxJIlf3ZM0LgxTrOV8Sdr7
65W1a+u7wFHkpOq85T2B4/vKcZW8T6L+09MP0xPHVFQ8QTzLqwPIJNoL79oUJqyZ/LSZi3NHWSLU
urhdDVgZYFCdBBcS4kvLECwvEfu0MmMZXoKGkdU/uOy3jZo8zIZEFAwcRjs3YRUjy1OtCUWb+OXr
EExISgp2HYVdBTyRyIfU74ZMiNU23JO3H5gePF9biHTSCcv5fV0GuH3R1ZAayam5Lk3KWx+bLkjU
QYGZEbmwKBSJkcC2ZrnQCkDtzN1falFL/ROPT08rFwA4ZXNg598b2bhi2s8vfWqxBoHh1Q7mSLSe
3JN5DELnjOmO8xo2HZZbaEbYjZ2z6lpKXXqRRm452jeJcO9e7zhA7LJ8bYz6YYBvXnlc71x+rJRH
0qA9q2WEwreO/gX0O6KuDzsl0mN9mvSazYrtjXnMz33PteqFh1XxTi4LF9Pr3QKbc+Q0DGlCZRJP
M02/9JY9/yCr0/IygZ+KN8sjzkGcxeW1FAiRgv92mEbmGsCx7KKyS0IvR3Xz+NnZjl0yR+cQYar5
w1GQiGJ/hbjq9ynbe8Q1Zcg/+9lDFsfV7UT+PGxIdSu+4l34x7ZDCbENIdHxcYtXTiWHGqQTHtCP
r8G3s3Yt6X5/BriDn1ILGLB8wrkgMD8Wj9LSCGZPoYylasDaAdvPd6HEbyoLqvFTHYXRZgRAPmWd
eOmcZgACcvVnUM1cpdRslpvbApfzLcxfDnkRehsxA+/W57kd8x62RmftGFjffV4dS6wpxgASiLAR
lHO+xIfDkmLPFbRpTjLikIxxJG+wlZ3jpV8VDRbzB7e5Rp6f7sE3uPy2PKk5C2gLUl60VpYayYJL
OHV4zsZxCoPjeNSn19mcoepJnICxZeRPf0o9zrn7O7ZYy+i7Deo9MUG7whvjcotWDQtXHxnsW4fu
BqaGqeNh15r8MLcNCZty/ZOfUU/w7Ts8slXYKnnndZvqCd4XPX8cq3UFEQ7fXIZ6BCstO8kj2W5P
w9USO9HkG3L0VLSc5syvgrkyw2qyWnZRjR+SSd+fxIHyw1ORsVOSbc95o5FkjqzG68/ziYI4/sxy
uKtBXDEW/mhL9xZYOok19438CyVXDOBuJ3cqtNDsp5wxHjZETxZu2CVmnqFwXZB8scivcfoBCNTP
KjxMd7zyTNMj58wBHOL9Q9g8pR2ZnDRJXFyXtJ9ciaeJHxzYVNpRZ6YWKZ+28VQitdRcVSPk/dRW
buA23qL9yv0JzW4TGqRrVVKXu23Cqxj6KHZnPtqPSmtPh9Ex3EWGeDIVqAnBS70xl3maDjD4Iwua
qVwH1oCRGuJkrixwYpKdkkw0ARdkg/rd3YSTOtJEQLKCXFW4s6x7nfL0K16J+YtG1ymcYHT6Knva
o8JCD1UXMytIXEkNM1/ph19xVxCN8NqZL+1Qiuo2Hl6sUO8+4j30+ZjKWYq7uHmh1zvoKEu8PsNo
ixHB8IceZsf7C7AqYTClUkvJy2WMxyBs6Bo0REFDTAq/hMEkZhM5Iv0QoZ0tIBCinIrT2xo1DmQQ
YeynGCUfqLMpqBtTwGYWphdnimojp2l9ouoxJG+vYiVcrulAuPoMDSm5Mmnabnzy7thR0lMAw/da
bgQmYrqp93qhlUSJLRIxFCepvhqudEL6RDDmQgxb7udabaQY/fYmhQ4qiYIajI//Rw+tHV1UPx2Q
/ykMLyV1TJozFMIkzmOh6B6PF3FBwC1wQIHjV29UlD+QxGrKx8fF4h5BUkpiute9efF6aDZ2qU3K
2o1wQVb6uQSKcP0DiAiiFgBxqpucBWDHOEYvCS4vl51YqbiVZbD9oLiHAnc4DvENSyzs7T/ji35n
4X/NXvEA2d1Zwr5FBOo03VEi6AtB2+0yVkvrfr9o4wmWrUQOX9jQneCqiWVuQKhOYMh+u0V9bEEe
7AYCs5q8gL/V8P8OsTqtssQwiM5b6xob9xgKJ+Ke8trQhYrzIFqHzFRWgxwvOjDIPeZVfrFN4EZi
v0usKmvafR73EEM2xRoz6zNVmjzItjmAcle96WaBonpk26xziUY9juE4oT3zU2h7oo3pZZVvPPIv
YQ599pQHlbqc4ish+8Ww3PCA9ClIxTQmSb7Hal4j5yGKoMfA0W2PvieRsnpRtqT+HOL6a1KRwVHA
WjCr5M+z6dBZgHtz3nV0fWVVFSEYrnc6pWow9TlhdXb7wn/5/g20YpNAv2ELa81OoTmX+2PQFtG8
6Bqa/RPzYDWE9nOynteYoC2M5EOwYEOwBhA5N5xFLtaig8RAOXRbZ/JA2fhbwWLXvSUjEqGGDZy2
QDn9c0vePvMlYr0TWLoRxIQer7J/BixYnYLydZvqWlfpzWfGPfE6ZlvqQKqzFKOXlqcA4ewQkWEg
WH3WSad8pvZowlbFA6gg7L8PiNrSNFXyi78wYI8G/UkLSHqw5WVsBtlTDx+0Wxx40wxsLwpTpMbH
FIiAQnsLjE/F4Y9BKl8Ck5RniR/jttjxVHHV7j8zEqpdR1SS2IOSpaVCLXyabVuI1c9JmDIxxCss
8gksTHz0vom8CIwDrt/LhxgrtWFY6fJ/ebEfJuCVwtTAwQL2mspm9TSJq/qXXKhYW6sjv/1k0T8E
cGgHTNeTYFC2bmwyyQZgko5ofcMUeGJ1kllzmQasDNlaOvy6MZzp8Oh+IF3I9/ylyFd6Pd8bT6NY
d28nibopkyOiFNjnJq8owgc7Jznsswz/20sbZ+UL4t16QqIxAlMz9irrTD2hSeXobnlOlXe0HV9s
HjjC6UmfG0WcO2a2S63LhUacwFDj+r9x2bBx6lU/4r/Kfp6iSgBdsb/ZXGD5m9qpayZT+ooQWfOj
oAqKNhJFfZR9gRaXKosoRHBOLcb7QYdcBqwV0BOvXozvhf8fVuFPLFl3sRw1Jkd16Jt3XhDH7hAG
fvobWJdbbApEahSR0jxXIzrxZOZz42lQc6Y0KZW30dM81tlDiz6dSoi797mjXZpui7RwZjVLBv8V
zqIp+NCe3NpOtnUQBPwFuiYOOFCQ4480+6frcKIaB62OYImQhf3TpfXplrs2tzXF9EAQ8cdCnq2l
g4IdQe2P0oDG6GnlNaxCbI0J8KhFi9niiOaPA95uDGOi6ORmEI3Zsm6DCi21WaADp9eJp/3GUJvX
H8j3tuorY0UAv5jqzAXNiQLDzZAAnICdwanznRH3oHFvyUbYDhYeVnkPVZft12Wx5XQSI3oOJLoB
oJbmQsWAfR+Z1zxmAp6AcxbxSKG5FBaHI9V3z2ohCcC5CLJNnU9nH5tWyxkFgi4yMnY4JkVcfmt9
P2+/Qnzcw3ZCgPF7ZycqQq9InRHXyix3qPpevgteXUNWwrWlyroSrYehFsk3+SaNjutnyO5pKs8G
kfTKPHXjnFirHvroy6UQG+1jBf0td6ytkT8Xo7+Vi+UaJzdKHsxCcrTxamUcexYvCeQZ7llEVkWC
+bs6M3/YyHhSWq/wdaDF+p7T8D81CJ4mKEs9LpNF1cs+N/QL2bMKqyYGB1WHqxIXifiwDaqibO+s
OkVocEdYW0u9aKGtHCCAR1fq9+3Fa1Uqg0SI3UeV7aRLdrtMl5giOUpNj5/xahr2Q3SMBg/hTT1m
Zc70EPqY7gecgkt892H2jQAhlBe+8wpjCqPLHXsw5Qovg08RTaVVnC4d4dR4srP1b26Ho8tbF9Ix
2ctdBFMASUp4sMljjul51waCYJDL7dD9lEwgDAmrYMfI58aDvWgfHMNxw1IM9uMYUZxrpWIPkxEv
JYOsyW2bq+WSP8nQ9g70ie12DZt4ZpNocwxzc9D6Gw3ps84b1Fd4i7LpiIO0lZJzTb6qq4ZUUEhV
481eSibeTpARTP3myLt9Q11Gj5Z9oewlRWf4kZAjedg1gXlBexzGCXLE5RicN52qMHqz5654Mawc
AhZYI3EmNZOV64rBdQ0aiXPTuZfSpsEFShHHM2bOZ8eVpBQaVfc9ATCLuNkdwuoSDwl/w4FgBKne
htQpxk79H8jOTKQgcL0teXRaWAU2Dq8HjZ2SuJMxfo3GH+eWW9XhjF50UuhaXeUGr6sSeJKJ1dZF
mZhff0JL67xNeYTy+48Z/WxVAracxHZ6yMa6u9oz6q1ZaRdH+04or/gzZ3jO+xJLBPzXTT3FTYk1
YRmKwZqemKV9fB9NYWP6d33Xu1syVY4uOTnSAPci6lvUUElHpD04OuVui5BBOOM873+R3Ltgw/eb
2Ha5BlYFviDfc7Xje5KgUkbCNawld9CS585KjEqjKKNg3JlXuUl5NKKnemoHV8UPhccotbjkQOtR
voHduyyTEbJihc3m4mmHuIES4U41PAcr1fS78s07diUQKcx+B0ReGMbqvnk08KTss+c8VME0ZFwC
tRsAwvjoSfTpG2UYG+DZOC3bX9ukL6Dq9kxil4IHDmj2/tNvz54tZhFPgphvR9XiwpIYewgKs0zn
Ov26O6A8m4H0K9LQC5qkfK0tuLH+vHtKYyqY949bbldI6TeZP0Z+OLOH1aKMp4m9HkD9xKeXnKmn
NwspRCp2lCVVDEPSQlWwohAl1sWwpQjc00Uxi2afPKjUvhMgwoEe7DCRHBtKf1anMT+A/JdIrHR3
CWuQBtPxcvW9UH9ileQdK0rPPJklOhF1kaS3EqHeMRCWZ4n7eh0i6IF7ocly54/90WYkzWg0jvzn
mrVHftLVR2+ssy6/02gbO63IafcQTuhxJ8I3WvBfEFUBp3ccimZitwdGX0AYuYvxuiUC+hUqr3+Q
Z5mtuu5fmBuIWL6pDMax7G9UyZmG4netTl4bUcH03h6muUk71sl+W1OvpB+5bhmwS8KmCOWQ7Dh0
XcFHW6qtbcro8azL5xdHGDUrd0TS2BUs00kOoik94gKR/xbiH+M+XGpuiMb/SIrL7Y0XUWcXZKa2
4vRRocIjW89Sdvtwp8IspWnFcSUzXdz3OCbfioTckeRq4pY4ZmjYfi0kbbO6ei/DKFw/IktI2VOQ
QNA/pZKf8Djtopy881krsczd0y0DPotpM8rcecgtRT8STmhr7ADR7k7YFctFLsQG/H/19KeF6e+j
jJuzle6V6Qs+T8ubnI9f/pMcBKYySlAjrDjM3V6R/7hjAnpR5200TcwDKMCvMV19/V7XkJum2Mn/
ryHNcqvMlVEA1bJuhqFghhtFTXzotYVZH7bVLkeUUFNp6DfMSBeAFqC9aDMgE7dDjOT5LoET3CKm
wBH1w9QRLBkaKQDc0lIG/GNqlBOcjZhmJZECa8O/5PgMOHAm9iMoMOgHAkAc+FssuNZO3lS8JdNs
qx/dfVgqqJeMsX8jS5rsMLT/S0/ZhWyG8MVgxmog9xt9pLIuqyBGtCJGoBWus5HuNINbexsjO7+t
lbFgPTCAN09rU0ytNEZbZR+mptKcev0sn6UULL/7S4jy7jM1SU0GiS5SBtvYWUPJ2Y8YZo9e/34Y
MbpXHjXnP4clXqYhy2mCOQcCCB+EkE7Gc8yUuNrz5BydQsRn9/epunWeBVXaU9DzJQGV7ngE3ZnA
J93wrxMJP2T7wH5WzLI1SQzBMcl35ihL/TF+rAeuiEPINxQ3zkNRyVcoxklrF2CMHU5Zt+XAVfyR
iN5MzB2wF16Ifk4PdXVqgr7FKHbfITTmhSRyhjJYSzKa2P0TZrEP8TpW8+F2alYwaeBaOGNzO/sB
MdAXWbLak2W/bp08vwzmX+vuAEOVuX0f+wgg9rhh+lJ4KndBAhruT1lQFRartTkpU5B9SZA7blZi
o9DSjdRWk2IH5jC6WVrm3fbv7oG6xckkZQqWZcQN47Qh5lXLaQSU4wLQWbClC21GKSGAeOfxdkT4
xBqteFGb3+6j/n/ZmQIfGkLNP32iPAjE+/on+uNP0s/1muHuuOwemYCeHZX0L13jmQ7omxnsHE2P
kBoGwAEvZYVrBEIUhD6rWW0ncHXQl8G1fm+kKTFPXENbT9XsODgD8v1BWSje9pglkIQ22eNmkJGu
1pmzSZ2mMZimj/bp9V4EImbYLhDY6HTV84O+4XxuKTXUikjF/BbGwoED/2CZ/nhDjs+HxWT1CXMa
gWPMMoJwUhRgn0GYh03r6uVh8/EyDgaXWRQ/cxsJ6lF7ZIKJUfYueuufd6K0oBedbEspYets5ioj
nE/G6ulHCce3Nidp9ZpxRfczUe3C32daKRHRCi2UP51sfN5lrHp+O0ocqdgjx9Wz3vW5kCKoHgcg
bIVdO+fN+eiHf72BygMfBnLP0G25tC2b8nIiZ8vQxd9EImaA1CyR8HKlVFnx0fa1nRnR8KJ//Vom
drmmKpvScyyP+bZvNzHTaqjvzPVh1lYX+zGTaBujkeA/gTN2T0fWFz/tYJ/Uc8/ScSBMFbkU/nBY
bbC5MF6r6WkbPk+1hFwPf7v3cey2bTD3NETB/+/wHyk0FNau6vVysjpuwgYAvzIuSa9a7VmcRH+i
HuFFXMpEW8DmYiaBRKZTJBdKHHEVWhDVccglh6qH30xKAun3VwupMJa84LosR/dYqKtjfl79Ig3M
Xs34OGVmtV33kY8p0yMeeEDafx4JiGTwEIb+4JN0xte3+24cgJntPbOzFwRkcg67QahP862L1jV1
01ZxLRBbexu7NPRd+ZFOOlKvXSLDMbqWX+s5UPFpssvGqdyV1l8oRmnKmcQxUhXJwWzblFDkE5Lp
EhWsSTEb8HNOpjK2n52+9K6XeyTz79W3s+wtIuZhZbqP0Z0YVNLV2gQtkAKZhzWz8vB2r/hQyztj
v3iGF3ckuvOOVAANWCLfRobTfakQmhcJegYKvrNGYKmXx0Rc/fzESf05mAT6/fc5Hc0j5idRNnxD
Ed8XDGfRS9h9l84BS6khpsO+2w0F4oIvUG+vaKY5/B0ccUdQvaYm8AB+hv7CdzuENJjNNFRjzKHT
hyjnTOhdAW3gKfk70JrXLKESKqwNpH5BYtfnUi/tcBCL3/CkgvhxEMmWmqDFLLLHTJ/LeU0k01GG
V6sHolonLeSE7lQ8yS6ics4eXa7a7DStaoqF87XHWD93jq12OJUt0Zu+t2TwKeKC4nBlrMERNqWt
Q5jHc6hJ5LWsIP+fsn77H6TelIjFGGV2HXsImmOeNMB1qzo0/7yIQChy0g3DItVQfvISAQR0VRQ9
YwnV9bkb238EtevXP+okiJdHUCc50d4fxK7IFZJWtpY5kRX7UaeK9wZy/GWy9Ih3Nikms6R/kUqY
pMFd5iFotLg3BjNG0SOHja5RumIdG1Jtx18mqJNQ4S00CBKFNm+Rf32YMSVeNOaynO/fT+MjVD5S
15Lbp6xPLOHv/wC44mKMVRtyPvb88C0he+dkckh/z2ogSWRNz3NBrBkFKjMoTTLGygx+BlRcHwvx
rAswzQB4Dxd2vYQ5ZOIC3a4QbmfheyRaS/a+Y4mYwhnl+lGhWnVlBhXZ06rrxoF1PZgGxqb2OUb4
SmO7h9O8M4mC3IrsG9DnFDLC7S0TKkyeyvJsiOwuS8V0l9lh/n1ZAqowEmXXuTi1QRdg85b0nRZn
SLRUyKjlHSeD0nU4AbkBOa/vx7erz5HYTOdh/H9YhGlt6mxsyNs+HNqzqkkY+r6yXlnAaNSFYfKH
afo+P4l1Hed4LuHrBWzWk4BmzPeNKz/iPEJZ7PNAWn/fRQJ0tZO4ZsrI7/lWrrzhLcVJA67Ea4zD
NSaF980VcOix9kohfzfIEm/bHOEUUXlUOKvd5gk/OpRVdv/EcL22oArVuIKNQSdebz3t2cyo0lWQ
WNugwl4NbH4aV4euksU9AHKOvjoz3Fb1SYTgVBAlBjI5Ntlcapaf4Xyjmtq0MZCh9baQA3p9LpsA
a7c8FMIMRv/s/gb/fqh6hEQ7ahAwgxXFP8uG2Nb3/dEJMXEeZiY7gQNtJOAwaItFqd2UOyFsSuA8
cImDMkF06hhgs0NmRXV/8PBM2Qw9lVmNf9YS1mt/6LfA+y0IQ+xkyv6OnVj49kn5djYLDgM2odho
X7j6yjE8E7P7FoDvpalQC87uurHrKg1ULFh5JUm9Ize+wi1CLcQuj5ss3CRcMmViiTpvdlFytpdI
X4ukoqXsqpQZS/K/DIB4l2X1WgtZAbm94zznNEWDm1iOILEbA4EycYlH0GUGbNV8dpaH8A+Z7gZE
3BPY0NJPNYUr9MKOiLMQk4TDRwflR2mxD11xLYb7Q0hqCyUi832ZqEmD5II8Bx3P6XU2zTVwxIzT
WZnkJOzat6Er0gw+KJDQCBvjKkTieMc9QbFRErG/8z8GvFGnWt7a1wWbd0oawSTW6n6lk2K8aqve
HMAR16G2ixlWEIwq/3NNgvBO+K4hZg+2RJR2JHmAbeBcIEjj82jtHboiq+wZHuMxDBLZZOauFB4e
L/3hOQKQdszm+kakbzG0X3zJphUTwBxwSAxZ108gtedgfMetPvJ72ldXo2FoR6Ebbavj5TUqeXR9
0PznEg0eF3l9pkTVg4dfNb6234dEALKDXgl0XGZjN1ckTKzE7BTXv9D9t/W9WUNG2whDu71vTrpt
Va2fRrvJbDPu3jHx8QQ+GFzXEsM7bicAfX5x6npRiD6hrgfWIWNbWv6lGiDMhz0Hp7Fmu6OsUxcx
gioPSMoWvyNk0SiLMdfMzrebagLUVr0g8Mxk+ydAvRJ1ecAn6kmCHwD1CEBW1n0S2OHLdCjilR1t
GmYUAdbNjzCKT9Fe0LQvesZPfx5zJjZARlDcsBKXw9pXVVZ9VJNTyvvFWEuCsMkbOOy3Y+pYrUe4
uIEHDSn2A1hqqrtwdvqVtX32IQQrnAZt2dlNvx0K6JmdVhbOTGfl4l0c2IHA5fp5WYasPU7DR9is
h3vOA7cWaj/udLdM34ZPBvYkT9kEa6PjysDmOQHLHG5Syqfv5o4QsIxQvd/0U1uFPiUzFiE4na+r
IaGHr1HxBuqY/Ez2loDS/2b3wKIQ4CXVn46r7FCeFAEP+HjlKWFBAy7Fb6Q3Qz0o12fExJW3GE23
o/cQ7XULA5qkB0e4Kxry71IdLRrwMGgPS7LTClWm2fHCQunnE+DYkUF31T5Hvm2XIa6WgO07ivxL
UmuKeLq9LyDKhuSA2WyQKakOjnfYxesjVkcuBwxlGLjXuLHDOd83C1q6lo7IVSzvY+Ko3mk7OGR3
auf30YBFV46pSVABPLSmbcqHq3lJC1cU4YOeS/5xeowPEpp0aIuVCyW6+DBFpi1T70YmWG8g3Cvo
zlrL7EgcWx/VHWHeB6SGjc5Y1VXRArwkMjo/Zs8dWQwag9qCVfAIZ3y9O6v44v70t8hLQtp8Vk4o
HBWADk7OJkLPJOf8Kf9s4IsBIJAk3TYb7wqElUdN3wRl9I0Vk1uSlz/qQJrjZIVFlSI2T64lsKt5
iNDTBg8xzl+xQb/wYXWP15iGJSHRSiOceVu8JG7d9LIv3VPeK+bmorOAPywVpUltqXCyHqqr4Prk
q0wd7pzqcep+hMt1JKt8tyrC4FSrtPPYNqsBgbxI120W8AfNkTFoU8ThmhsOdhCLD6Cl+w6N0kO7
zfZT508oukslE8PMYmpm+uTuUVaEjdJbTQS4RYPH9HTEMv6yLpbnlQkStj9B0LAb7cB2mrdC20td
pNZH+3nAZGZZZN7qRdyn4n+nNDme1uLHWYyiN00T4cw3VMZtSkMOfK6zVn967p7XAWDqbZBXO3vX
3dECRKTXKBFX8VDKOYK+dFyxicyhyGea06x6uLiKMRmAOFRx5J2+VMGB5k7NPFf8OXJBc24eEDL9
3Qm+Wkp4UvPogKPctkfR1ULrQPTY0My4/wBhHNrIKhiEpJi0K+fkVSiPynUSoszIIepWVqkBso0u
1hoLArJXl8jxakM+Iqoh/MtgyySW6A0RUVrZyPazdnvmQL17vDxO1jBUrMzLHrIE31UeDyG3qj93
adqDftQbuDqRQhVYplmAn+ywV+OKMKepyBWCSTu7PCAGthuDQw2lo0FL16LwDWzdkYIwwNHc7tpl
fasE7naTx3WtWAz5FPUaZwlwxid5a2g3CThQsDopY5sC1GFPuHqPggiiVq31ET6krQXdWqHG49MT
Xkj0W1K92rTX6Fc4h68NY6InVv4SpJFExDf3aZjlbp42+dexgsxo3i+zOzhyBt6dc/49PDd12GwF
C72RSLCPLkUQuakIDPMWK2y8PhciPWQQOV1xvaX6puu7g1xzOvUhraajLz9jzqk9Ss8ypweEOOdp
wQ8LXKms988keimY1FqHADoGbv3M8RnaG2B2yUi2vhKFuoatl6ZJ7SDRq1m+uJmCJxwY9e5zGgsr
EmyboyvKWDY+9+gRGX61ME1+Izh1QU8XG6xUx9nqIm8Z+jPs8mNtNUTzGOXq3dkAr3+kYn96mgpY
PfmYxtynLpYvrjBNNybhbzq02xUvrlnODhPEzSyMJQ3zh4+TDW2zLCWRI9FneKaO01mJNSFS2kpM
R2a+b+4rgiscycNE1sujKSvrz0mWj+Im+dRMi6EiAv1KViObDnY59e5Uc3zFJ1csrJJl1DPMkVml
/r+XQ8Nc0BKlKewnaDGR0BeKRu55tFh15sRNuW4Z2PsC9XkkNAmctR2KpmT9kJI877iX0pHGoM8z
YwgjSwCXfSAr7uaiG2dWxg5LN//BQLCpMMNS2y1cQlKXqgI2+26vT62NKlgTkSFlasTeEG7Cvsnx
yXgOW4ANdln9qoPbJnAMB0s/PEv5yd5+fuhEVljeotgCisnQON6oAV1VjUwzjRV0ooVncNqLwcEp
8xrFGlSCs6AGFily0X/rO416dcxEpd3Alu/X04A485CCekIBS73OlwMyZgGjGjtu6TGcpuwGW1px
cYGkEoifPV5DtfMUj+RY49TKOyTSTQ7AfAK2grVHLtBhvpDLxxtylaXI24YfIeHQsK1cqL2zG434
OBhWY4st6TrUCdXp5frei+3LX0UDCRrJKczazCfWnPVvr7Gu22zvzoSRMzHcBZQk1kRF4ZaDFey1
e6107DFQm2PQbdKS4T7BNUAj/Ngt9IsfRb5GyFfwtqMbLi05B46bgpuUHoSLjPHUpICF3q6hSQzr
c6GuVCoCGt0KmNpuUvnv4RlrAfkZo14Ki1I19uSa+3F1tXxMDEXeO8Y50mOzCiNIuyCw0f6FqNJZ
rw/yPUDw2jsJ3IrBsDhKpJtoxCn0iB0UXYxOT8KHV7xPaBs75TBKsj7rWNEK3NJOyx6sbe/5Bwjz
Zjj0T0Lza508iKPHTocjV7cisYWWEpeLErdLOkRRdbjczQC/dmMlgYRCSApyjP7YS7OCld2mwZ/O
SiZL4XrgXasby6MULUO49eITnHXbePW+bza7eNZuObJ0EGHmQA9asZGQtnYVU4ZNGDFI89tZGtuc
9jXQooimlm07jjj6mAeZiQOge1vtsro4C239dIPiU0CXEE4B3iX91IN8OdoSk7kRjMLJZK5eGMGI
DQ/fhsLZT+8NpBnamSkv167CO9zUwOJ9cvtmpnmpLMUDvmP6UyAiYn1DefOfldLvwDVJkY1nwqnF
3Cw3tDDMg+Nd3Z7aorgo77/dl1szHX/xRr+A7057x3ONEYwwF9lzclpeTyIGvyOBVv7UOHF+Kq5q
M5H94rMjWRCw2lDDx2r0bkcYAsl9Gub5yaBBmNZr7yFFcHi9VYvnZ1WwtsQyQoxWovkjSTlnOP/Q
j+d+Lo5FtkXD2MHRIogJTyZK8gWy7frntF9RXZSDZso2zJUprHF0mdUHD7zbbr6wxlDQooXhqPV4
sk+Q8ZW052fvcLVWPP5bOP4ybhW/vFJB8fOkUVExNRFlCjCLFkdsNP2MJpO/I5xSsGjrULaiKHMv
5SCmIdJDqOg8kgVPAeJhR99x7gTZVEWp0oWhkHo289Sb8V5f8kExglYsjDTHsyCUlWcQKl00L9Y3
csu1uHHue5jCUUZI2DTBvd+HXcF2Z5ZUh6/gAbJLYyadrgE66/hFQqn4PTKtmRIkY9ACu4r13nXN
m6GTeWZPM0uRnLcpQotGvYNmG0wzZrmXv7nnF/PIfTHe0MA1lLlJ1lT6sOZCQ3AYzu1UvmvTMJd+
mqmgqYrgidIQVgiW6UAuIFx4XHkMfiliE5KguRjxR0B/84z1ESEOuA+13j3mBkBXp8HKCfjKEAjc
4pAaf2f/qWRY4FiQjiuOiHOTrmSXWD+4o2IKLohrZ+WdcTtJR94Jfac5oUUL7x+Ej6AaKqmVfwE1
BWbsvPbNgq5whrgx6N4eZ7ODUWPe3K2G5Ox1GRFUGuF/ViYjW3F4DbkS0qwD5qPkz03kVFcUFmEF
tJ9fjYmY4Cc5vQyuCV/5VYGgXi98xoP6cFZve8WDO44eK4Zr19jy3O2shATfI4HIOiITFCMkbAdh
zJEuBQcKSzQwaouWbbMMdTBVf2cGPeOy25xki7dc73UFG8A0r0o8ocv9IgMdXVN2i1thSKyDXkJY
m7sEUhMg0OwB3SntatLvwR2BiioAcYe0Z243VIC+wbrNZILCingVuWTl/2RVBUXOTKN7fAuO+b71
OZ14//euUbUOSfFeNyQr+x6Xuo3Ur39jo/9gi4VC8jqAR6Pz6JRkY2tgkXVXF/u5pHmoMLOJtKMh
zetzM/U/WL0GqG9KLkmgutVpFJ/HY9erL1LjEHMMcTW3fImdIjut6H2WrN3xOUGVnyv+Q/u9P4FQ
1lWkRM+FfzAEHrLkhU5EVbt1UvQb+r/IoMjTT7tOyGQrjTqPpbR+xjP10foWyROP2+kzikIowVQG
lzY1NCXPyWIpPvqEE6pVGtIkdJdyfN4W6WHKu0q81BnrEXH95an78VesFdbvWvKVLIOAwg6R2k3e
P+OivJXv8u7z5GWk2Skvpz2PKYgpd+6ClJVNMPSC+aCXvZI4w5LVQXVf3CZKMHj1cbHNMc0HeFqM
Izp68ROBDwk1EjwsOQDaqqfXRogw61IijTTQ2ls6glfrsC9lTR4wb8z4bDSy7+Fs3HA7gYV3RaDk
VtObSKAkxR3iDpH3BHzgKo3E4GBje5YCpL/r0Q1G+lqJ6sxTTRr6sTd3leFYT/B8T/cqz9JFn9oT
MSCmfY6yQe3/0PERUa5Dk2EaEZFWoQG+8w1nLb5/+7McSb4q5U26D5G3O/rfFFiEVHJRd5FgjiIm
3CHBUrhAx7MlGp2W++HxicoXSp2rEpSvGIQJV0Lb7qYOBNeQFAW+v1Z8G51cjHjb6IEds1bRWe9G
iLLhIjhDG22fgv+hSSFOstuSnqvwl9NuHzqhkEICl6jd9brBW+GV/B+d3n37pujEp8BkX0cHRAK3
NZlZtC2lUKDxMnyMnOT82MZ8mcg2tsw3KLSjmfkE5fvUURTPAtaA0MIhQ4gBZBWi3NFFVoirPTbr
EjR2kT4VVaL31vp9HMqEU+bFjqUbN5P3lKlh3MKwiN1SzWIXlp0MVB+bbDcmCXKEgajbM1m9246Q
f7vmNUEW/p2V4CCVDI5KZcZG6mCUPINwq95Bcmq+2r/mH3XDePBxESikKXUmdTQxz3ZGxuUo/TF2
NwpIzDEtAfWPdHHjx3zmR+LtJ6vuF2fFXqLgQDa7amibe6RiOVDC9b2Z8PL1lUZGGLocHNlXdzGR
AZuvqDgyGiszBdOR/1NhiPUKLuaK/e6ISJSw8BmLe0+sNOv+PlcTynZx5DJWcFI2amqt9RuqnjF9
sxFYII3igWvCrz7iqAXVC9K0kqZToVN1NXJUekA3AWb2YLkIh+u6h5IuKRc61KOZn9DDefj9J4xc
/GwuCtHCq2BpCYmLT7lbpHXFaIt3B//deWB+1mr38bgL4Hr1wJbFIqMG2O8zFQcOmc46sHn+r5uJ
V9iYLcl3KDmDtc78SSH6xZQ2FuaSh9NtniRrGW3kDrDEbEHuH285A227PdiwjYJ00BlRffQ6E1no
xJFXczW3WxizpTDd5Eo51+TpZvLzTtyYMSl6sOg/b3yUBcotj9cVHxEGroja22+TKa17cFcqJsI9
2L/EC23mKnlDr4BdiWNLD3qFxM+/XthHasF5c2HJQQDvZG5ASg34RhChrh75j3Vq/++hGPGqNd2r
9Ttw8rx8gNqtFKe3VCFb27rN3wxy/HM/cRR7X9GCcWWG7wnCpiNckrafFmuW9cb0/rxFtAtQN1tD
pA4T+zRoRcpv/ham14+gH7xbQAEHmqLXWgTtU6MAW0XPgXfVhk3pkIeY3zhIvilx6QnzodtrfQnc
5RBzN5jpJKMQbqb2AYlTw/fKL2lc2XIUHAKDVCvsJ7y6y5+m7hnU7fffie6m1TPJXW2+KopGclma
0dcKDI8JkVG6lebmTnfLptxzrGWRwmsxbrdRu2NJc4pGv5SUD4C2rsoSRGIY1DhlN4CVMz4qAv+Q
DKxfQBbRr95MJbp82XXrz+41LkVBKH7U76zg85zcwyrLUUawS/Ur/IC+lVNSd13kBp92lBbUaa7m
B1Gv6BzO5prYHVS2oxA7j9JjeRtWwXB+akwN+Xot2BfbqbjS+A6u6YKE33DzHPlWlhINkP6c+0RM
XYoJvOePDnRkrUL2KDO5O+5PmfP+eiaharhYeDOIvXz1fDqg9Faq9U9beIFn+ahF6xfN+1IagaJV
O0eUloUMX0iiK0JhpmCYmNi+SNAhHxiGfQ7u9D+wErPMd6o+0lOWhD+x9R7C9NIGQtvyuk5C0sUm
+lK5itLUSLfkrxub0VNkGYnrxXsaVXKrilGr4wC/8YRKu+KFqO/Yn7pIqoF8Pp+zcN+5M+Tsf/9F
S8YKAD09/XgKnpINpuisu7wNaykqSg0JkTPReY2V7yReQouRf8pe5y9iuPlKtJqx60VLKfWV1xOs
pkmgEzLI8f7d8TlhwisNLYQxFd08daB3qgqIj/BB60ysToWo2S17Z969Umr52TZIQrVW3q6gdPLa
DrMpqwmqxE9WNGeT1aMgNvJrKw84yvwGXyL2/TL5MFWXJ8z8bwrx+KulQXBW9OyAhHY9N3B7aBq3
v5ODUJqTML7RpUc3vh/gK/AoZyCRhS0dd2nap04psux68e3gI/YlO2A6SWMZOtnL8GezEPHB20tv
5BhACnzUzrOLL9WUHUIVROMENHCVmRz3CHy/Aku2ouB4ivsM5a1w9i0cszNTd/0+cn4GNx/L1nyt
LEFhfrdaCdMQUfdAG9QcJoCXOI2mOTk7S7F85jN/BI0AoWrwpclmhIxlgAGaaqjh69CavL0XpdD5
BtKVpAFri/wH338YAp4Tafvgcxk8F9+1fuY70SOvkMTkJ39OLXoCSrQprvgQ6wUd9GbxK7no8Z12
inQ1eLKitS75Az0oVhKsyn+6huBFYOeucUKe+kvqXD4ctCk000IMOdzTeEXOQG3bmiTBZ/9Lv0hm
pd+Luoj8SkeRCRw0mdhhaB4G34H78s/qFrrj9PPwza+P6ZWHj8r7tEgwNKOog85G1+deXQ+TP4om
iY9efFYxDMJl4xSABJ1/ZgHRxky39EtsJJTiBPN/BGJ/uNRnfcZLLSFXmGUJCO0K06jAnquL9C84
pZ+9qq3MTW9eLZ5NmQ4ys6rz2vJUzUbf/wpF6aS1bAWBWVVhaz4P3O2qQ4J+KZOUDp+qNUdj194j
fSOYuxVLHmYtXx8kjv+fbHqPwBl/nu80vOK6XI9D2QbsjZp3G3M7/yp2FpmodIaYudVrktOAXm7A
ppcLmC4nJ4iEQbxxYlA8SU78azBPpKu9XdjScb/OYbi7I2DPDUkFI9d0CnrRsDWABtlPM2hgXbNN
gsNgJYy9ix6v3qflGEZUOZ9vDIxpAJ9bFyRMAHzbMAEzeuMCmf9420MrlfhwLFRqKF7TAPXFUJjf
um+DndzdXL63tmIKnNDSr1SMmXDed/Uygheqva1XtT52lHzmhM2hoVX/ZSvdUlndOfEi7HMNPhag
vkhA4a6FuEhVnTtcrfBbB9B4C0hi5uIA7hzw7dekgHT5oyZqRnuA4msr5XRqiXNbPy6AVG8XQYg4
Cq3L4wxtC0Mli+xNNHNm+vjecjLAKoM0880bT3nuOLPJ+beR4w2VhhcwBmFczsArln9EiCGgC/Db
91s3RMeKGBu3+mR3CPC2TxVKobLySTLuFLDDg+6KL2CTJTBGKN/9wla1DppMTHx4wEjj43B5C+xh
hrIjAzfpkZk+PL2Iuye4yC8DUYmfzACBpie85PQU64HCewlo+EKg/OGtEx7I6cCWVRWKkm8B3YBL
X1woDup0PadEP1LvggAtNLwQoUyITdCiDjM/x67qFkyoHatwDrk5F12YnYDeSaTYSqbRp6MSdj/D
BR44GYkBLWfPn4wXjbJMJ3z4sMu1jqqZn7ELtdwZLBw7KquD0lKN8yoLJMIeRxUB8YykxmN48fQ5
9vI7SgqSarA8ZUeIBHFUTIjjX0ewMmUWVfVaaYDJ56/SL2OgRwFv0d9tb5E/U4aGZO33s2pS+ZOH
gT4VIRmlA4xQKizkZXSm9iheLLrZ/fykQie2tXk3JjgGY4glpnd4nP1VhgH6qVuhIyfrRjxvlJOb
cpDFvVEwLLGeofW1ETByQ8Gjy6swfbs/VrsJqpy5/f2huHngAUHEIY0lb0PrzKvioJwqT8CjV0Pc
Yox1lJLH+NihuBExh/WhkAEyQYJLviFmsJGBwbwxTmS7uDAG9q8/B97NzVwcknLPEck9kd4rlADl
n3lPKzVd36TtgFgrKXD4RCT878YQ55/IkzYOsjxRBjGOKYpmefCKDl50hzBUs6nbWOT5l7x7qhUJ
CZS0eJq0v5gOklpU9mhtGrdNNjSkTB1D/6yKsxu6fL/iO0vMY9c/Q/5qG1JixdXoAOa8C00cRwxJ
0kxU9KzuKj39aQySwp2XeHCeLMT6rK4++lJhwjpaIbn47WhSdyorWASTq+zn9rc7nFpHx3laypI9
DWfq8XVIuJ8P36bohvyej1GMQSNX/o0hHQ/sL908p0tYHqsaOdCD2uJo7ZrGbWLhFm1S60ah7f1J
cFTatASgeov3gjraCMABtjAqkefcsoIti4MjVZsURC4hPbUhn35MUttSFgEmf8RfRLSt/UX8FYvl
c/QRSzglQK9l74nBHrrpLNH1UWSm61cgYVMkALpSfHcNCBrhTXSaakE5cc+zPtvuTb/MkIZCKsKn
xqE++AbdZTFCEIuKcX1MYq0fZeJmmrHafvMjkT1glI3Xf2wUFdp6gUrYGCB8IB8DSm5wn118h4Pv
XaaI+4U6ByF6WibEOcIjcFW2IJDfr1ybFv7UEuainGU3uuyEhwRQlIBEzF8xnGZLNNK3U15y/KtF
z8Rj1T5IutQT3ejU2V8wi+MSfnEt/NrcQbOzySPZXxfJd2tW0xLztO5BVX3mqEXLpGPgcwhQQT9Y
lpcfutwUXFPvBBMMfrOk1X8gPcjdsXy4WEol5LfpYXLY55GYFvIy3muInC9mrz1Pm530RrD3bAYZ
pda7lSA3Clq8wTN3bW5ke/BXyEUnP2qVDZ+F+Ictnoex3J6WnmK8um+Wha6ZTxapaAdY35g3aIJG
kGJ70TqjQFwRgngOBjQgcn267XMc4Sa4rh48eaX054H/ODc/+wBpjeYyfvUfZLk5NU3b2pmxoGUX
Q16rQBD0T52kj94cx02dT9cHwZ/IMMAY82EnClgxxa8cJsn3xzJXW73VbCerR4dCGDRwJV6/BWm7
Aa8o2buKQ+iMColpr152u8GNyySW44pd1GIx6n7bRiCczvO3iYX10HxTCW/xfozil/mF3BoYUISW
xgdZ5UziEur4GFAg9vkF/5DrBwaxqaIMoUnZWuFYtwd0K+ICQv/w5GrWVFxW5tackHz1MexC3fee
I62B4SCgQWoWU9pUhGTs13PWreohFxzBqTaniSdQvVJlG+n2mWcFvzXT6t/fwTi58jGXncA3szVQ
UrVkhkNWQDpPKO+chvw1jy2StUrPRthhuSAH5MGktTikc6sGPgIGr4u8nbPQnYRAb1/UAmdWW6ZK
2YFUiovu9oIPXAgbVoR6vsPJqbkN/t9aIeHK01JzbLeVB+14nqOk7N/0VVNSRaSQCk5ftYsvsrCo
x3p9ucpvcoYjsXmztSfaONky1ujxoiDoYxL/eG32A2dFb4n08//kJQuz0PTaOJQMkTqw6bw8bioD
ZiqzfHLqPdoQgQ0jiI2XxeTSQRMitO99cYMZ2YYPWB5qzphQeOwHlr5ixqozIUcUeTvo0cliqr1O
bpuzl/SHZaXiHpEpfwhcALJR2qJ/P0/f6Vo+8mlhbTuwQC7CIL+42X574WRqJrEBZr9JOu+/CWpL
oxmSXfieMTtVjRr6Pqh18viXfQRxBixYNRLjSTD2Dd8H1V3/6UVIIU+q877O1U5ZXhJh5NpQkU+F
TmrMNJi7fnF+L/LDhj4y1AP9dLUSI9ITrtxPlw1nG6J0i06ULbMxnNso/d8SK9/2Qc4zW6bHgPTu
XUy43gGc7zX4FSPy4gfBcnKjfMccoyZDb/VDTvzEE/97oDlCVT6C7ybgeAd5bEg9Lfh3h8NqYe08
mCVgrVBtZSJVo/bQjwqc2IS22Z51gMWAMYZNQG3LLtwFfRcYTS+2YmF5Q2zbg7HykWw4rQiOITA3
ZgoJcVbfnT16VnpXubhRsZMuetfsXIUGcG/6abvPR4HoVGrTQ9zJulWWL3pZLdcbvM5JG/72YWYp
0K89rc5yutpaeSIJbYoINTzYMqA9g2r4OY1bujz3q92X8rhZNYAxCTrWhr1yEWtaHkmAc8L3Whn2
WimmZSfnCWxw+f1q8tVSaUsDuTU3+Z0U45eVs9hWcsZ2XajcUxnTABgCoBKUJNVFa+0HS4bxHl5g
I5CZ98T0s5JPLyPsCwPRZU+MbPGP2mRLJSjw2rF+Gdm43B1BZRULcKZozh/9PGjjSANvt+oOsHGx
UHMeByMfuVkIfeIux+C63uIPHUPL4ejyZJzjFVJ8Q4Yicn1wXZooozq/1fVylBBl23iW3TMJ/8OB
WsxlIUi3nWcP2KOM7pQ5yGf5PQmJ/7E+W+Kg7QsyolrQZqTop/qhvet+BUAw1YivE33LBQVMZVYh
U6UNOFZ9L1XwE9u7HlXTSJz2llgdBF4mKtdimMbrgYv8wfeNq6JpjPUe6coICVNUSfariuB+g+Am
0S2nqMIOnoO2pHFOYdiFWdQTno2qQ//DxXlHey05fWsXCEHDpBHU+Xab01frG3pN0Ud45+q9XpAv
nY6ZQ+o3x6QCrfGHRuj78A/O3yTINSHBMZf5E0RvWLWUIB90or9B80z8MKWvaQrFky/RKDm+Bg5v
CAyEkDUSQkK12GAfATl4zosx+FK2XHJftpIRV2f5lQeJE+qPiTIsFvAQgAjkk83Y1qy2DyTRR4ax
Nte0uy6IDz/VI2MgdZza1sVv66OUY5tkqY3x9Sv2GaM5TFj0sBblltxxElGcvSF/gsthuuraZgiS
8UofdQxQ7E++LUknPYYkMwZy/oxFpnv5nWZ6RPkqPnmZVohozPT2P0UC8im3RMS0fzwhqKlCDMM9
04pzcJZWyHT6hEyPXXIese8Ibg8H9UL7HDUWxNLP3fXBOYEfMZvxTttnARlyQ6zaBCkQFpqEvG8h
AUFtIx2Gl+acLh01RzFV3SIzXmNxZZjFpdAlAgZBKKIwtsd/Wtih36U91BjXZC4zxKaB/aHGFh2A
Izy8j1YBb/C3uYsM2uKgKJ29G3LnDrrtUaNms4ohXFNVVbIYNRSiu2J7hnPLfLO5+cZUuG5HNasK
2VIAN23MEBJLTA7uI9sNuE8kYJSfPTzXPCfrurlYmhNqhvYnSO7J3V0zEvhW7DiK7nMNxDFvK3M9
65+zmg46jR/RGSwIkHTcNbRWGHqN1ByH3+J2jump9RAEdm0FUD8ukdOTfxBocqqC2oHDS+3oiiWV
44Y1VgyUbBMjYKNroSBX9c0tKcvRiyfvYFlR0FNcAsb86MeV0Ka+zXpmPRouJZ6mwmUhDMCCJDbt
z4Ub61/TC440EOfi1tZ6qszVWHy9AzDEx7tOxLbjZHl364Yn7c9gyiD97noSl/L6hPbzDLIq6a9h
Iy0iu4VgJZwS57ybwuremuaE0aEfrJz23H5HbKzjzdTQdbGuT8KafBixjTsQ2MKzVBbVnGbz1Qrk
6lHO/3hXi79U5Gawu1h3Ik9BuPOfrPmExoPMAnFMm8sF8E49wMwpx/MBftJbZG49n0rlsHFWv8tC
7o1o88b+a0Dd2A0JYpIb5M8j2WLje3t0qZkBll8DakJ53AF4WKtjhn69IYMHgpFEZUBS2vmwyQiJ
+CqD/z7YR5CI9wAItkIdjdD9luBnbbLJ6dyNYtg4+TMlYp865Hoz/umRCkGja4Qu62I0BMxYzOmP
MOPDjUuAnxprsB53bg8YCtsTwEoWFpfaXJBvYyUrhcdLA6m6putA6J8hD1mF/wv3nSvNX65smQrr
NRuBFqKslVOi3Ec1J9Y7JSCHNVGUaOsC/u3oEO/3A87bVUA84jE7FcbQORqFJdk3EL90ySrp5XvP
d7Y35hp4QCa4CwrfBY/VFG+dYJXkU8xTw5lb1cmbJKBCR7kQjpBWsulmFAlnXq2vnI4r9ySFiF6L
Jpv/MLIEPSt177TdF3t7vcZIioNfBC4e9seVDJLNlc6WPM2I3V5luKecBemzshTDOrJ8tYPqCmRj
ZTC2f7GwWfWMBLUr0knRPsdHFOV7lrRpN9VyM65A8NG2vbevYg2EcaW3YWEwBGT5/itzqEtL2zAA
zsR3MZ5mXn74VfSrfo2nnQ1D9WbYMsyvKbojtluJ+YTFnWeVUpSc/MjKrCJ0J18664j/2UpRhPuy
SLyvUHDmBrkHQWSqujlDzDORag9U/N/O7QHl1UtLskfYxuNczE4W2O/ZRqHovJlyTQA1JmMtWEUT
VvKak2mHsoITV6gx3KDTr8RVg3O7PfPfmzsINWd+O/J2WbvM5cG/zwWkN1LH5EIfSPu2b1Q2Xq2G
wvlhriCaosZ4DCc5HjciRYYh4FMsINinotXxJuPQFCqeMePgORrncb3FmMuZqCNTt7AdSc9lCH/G
G2DsBoOHhZYVs1V25Ztok8HpF54o0NC+fs2R54a19WfrEcvZTkLfYEA/HfCmG7/giTJ8RX91ey31
y+JsriZ2LRQSFKDj5pFevAN/lNIrlqk3uibjUYCU3OOF+8OcN4TGpT4JMPQYkcg5h/2jkBEOb0iW
2s+1f6d5UQF7ziL2usJeQ2GIWudQHFN19UM75YXsrNjrAbh+5ecBsV5WA6Raa1WzOipbv4ri70+g
Nb+GOl/hV1jrGJOuWgtWcKg/olBpCJooAADuVy82LbACz4Ujj0SRSe5HSeZE+YsxJ01/RdYwbRaB
3EZ61Fyin9zHuECDmyRn45TmSPc6BAD5lhddM/8vPXs5wZ2+guA0qwOA6MlJRvPEoIvN3kKvMGCs
r31LXgS7RjcOCtdOhbEryx8unF9aKXqF4MlGtKrn01TDhouJZPB3lb9f2T/iOc70F2EggPEkqaON
03iPObO8ZGSoFfIZMsJUthGiBTmL7Q/87NC6HVCMmgvwg1MT0hrnsUVA73kOZ5t3DITv4puGPfmO
JnCi4qt8HPepWlksmkgZXxddbwBPK2wGmT9SrpNrcRzKcl2dke7qeqpNTtc0u2SvUQ9rHkHMHVP2
SOu+hCsAnEygwlDxOCYtMc3B8j1mEQ4n7YrV4NVIdVMV7ivRid0D1x1paVqsybIXW0peKEMk8v5K
IbSu8BDOxBjgp6Igx3Hp0qWmDA54L6FQjLVIzllcX5NPc0xTiEL8NuGYOA3GMcSHnmXIB1HWgEEk
r/tymzZucmSHhMGvfpJ8Z2EhtqJaZLlrkzq8pNEkHwP9VmdwAOqfAziZ34HkUY9jcVbNMWT68DF+
2hgu6gpjwrzhnOPI9UnrSUtOcDcowQ/ha9PuCONQOCSmafMIBbzXdYxh5z6Ieoi0PpYNDR5Kzi1+
aj4gGZWqEsKrXgbm4m1DoCg55H7wYHN0cfhh0UtywwH04OiiaekW4Qm8hNeloJgIDnuzTyj5oNjb
RGpBGC+4ssSJxnFgcsGcoKhWcCbMVKFxyDphHIMwFGCsbrfp7ofyazF0kwDN8eUYN9fthuRwLneK
HPxNFGK9DsnV4qyFxzYaRQYY8iW0BDyErd51XvqongZApFK4tyGUHhdCaPCJJ2AiCMhNE9jN4/ST
Gis2RpuezYO1N0MxMS+MkEzE+ZZF6yNSxk+2s1RIfffLE3Gtz2ZKGf03B3kjbAFD31GLaIRd1SrK
ap6nXyOSzkCPLlUqSmkCno9iRE1JjZtbFIu4QrVl+UQ19hfNB37heVzrLedKXNd7a5GpsNlSUCsb
c1P6li0+f8OsBUtMG5t5O+rZpTDVw7iwDX+X4zXo0d/Loq2SPYfT5j5B6+yaZCLWhDaRtjyijqWx
dUQhTmX40X7G4ej1unMEZ+mElHX+IunJuhR4YkrBOyTPSE1UubUCzHK8PmGqMSua9pxtmeAy28mD
PQ5AQKk7oZUiVIQt61mUmhC7n8wbTRtNbEeXycDLLzH1SHThiXXq8TbIzot5HtgNnDyjGNa609gm
CwujrqXfa+OmybpJ7labxDhhUlru0ZFtolXVITUpkbmrWKpDvqg0m76P//4wQVGewT5qvUEnQ78n
BcR2CgiFbbCraG7IkjpLlk6cirRzm7gAoymn2IWgrEVmAdfkVWF0nJsToFHNR6i75/GNATLAFQk2
XweRMmPHPvcEP7Wk+CQrYQ50BRGKDn1daGvXOtF/tVuLzmdsPewBrSCYW9ddkIIWIFBfBPVhD/OD
8WfHWm5JTDuAQQGzJ3XKb+5GApoyXtl0J+s0Kxkhq7DE2caqR7d0RM7FkUJ+2OkYCkiB7Um9lBOH
Gxgd71qUnNpghpy7J9tp0L/HHMVYUmpCF3Ls+OtO53hGRYlqvdCYn0C+we239mWINCYil1y97utO
pd6s/s/HsK5AQjyTiOHjVy6NWcWpFEdJAGxkHk7TgFaEpTmh2nf1lJsMmW6VZTGXO7mOhYK1a4W0
lW4426B+iLXRh5Ybwb+Q7wvCAPy2uY8rqi5BtxhwvezvZOvsTBFr/NBQdBIPjp3TS1qn4Jk2zap0
uLKcnrwPLRBLh6wZBF3UF3b48lfJ+vjPw8YHDO0MiKAGpFyiEyIe1ucOy3/GQClLU5bonZCQGmoF
dKIRe2Un+X/3m5rqvl8osO4wXU6UooYZDuT0UmJxSOgsGb8OAxWMWDLEqyrCTsgwKEN3+MeZjTtX
9IJyg4EF1TAArm3AsItM0uIOf1ZIX5Zp2oyQwp/H5Iix3U1ANcTDEnilbbAYJZqiUkkvEfkZ8tTg
t+ApJE9mKXIBZtfyOYpK0uVsOqXed4TCkfHmvVNr9ZhV+8jGS8QoHIrbXbbYM8zWlFqeVPq3kpNO
qirwLycvgQj4ZsFSRBPSQyMsTd3Ulp1PXdxJj+ePqFiuQzoLLT+zErElHljfQfLIyuEeRbfxQOqJ
emDbqASBOOtZzLrWZfVmq8NxX8xpRcb2oZ9UuNIRb6L7fuIJ/uaCPTO1RCi8dXzXlgAa0Vpz0RYD
IL2FqIsaCMFf5CVC481tx1PY3m5R/Bl6aUxCI2xZ2c/XxVpqzC9gaI/CPsXXOjqfNAkGFxSYr6tf
clT8uEl3TEIiFHSzriycUqD/6LSu9HB/5cMgSU4hlRn+H9O0yrQqFwfdZPKW+Jw9JJiyRMlAwOTv
FTb+nQ2Y7xYPzqz94iJIz9gtwVKj7zToaTlgWKAwyPouRaz0Y9lMtdW2fL9TN0b7j45JsQbrpT5z
zwsZMb99UK0ozE3a9aCnEWRmB2vISYYXlQJ+kzI1q3YIPQzY8v/LOTS10fX2+aSX7BsLO7xpiaA/
7wQGD7Jz+IdMrpLP1T0wBRiLRUPqWUqSD4nbOisOLoSbjGKr7pBq7SE7Qvnxl5N0n7m68M7nuCH3
Oml51gB7iURGSH+z3RNRrhDgfWZ2lqEshQQ531rDCl53fEbFUAHx/4n89jANnLe89Ot83NrZbvs7
qAI41+UyAuEu+Pt3px1fyri8so2W2I/0B6ALmOE4wA9Y1P3rIDW1pS4iqkYORZMH9aa2XFdkBv4c
YHSq+VXnKX6P5Dk4f6VvVCBDacK6lP4JzQMFKobBADeqGXOhgH/fKar2/aZIW4rWbJ/tX8GLaUnq
kcJ2F7z6Ftsh0tejY1YEWmqDoArjAVtGuCeNXIzRAkXdFqtvA+wnzFm5Lclh9vbGEL/z19sIEOUy
4tUjgbhx1aASb//RAVnqvLN8rk7m4Jt/0XEvdI90rMme8hjovawIXSlmETBt/c3hcY9Y93AzdCKL
kCU/k9O53u1TLxBfFFp9j2o2LwXZKJtaJPFXsS8v2CbYWdBNnILZKcwvfjIHHpajYEg4QPwL4VSt
GFPvcGXhyr6B6g3vHInNcQXINelHngwNgKwtqsOq44ptEd6JS2ryKSdfwlVPIOvC4uHvVxzpJRvo
VQ2ErPm396SXXgXFu727O1JX5Sa/aLEjsUaZ26QfAYy2yqBRd4XJIGEMGH+p7uwkn9aGm2KCuD0O
4oHM6yWVSeLKxl4yGLlRWTtJ5ixVFRulDEa9xZEF4q3qYCdwLHKLdA2DA9KPVpDk9r12e8KUdCsF
oK47OJRVD8K6F/MqxscKG4WyZIJTOwSTvwk4/zd7dCsguvZQ7+w8sRAnGgt5nzRlsbrqXiWHUnl3
88SnkjyDncBYElRsXZh7w42Z93D7aoZkUZyguLVpPbPuM38i0PFETMHWSAvjjzT0rA0l/GXvNLIu
brUM3KHXfBcUGZulZpIqLjUstJKyk/3Z7M2w30qKN/8FtPr6FeefNSiysHEf8aMpx4IvbqRwWO9M
sYFkMrO9R8T/96L3e6Hi8uhxrKj4WhIDAarIRx9XH7NnelKkv/VH9wcH4kREvT2ai23r1XRnDZcf
QorbXmsJKGyIeNVSh1ke7Zzo5OOQudNTj+EvUztHeBj/wgcBNU2dnhy9mGCClyaz+QniPQe+eEzc
hOt3ermGRhH9ZFybz5kamfeoYoEhME2tdBK5Ff4gc/h3K60xrL5bM8AmTU05Wr4YTk2YLU+F3I2S
xDCNAK+VHjT2o95IE6lCpFZmwSTVvWP+RIuKDvbCMfczvDlm2e67RSZiJw4rR3YnVoQsa2O0/R8v
7SlHJ89iNUqS/2pFt3/Yq9bpZcLw6EEwrPPNNhOsmIiZsGd/JGxdLLXBjkejEJGauJFo0RXRY+G9
0ZnElKb+LkgfVZKBpvXVHQp5nm/YEmk/NN0rrNr3S1/aBqbXTQmNqwUkYUzdFpdz5hYCC5kqr1hi
3KgsYr9XtXpf+ERmMk5sW4/Lz1K+ycfxnQUWNgJX7GIqOHkyzMGo4wyaX6uEPumNcWTHNMTtYjVa
YRyFmUkXwLqRGoF5ocLhonRu/TpLvLjqbnEzjUMCBcrEF5m+/qu18dsLgUn6Gd53oG9HU3F5oKSn
7Qk6zT+jBRTFjEfdg0XbTx8i2S/SbR1+Lrq8oLpmkLHlNMniMVkwFx1/EiKqs0BR+rWf0cemOu03
rBPgtwTM3kDDX0jErKHrBRFseQGFjT4RntD6uBlM5zwVgefwlpIhp6BEnBH8FrGpOV+2AmKxlGvZ
CNn7daGGpY1YA8SwI3/uURIwFPJT34wdS6Rr1yFL5FAxg4Wf0m/0NJtzkUpUt549W//nUyRVyTH2
F2V/U9A1s2nRHq1olIQjpY6EcyvHxEjhbXM2dr0ajcPVTYiEx3RQYxB+2sXx7sC7J4QdZwsJDiQX
b5xKjBGIzJRj5KuCIG6eJv3ffPKo597Uhfkm15LK9oCLoPjYBincEXYEgg4EQVAuBWMyCcZ07X0k
TAODvo9Mq1dedbofNG11pjNm+wKTfT/JLTAcOll9MFiQAqhp5HbgeZ8NB0QGgLrEKoII4CAt3/BG
pDK+TPZ/E5XiZvRWY8rHURx1FW19KD4vzXMqK4UhsDi6vEjKMzB/WvZcRl19/ij01l/x+eoqdtWI
idLjEqDwtHzVFFYTjUFnhbZXj43Mh5zeypI19ieEIIjmXxsoiVxR9MbrmGgEsNUEJenBqh5TaTYE
hNH+CzksqSu1wyMPg0TJXdjJDBswalhx4P66uhQ7pb26G0ha7hAyKhWJlkcEpOShuMu5FfUp9Lwo
lzJv2VgFnoXRh5zW7nWS6XZ6hvwcyXB76/6D9pS8dPNmpXPPG2xngub/rv9EbrvcxPjpz9NimKL2
IQ6xfEsT5DZ78limQowlhCwgBqCUQfiuSSCZn6qacrNLdzktaUypMEcTkQEqgLN7P+Ygxh9Z4qb3
vyQsuJJSjCc+ka/rM0QBiz7kwmKls9gEv1wC5Z9SrCOCDcI14O+wrkwTk1rWAK5jQVwz9g8V2frx
AGNCLHgjvgZJKy3ajATRV7eGpc825BZnyD2Js5OgnxFMEO8Jxxaox6r5bu4c+3IQGtc6w1v1GdRp
g6t8gtvb1jYSWdoCPQp/wOriBA+lkgUoQm5QwnCUZUY7XfLF2yguV+jB7UgZR/xt75I2neQiFoZs
WqMlVmTxGWC0pSUAlOLNTGS1KwwLX9U2hid0W9zXJYwSw3MqNTzGdtu6HfMX0d5iVGqoQymdJgYr
77/reiohGxm9ombqFnNzV6ECeD6+Gc4j+Fpdj6qwdxaDVBuXnVpt686/jpm0lwkn93qjoUUy54LL
LdnBVwtBXRCbNZo0Cc0/MgcoSKIie6UugIpwdKrhvjMZQSdFIBFx+TxwoziIpJqgq1J/EVP3hdgq
6uiLCQCVjC6c4e3PegKbFdJwpSJtAOF5eGbSRDWnBlnPeSAv7hJU48+M4egGT9mLlYxz3e1gwANf
eV1TLJBHlrqM3orJxXYmA9MtKk8ATn4HCXwVKYr8mmnNs7NrT9VzRNRXpQGrRGQPTZILsSfL4ma2
hvQ99zBIqRiPKCgCiB/UYYx+iDsZqzY36Kkn7HVo7oo6lLa/8W3xbaHXTNNB6kvy17RJp15aIoCl
vWHWIvt0avG/cfuhjv6dyPg/27mfHkMBAr7nzCrQLgHVHrTLZqf0wI3fs35bDMyMc9nvdUG2jsxD
l/LPo5YM8QujUhqQPTjj6FamuPztxm+/zt2BircGu98QDiaJHU/h0hks/2fguCWo6IIDpdhDht4q
5F7BOWFDR63v3gaI8rX5Ar9uwKO8txq67FbIbdMVFof36BXYt0XR4yHKOn7VFjhqktZM6Pcnyc3X
EtWS17J6u/wUgpvIhJB9f6LwHF+6t7JU0wo/CCcOw0mb2iK3p0oiahwo4h82Ed9ufL8c5BcbFFBY
5KwvM7w38qVvaL5zQfiocPU/dOvckEnx/1wFFYP+xNxDro5sHnx9OMRlHn3o+MzthHfK52GBclij
YentFaAsjH/O41QMCIUz7dTNaIIOaum1oelZtOHYs1kQghaioVODDNL89+u4U0ozwPz8u0/Sdhrv
6S2CqZokNG7eWFBHXXZzJbPPlX1ZZEDRplGP71fbaZHlCfVc3vt+he3lkN8BzhCNwo+FJbZn0Pej
mmZn4iPrVHkt6XSKwCaxEwcIur9T8ibOeRaBFuLXd55f/XbaUUVqM8ZanDPCX9NZpUtlavVuJ8t4
GVzO5xN3DF4vyG5QaScX1lD3Q0EnWAX9kTStYYIGI792GCwv83jU9qNR6llNE3MD8Wup3yU4NFpd
VVWp+BxDj3xXdym4yzvhpfdhmfOdFjNiUZdqy7KMJHBdGLjTiofLqH5HG+zYUn4aywICEmAYrVWP
56tja6kJ4ypsp6VoEO+zJaLEopczsGVVvQxUjeEf91clOJLrhilBcN07sTzuweoB5AWlJyWswV+t
36xbOW+ldzC1dcA1N/7qkiY+vzroYYMKv0lXQs24SiWCL2cv40cc2tIxsw0l1mlLaEpvzXYdmCaW
GSbhEdCbEqAWvqoDuNBW/w1g00Z10RitcmTD6fwbHDlfRqGYzlDwxjTGzDmO0y2XctzRVwpQAyzj
2K+8cqWzSnx5tsLzmOtknILRRnJIfgV8EVXzO9LAKeRmwulG57PhMy5SPOch9ho2ybZC8i6o+sFT
JtW0blW4f+u2gAAUk5wAzGXmHiOr4SxU296iXX4ej6d39cktvcJNrVdGXmMgKtORBFsHdkugK6h/
oDCfqw7APADLkfN0J6X/c7KgZzJ0UplQza/728ezCQlAD+O5jrV6JwBviUSMPCNwWTi+rhl7rYmo
HSTtGSFsO0GjPs4aoQLqbz/zKz7CdTdTikui8EuYcMfO9BtiicTcbGo5gbAvSl7wLKke0j08fXl6
nEThBkfI7dVH/OCXYK9hZkg1VmZlPA9QtB/8e/PC1Jy3d0fYWnJZXIzl/P64BSUTYQP01UB6//O9
pctdFsdwAAFcx9fbcp5IDFpwyOWZe8k7ExDznlDtxA2konHQroLuWMLOGqsojCm3tHHPJ7wBdXVW
V7ABPyMYr9g1X3OnltxtmJtleQUrEJ9h3SEVJV/b072ovludut2L59FzhZywzRK4jSXfGbxpudzh
jVmiGbVxo6IkPqPlmm7TYzwKsNoUkpKxQ/zpJKMtgfByOb08SquFhacGM5twUIITvHtcvnG1UquM
2CPSJsX5XQWsudXL/X8PIHowy/V39J3IbeFqGgCkONRqpbLyk3OdsUE+bLMvFMhITana8r8w11Tt
/40RBZMedGxDJqGWFZH/sbD3Q0GsnEPLLAVDEQp8wJC9TyQiluemAOteB+QRhpP2nOolKMEbbbcK
cLpPhREofnxDRj2DDCO/avVC/6LhdoSTaOqkMVer7EEPyrt/A4Mvwez9f2YzNCbA/4qVbZeYshBj
8h0+cuKeCJn8g1FYc3/Av3hyuuFLiD2JUri4QKv8sSxYT+TuMJ5lGpZsjPMVehhTBS/SMzVarCoB
GRk1YvUdU6jIpWxugydDwerM7Q7V8J1EK7ejkCX7eNmtXRJUipns5WzzCsoPjVaXsZmUthUNzFqC
6mWVTqrw4xyfW6tYvExjvKbEoDFJqL78veSUCOVV/X62AF0hpISvhOspc5ZpraCHSloH5qdk1yWX
pBVp4AS5FwEd8wO7eLXuXwvbzo3rY6tiDcE7xPzRI/DP5tICCdPa96tZwX5EBwJDFWWcPOFnvOmV
W0unikoD1yD0hleVHfZu88g3PGOkPv9r1k9O3egcd50ZN/uXrU3e+twiamkxIvcKup8sjvy1FD7Q
y84ZYGiUDJyKuP1QeQWvoghfmOYx2OLaaMziaPc5/+UI7wn47RmdSBV9z1E2xGX/OLe0xPnLpPM9
aNRJ8SKA5GtTjxBkqi8Aha2OjSOJsgjT4KUOq00TfYlcDxZupAFQ9HxWjJf/Z4KZDLbMpA5TgHPQ
ei0IG6A2+A7mz0axb6xoYGMDy/noZFHMIVkg/ClotlRJ0joGXuuO2tfrtoXy65etcAfOOo1PXKoL
7/Ah610GtX/K2qgjpmKgxv0YNmGw7pSTxBKcm6AjJvhRt4SbORsLli9lY+irBtSdoSotPrSjZNl9
wExy8unovYif4MkdWjI+Av82jVC17j7hSwo7z9sTriBdYUj1wnYV6ENLPHgkKCcDF0qmbiSv9uAa
xG1+XbJNwZb8FiA+geJnShVXQUzc2vo3miSiy6B2mVcpOKuZ8skIWkQ5aNXo6wljNvI6abhHsCf9
9dFXYGtUleTzf/XmCuV/3Biaty78Jze9Hhehab1tw2bDXFscmX4dprJB/KEJHpVNUav3Hh68PCyv
JTX2t/0G6ToKzaOLVl3Qd5Ga09bbaw9jAXcJymomw+S9lqraC3pDAxImS3pllbpqm0Jv0SmYpWji
R5Z3kx3baK1Z43wyeTSM9wZT5nqvvieSz8LSjHMnDDWMQ9LLnKcigtPmVxduPMEjcceWQpG9B1Qn
s4zfXEKsc9aHih4s4D1k7Ufpy33CaWqEfOLcLFrUW1THJE+NU3C3Hx2tX+zGZiDsm2QE8pFGaX3G
ndJjAq3STNjLUeIpRMk22IJTdKXfbk/g1JlUI4YfLYF4khssTC71RDD3GJto97w5WdV4oNqwS6SX
qI8EdDCF/kZ6Pr2QGMDYW3ouXDcUUidsGGBLMRy31GQoGFqisv14AWwWxzg6pFM6Rl1Kpiv9jBEX
W1iPShLXjfZoMYC3fyk/FbBujjcjPP6qfXPoIq3RYJB+GOo/PZhc3RhZCoeyuZr5WcD/USkOoeMC
ijiY1lCKnC7b/RiR31/u0ARdhoYieTXMi9ykuTv/Jsl0erNI1/4lHWTsHSOfYaGt1EwfzZyYhOK0
wPgNJ7KyojzwM+QaVG7wLghV6DhXqYESXbXth6gA00ivvrQUhoRRe9Y6/+EnE9EKKe5d0pi/mqJK
B5Ey9Kjh9cjYudGeKzkQpvJIS6oVVQawgyWtXJQQHw1HdXfSTmB1DJK6DA84oeHgOL173hBuLXBX
hCuOIj9/EQHJLdadWUAmS1YsQ9sHipNqJafo8sBiktBUu9IVSf1IzgR+H9Yfh0ZxM8j7kBaRI4Jm
CU1JSogm9+mCMXy5DhREB/JLzBtCOo7OOqSDuJm5i7uJTuJgKxlPGI/WTIBRKhDEfFtC1ZBDG6DL
bP9Dsej73zf9FLerdw3Qv67KcQBJMoj/UK5bOWBASSV8jv78zSFy5g8UQnIRYUXfe9e4HV3nN/Sp
LSK/eGeiInBB73VJxhSn6BLXa+KjA8DaJY7FUotyYJglqBiv52msGH96mL6ppioixzNPCF902VzB
QrauWFUYSV2q+RZrYq2YrjeuAberhXTgHHDTGSdoSXjzF9u/mFlMn8mh6T8DETFg/lRkv/UUHR6z
UmHA93LfxFYntJXtyst7OcXoGGhMZPohcP0Hw/Fm97sNLNydGBLApP53/Ts38xqA1/dYbE6lATiP
fi5nyTHDWpj/34o3vbmEZaMVHgtnzNkaXgq7+vmo3d274HUXYCltez2MMOBKlObph0REJpUplVh4
m8ougT2MPXAXMP+hVDUmh8gkwbZBk2g6jwr3bQwcOFzqTNu8/+Ik+q9//IHQAoHk6ThUXEE6/BJn
3atCY50B3+aQzmV6rmbC6e+0j3DAw4pN0eQb+R+yQutFiVIHWSoyVCL1HM/o3Q17o/VvN1dMvNk5
I40qBF/zHGfVhvmxmyxxbO4nTavl1z9RsJTo9y7bftCH8DLgl3OKh209/1wHceLrGP1zBCkvXKto
8MQ5kBNLA63csVQRdbEYLlIVvJlB6CREvZ2SNG+lDVxlHdMeXQ2DzPZ4SY3jEJSoFJ20/5z6PHCu
Tr9hYRuB1SGdlt4Rcv1r0JnG6i+c408xRULr+L5WfO+r7C1mjh0ar1d2P2ILCfZnowvxLxlrdhtw
WvKi/4oxhyD6HzbTLORTcTGXlMQ+LeK24tth/OYOOcu0s0J3HM68W1mvhmoIhOhd7iviwVpMOWi3
zq97cwY1t2aWvu4ulOYwndrMlYtGSB9pVmLZNIp/gWrcZY6pKd8+IkZpM3hHPEubgfAqbifWnCjo
t1tNldV8+USS3GG2aiKS2mdjUtTe+k3S6WUEpaLvECQ40yu8enPExjAmIfYVvRAVCBhCTMUJ3+D0
r1TwaAdDjyLWTezGjMT2kUeTTTYSqyeRPBm99TlXgq1qoLDQaFLGSCjmjzT+a4Bakw2OOS8vcWgY
LRgeCa2TeeK3INf/FrgXolZ+JC8ZVy13PYfN4b6Mh03te3A14sppgs5pSziaS7WgYy9dVdCzTv4K
pi//OH4OPqArUzHvDOjHv7lp2zNAZYz36Z0TBQx28ugzsBp8ECxux+JxBObmL6qM+jKUZOOicE1K
kGEfHSGHz45/ARP3TI/70uloOEpu+3BFHjl7C1Ff7KOt3oJbvN/cR3ZSlGtiUvVfGT1dxlsTQuN2
P1b2sd0m0yR76j5EKZ1aXqb4+r86rZnP+2vheW3zGRJlp0RgmPmHU0c51NX6KIVfgw7nQLN4JTzl
dxYO3D2gML+OXmGq1oFSUwL2vOTiUhuhlQLHEg2f7gy18v1ilsgNuR4XqDXtgL/5SF9/4GOl99pB
EJkpL3xCvK6hhZPV0uACtC4LAzImdYLs70a36aWzm0MIyhF5PZlAMAwwGZvSjC7KTx8RQp2ARcH1
iA0Qn0qI8TJkGQrJKbCUhzhKoZKNNjMV+Ue1gIKV6AKXHvKWQh68oKnOjBHUdLCuuucxObr7kdO2
NlqKO2KvSxjJLgFUdf0XB+S8UTngIIFEpee+MSjacPRNhg+9+X/Y0XEFeIaUhA4u6CDmK2q6DN6t
UmxIHZkRdcDVdkclCpONkLelIwl0igHfZVgpRrwObh41ihwukq8aEbNBCyzISVqS+ioKOE0VyXzT
/fOn6w9QjyK8/i+rZ7qzb5UnNyiAXio7Jk6RYfT+oxzxT13V2BtUaZuZ4Tj15CJYm1OdiZDkO8g/
SQ8xWVlFiEyLGFRT1i2Z8cy7ve7rqPlTT1kDxw1++gbDJNeXKXh9EQVvwOKoKJKLJ/L5JV8JTil2
CtCQpL/ur8NWvilRDvSx7aFwkCJnI4NbwesO6OeoBoqnOzv0gB7tRNIbDn5crorMWUNze4Cpmo64
Ob+xETXwNKa2e2a4HtQm5lqO801IRpsAAksX750v22WUUj35AjFXWi/ATfQdPM8sxCCRmHoc7AqU
DgTL4Ggic/n2W+qX0KapsFdEP4MQF2pew9PdQXxC/SZIVrHyljWS1J2gY7FhJjoY9ksVhMA1FJn1
mTlJjSY3VLH3ONjeIzho7ELg8HuqmThjNkOwhLi1PCqjRQdXlG1hPR6TLQO2W+TSlTXwerdHDVGs
Op66DgcOumquRatKkswD7uLgUPEeJk6EFryPmDEullRs/C8lcKuFiOSOV2AXsBP/kjtnMUY97BNB
CYzOZd1ELoOR3bmo2MLJZyGzjV9gbZvQKk6A6onNPe0JRBlyEx7uYs7G+pt6oi5OrnV1s74tXpWb
JqU+hkjMt6TFgzNn+Uz9EMbxxZTMNflV5Wrp3Gxb1yV4QxsvUW5WlycWppHNfihno89U7FP65aO+
TjD5yh4bxhY6kr5CMbE8ikwanlvvc/X8xSyVBVZjw30Mm5gUuKiJGCBYqURlwlT52bFzTSj3giLZ
7NJ02qN0LAH+Uo65t58ySjSmpwY1PKci+IlNzO3Q+hn+c1K/gqZHOOsV5GfkFYoHDa0ycWlBtvL2
6HgkB2eN2yBE5JFo1WwTpCXdfrROIgRxTKkTot+kCic9gTYQnGGdHcHhpF2eqU2bfbF0cyXwySAj
Kv5KYc3syS2jkLSWNSn2Dbt55AK92aIk6xKlEAfQdtsjCfv4RYzcN9x78enEWgX2l06LN8vNO/VF
LDJJUfUxvd4zuHs4XwtgXkILTvq42XR9LI6bbGirH8gmxriFBxMkclQ7vXbtQgxfJcJ/4SnBvFf3
AW5+LGaWP+IIWXb7dWZ/k6RuOtTs4HquPc5RF5jm9EZALxiO9RONAhRARABD0eDZdxQvFzQtnFKd
jl/x4DuDPh7VOMJ7qYbm/3x7ACbeLcJp6cWU3zlhBrVRP/tgzdan8e0BYZX0OTnNV88BFhTcYpgd
O+86enMjJ3e/h5a6GPnoq9oqpUaPafCQmNce0Tdq6UYSpNzOjfhZxmnGC6dVbxGCEODAnoOlBXPV
uZpzj1kuMZQ8FVl7/ZoqDxVlv12+UKpl1sLGXKJNSamvme90rqLp4yhH0OWj/nd3INdf9uVxdWQ/
1v79+Rgq9AS3C8gkfrxNDRdQd3w3wGIDEtqiD9l4x045QYJY3MPxH/qJo8IWQARo2XHeIcHXpmJK
hIwcdVzU4CVfF6+mAfHJK1fN3xCNK7Jx5IGrodqekQ4ivMSCbxyjJkWGpaVyNXPbJfsVFsqe2Pas
L6I9PO1Nhy3CwBTlYKJskThU8gBt0OInSe682Gg92iAPFuaxd8MzRMnpe3lUyGUAEQnOEIApOYTN
ebOZ6ECI+VtqGYvFF3DxWe4FElLhCDwsRkGQHCWLoDkia+iohqz1m3hN70XvPO+dymzVc0U1UuFQ
P3rzYyeX6IU9qGDpSDvM13wS2EI/fISXYgsLujXFUWCupsWgf0uhTBQ6deGyc+L/Uwrp4PUsAQ3i
/7lEWkgAEffXI+6HIOOeMAH0RRHa6wyr6dePXUagV6Yn0txkRQVOfwNp9MrUhRqEg4pEqt5yJ6UD
eMnMDJJi7NBE4JqbMFNKa90qPI3H+ZQPmzJHP/ToBUmxbVtl4kh9abPGI/5AnpPzvQ14+wM7mihG
mc82lmGJTS+uISBNzcMGgiDAMU6eesuxqikR+2g13v8oQaHlUOUsbx/N9i+qQ8gfUFUtrQCccYZn
dhbM726P0YhvO8dd1ohwETYmt2jSUNG8u/6gIWf1BzAd8mv+77wzm9qKC7Ss2X/e3OBvM4iO/4rO
6KjC34Ugtd1Nhrl410DUsJSxpQ8yeRBu/5lt1xaLEK4u333kZVdf3OxGdUyuhIEJ92TCyRRHnZo8
+LyiB+FdqhnIy4TJ6G84FL47bCBCecnhCkSGga3aJmN6tWapgdT0DVhrcym/XcxKh+qTqMtCa8S0
72d/pWLBNj0Stk/tPHozt48f5wShjcsiQjbTDQ2MWw/MCBXPC0lonB2zFGt5ldORGRIqtj7xx9SN
FFxckrbc7nQFbl9TiDPcuJ8EsdqGFAzBForJzS3hvuwl6TIOZ/ftlnYOIwvZJE72MrVyRe83JV+R
EUN8Ve21j8RFFQHBOrIRusLmXXwmof+qKggdT7ouXDp41U3TcoqGx/ADYsI/uAtxRuPs2mgXj2+i
j5LIE0sBj60BdkCZqrBQQdKsSaP3NV2SmbKXzmdqhZ92rX/24wjQdykbhP1b1KypmC9Co00nsJgC
dDV+TyZ2MkZUXrlTBtz0aiRZyKX2XgMlYDzfumBnTQ/Y1bqvocoJnMQk8lCTUMXhBkDUzmFUX6nR
fq3yF1mTeQEPAxLRHSO/8gRR3tMn9BM+ospGnFezfiYLYeLP1jd3oemWsySR863Q49X22AfGKuAc
js+Yqn9oOPFrUxoiQnYcGDAa9MUheZUYDdI3LuyP/FJup8NdRCxnCxmsPHKMWs7uN0zGUkIaZhuZ
wvOp/EUyLTzTxcCpPxpRiGcySwSveyom0YDZT/o2U0noqId/XYxp0bQsF2WxUHZOwLjEX6V/BMyL
FNihhe0hdIltXl5VTJ8W8AqAuEghAkbjTQShIjO40kSlMLLDFcxlpkx77ykl2E6CUdGRFZchhaL7
2fuOLSBreyM9kKQ8H9Br0lzVy1hWP5WlE+tn1BqR6BVKmeF36tISZ/Tm07cBXnZDhmiYujt/v5eC
VGqulP3f+JWJhheytKsm1o9SOdtKxk6Iid8viS+RUR3Z2BrNKwv3npgM8JFJSfvufNAZn1HsSC9e
BbL6JxaJT0iwsWf+QytG/IMFdjMa+CTsy03AGD7L5y6CVxDu0nbshmfMHXfWR9XIx8xJiBuEaLHB
TzMY8Fc8Dfir9zuaeTaxDH/2UIStI4jDcEZ56+esBdDXRkGEmSjxMcBfe871XX9ZTfpdiqmPmu4L
Sr9n49Tei4NDD4dpq+ie5GG51x19vyRV8aQdJevPJdHCLlb6EewWt0+jg5qQLWtmFyHvuUMNKUOB
/flYlKN3xpLZnWm19w6L00zm/y8JycHAu58YM7KJBvEPFgqvu0NdOMVhWw/a1wm26xQeFACmlwY/
Gt4mo9bOKV1gC7RCgAMvgmifLiB7Gd0rVbzjcwObAVZaNunztF5kcdWytyvHcm13NIL5H5pReJAx
pizlXmo6HBWeACP6uQdOwAVnEChggpbVyByuZHEXtNEPq+aUGLga0XlVCAlCBQWhWTqfwcbmBIru
koJazIYtfdgOlRci1SuZFMzZdnCPet0cqVyho+4IOsNogwaBWxajUWljT9Rmo8A64YsEBwAHxYgQ
ulq/tElY4t919dE9Nu7Byv04TIBaLqk9rhlP75E+msvWUhPyzZ+0sQsrLYWlbtVyqmw657Rg1bjH
6ZyScJV35CI64VV2uL1l6GuTsVBV1xNViWBxQLmOFR6pCHLzrUlrpy4uoye0h3n+gugJF3S1331i
byMVY3Lfudef6x7f8Fn39BRNlOB+7YZbnTFdT/CFh92VB0cG6JjVoN5w1GwxuLW5Nj48XeIVp8lC
yrkiKxg9GyNNvfcFeUkdLvXbTHyCVDgFz/X5u2ZyHdf2BtTpbmOFLCFAyrlSbKjKbpr5IgLBti76
Du8w/tDbZHuE9HFYMHFnP9vZgS7qJOHFQYX+qZvAbYHHxOhPuLpzh77JDo+VgLNWzCgNJ6hwZDaj
VRPbpSGeHDg5fUVXr8bWYF7jzXD9zXGVHYiJOZRJaoisxH/9BxaPEIW5+sReZEXcBMUI0qEY8+Su
M9e8xO/kyZMcYYD2957xTChVJSS0fGoQ5Xx2qaV07Qn+uajBjwetWjiRHWwKJqBPSGu1hIHEdPQJ
rDsLLq6IPVXyz3HHwESgYNAuat7t8DRoKt4Y9u72uwxSGnQSpo7PMKte7AD2gDKnJXbZJqZL0Wy/
3pcC7QKqdEyJjR4sO7CraCQm48w45MAKsKABDFIeOw3/6SG3JwHvQftQQ4hWcF6gJ0hXc00NtIhY
Jh+YgH6OiprvpeS/MPMZCkLTnO08WHxWidJNQ4Ow8ns+7RFuQVvjmKiIaHd7LCn157FmTJU4BmHQ
S5IstJjGxsCEmdJMo6xb3inx+z6MoL9lD6rnI2Lr3UQerzh/+8ve+8jHzJphtl9JUk/JoB80Gc8q
ICA2tf3+ozJI3+H7O4ymiKVYUmMxPHkQ/WZk0sHRwDUz18WU46e3QVFR1tioRk4moZsrvqxkbuAF
KVf/iGPMcuPAPnB7WkOEda2wEA/SaiP2DPONrcXBpoZPSLshJUvBE0fwwGzhYxEYcFUQ/V5pFzXQ
9zIv3z4oexRcq3BN/ok2y1s57Ry8RPoIyOcrBA6Td2p9AECZAUoRPe88HFCsiRLjZqyNR6gl453o
wvGwyIPrA99RBZXEVVLjt4p8EZEULALsxX3lKuFktaH/w030H8x44C1H+OmgFNBYKbEUXpdZOLec
sEw+fFg2hNT2YIE5qdECNcOyYSei/zIsA52LopvqVXxr1m6InFF4/ySVwY6lfVokISZDRL110x5h
AWC6Tre1UNrMRL1wMp761FjLVWcQLVIQH91iNgNrVZsokoGHXaWURO8Jb/yWpLDMg8aVdwEWfoOP
nos+H842Qz8Oiv7VTOSAmJB7W8Rk4zOT00rIZTdGJ0yhl5uGikDQXZDNih5gyXzFE3gK4wiLQvxz
p1IEVdLbSjinfTghX8Y0bRax+Pvyw4fiUXtBLiz0HU6+jizV+lx5rsgFih8jp+ynnuMW4cztMmvm
XAB82Thvb35LB+zTHFPeeIEsZYtNswqDXGGqjVfI06FPg0fV34/CqzlWTbnjPvVo3N1Mde006oMp
AHPXqmTmnm59dHHBxW1+Rlrx13ZS0U0yQEQHh813UC+YkcagCPEDElcEPGPxWDW7Z2GGkLvJzG1C
u/Zqrcmmtu3oM7OtVVAyYjtjm2v8fDNnVn/RWeqEP7x7gmxrtunNr0j2qwnyBHAuD0oRhBHrgeLd
9fhM+VuspwX51zkfFIYKwQFuoDpH+WnikNcWlFJqIb6C890QiVSXNkAvHOXWKcVtBUhpmIQz8rrG
l88qYniNgAmuyAUR/9L5Ma/ckAb0boIniFPY8RMtFKI56DSkbbRnKlZxwj5ojIL/xvzfgGwP4vma
G/uWttWSd7ZssN8CrK3dl8/1d2bvCVQ8mY2ovfAkanyIMSkhkW2aNAb115Bqhbe9Ky9jE6v3AKjl
mfINJfXfwCVHcdD41nx6iYlaH2d7FBb4H/DRBDpegsor6SdmwtIF7zLCXPtcMuigdZl1iofb1i7m
XpviFoqlLZQg6yJ4H6nk3wLARb1wB7+d+9bkFOAH81ELz7ESWlg6N6iXbEzF4aoyojg+pyNWRNH9
IeZF/VLgr+GX0rdbU1nReR3r/A5bKqijRb8D3QHEexfZs4RhVnkH5FyrpQgnKxcw1TB4PbFQQHpk
QGTKBE7hj+ESW+cJPaKh/LFc9I9tLLUI0gNUY4MIz+DLwAWJT84wr2teiccIij1c80YDQs0cgTXF
P+gRbHO3Gk6bbe9O8sw09s33gOm95mplw6zbsCQPJ2gn3NHEHBG6yoUc9c0GDIHi8RmlcjpFHowf
cn7f9ZD6veMtMAn+dM4AfwLCYB/DNjscCoviXPXNxGlGAFzBhP7Kim2ET5LSYa7wXKga+pbvf52y
JATkx09+aVXTsdj7MpODUASW0xqAz6Zf833j5F7q6NCMwL//AFSWrTdFzsJr+ZYxrSC19MbG7IEI
KKOPvGeU/xREHaQUKQmGxH0tsJBHf0M8S6zuL/oiwVbscVHGfDFYwWO3aMXRxA3oKuDSJtTPbLvr
9z22v6xwPeTdOWnlqjGJaDMu8nvY2BhZTEWmPgyjVWVzRmXjpmjAxHitgxZEKRN+DIngN1pVvzO1
GchM2soRsmPVh6e+fQlp0nnlBIx9Xw97vNm03uSLCjom2zmAbwxapWhGl1WdXJQBeIf8Ba+iP+fN
RO1Lh/B3K9iAjkiUpbhYV4uSefbcz2aIECjvuhew0llVnnU12Cna+lIg3Xad7RI8LJCgWUlNpid4
vnf40EN1ZBmSer1XrIaIkgO8BhZJYhXUVfairte5n8dA4UEkDVXJ33IXixLKKxCjpvmOhiC09wPX
+jfizY3u4TYAFmovmmPl7jlbmBOayaBxVFe5eBfOJ45AEIEhJz+Nc4cWI3xOFYqtlG6lnU2UfZSY
0Iv29KeSyuZRKmSVuCcxjqfpETw52U2jQP31YtGqmpw8Xy+Sx+XAduA7MYJS1DIW27fTKHuFtXbP
/gSIfyLUtv6Qmtm0FqWaBZ55kF95x5wNIFI762B4r8C9yfovAMQa5M7r0kJIlmc5Xlj+dnfxHCTk
mN8i57TnaKlljYTLR3aAMTiSGdZvK6qhfGPnG9OkS7pId8dYwlDSLJZkljmShZA3w8wOCKpp+1FR
hhZHdraAxUpef2X/U5InYRM/5ZhRl87O+9nMsdbw/QmnEmzAYR3QAQqp7D6ObPQqkkqtvgEjXeWb
wqxO88TI0B/vj7v7A9F+UrkIRjSVEL+RslsMm7+TOIwYvKGawWh2OyBomY+coneZ5GYci+/7N4KW
JmNxx70yUJMh1iDHZknW9+fFa2mkhtvKHAKa9ee30nSIx1Rpj48z4S/LjORcmZswKffuiVS8cS2/
hqYDUWbtqG0/G1kkrtCsIQCXYYlkK6OEwKr/8CcWVkYU+sera2ZTNBTLgybbKh0FHSQ2sfIXbg6c
B7YJ9X840Os7ecMV3RiiNnlzY3UrnJZumXdFR5h3Q16rIcdZEAEGzxrEE9I5Y3kz/yDUUftj1vq0
+q7xU59ohnXNk7lonaTuEGXKb9FPUc5K64D6daluayfKj2ajEe6zOsBAYuEouj4x7Zc8SEiwHja3
O7a3ppKki9hR5qS44LqS7+qppkw1kaPe0xYenfc80IkQFvPCR8U9gBq1jA6itLY42sEgk+1JJ9rA
d1ixzKWkWb11xRTeogVlCelFPIDlD+XvGBtBNyk1BZa0fSBKQSudNTGuwcLrN4bElujzamEtzpwZ
WtmIlJa3i6nJN//Sg9xwesLMGXUbP5Xoq+9mJtxQAkMCCicnKrp6oa0u7JaH8IgbJk7pIZsbrihX
6lMSbEW9pBK3MtBR/0TPZAnxBe/lxpmmJMxeOsQYkDnySmtTPTmWFArHfmgeAvmzxFB7zeiFUiTZ
YqzP1XLOYOZMHYuw2yn0dsazH3lW2EGf4VF2JtXymeX+LbEzm4hkfgG4gJH3OOImqVs7tB/RAXl+
LIw4f8WDuu+1DUEL2W6tnDxV5XKdMiZquakkGbTPz6oM3CFD22ZfkOYNIR3enuj+/v8xVNyyPfv5
JarrWjCw2cIGNl8ekKER/0+J0HmErDdYifqY+u6aFeXF+G5PNG87y0aNU1lhp3DwoGlwnqzgJKNn
XghTw4b1ShkgJK8Wdwy/IiVaatSChv6dQhE/n5JpavqiBJtQMsRI3kuJCf8FiQEmKVWUhjYXVxZ6
qtx0hFQTh/siluorGdLHBYMpjkPy4e9BsCdVuOEJzau3f07VBjpaPC2YCoFVvTaTj4hBrQHwlDDs
DPAc8v7AOwGIAgFaJpc5vOt328YNLjQbZ/Ul8+8orpfaTkfmr/57/ggWGMEMfgzeW7rM6jZR2OmT
hq5u3X76VKY8IyEItzPfKVflMIQGq4ZVhPNaEsWFQj37/FqNyczvRL774dwpWrV9UKOI2hiBfqzV
fP3UOvtI2aHqBmbR5qaCaVdVk8W+ifjpDUvwSvfpfXY9nVp+c4RyF8Fps984Tv/ozrSxnSJg9x3N
6TTbT4dgYhOm+LMqJPtRnctQnVOVUhyWQq+WhHj5I8daZxiAWIQkvIaUr0RRUaZXfJb1L3r9xbMf
n+/FOm6NCf4pLCKWXIlmHnQOiJPiXES6PlBdeQJW+AMOhddl/IFs7UXWAWVbF2uhdC30v1QwO4B+
66045nFhO6FXVBzoQ7vLDL2n8l5HHRU7GFExBlPtxW/ZGQXTDaI4nF/GrjcaJ/WSCFp7CN2GkGfK
OZ5t6nGRuWtvwu6BpX1284cX/wFqK4k2dABamfvs6DjdXJPpqElPzwXinav0H2ujaTpzCYMmtvfV
CXTOZ9MWMR6W1FrE9AHNTQzZRm42od5VjPfcvRxBZ/fY4IKrMrRRNzfkjRoEBFxhNYX5AexXwWIO
dfjK8lpd0doZN3khi8X42ypWZ6N2PaMHrFr5KXgCWzPuJRNueTjEGOrVUIPlwfnDpdeRlIbEGulY
/FoW9EModFm2Ol0E8gfXFyJojHKYLF+YHZt48q1eGqU3VPgY0utZygD53dU9SwzL0KKTdpPopeE4
kTc5nT782NVAK+xo2qsX3KcsHt6H6ws79SY+4Qp8Kw3IFKRELuNRvg3+4kuRd368yX+6P+U3qD5J
UnVedWAY3BTxbxFvHgLAnd3pY+USSJe3DH6P+xKfdsJSlSpX9DjejMZptNiu9vMfzAYwRhjgPrCO
gDq53IkPBboyjcXmpJVd3EJuQBrnkG/2oz1hvWX5wgqJ96mEt6uJjJPfyN/vHI5wo4Vz/wr4Un7W
tmQZM0FuNfyBexwAFvOZURdUcyEaxLJcrAiBEizRhPNXPQ3k8LTGYoIJPsg3VqBSlhg52gNJL3UT
2r/ZRO7EzbVACwy4eo8oh+MwYNrwsg//mlBmnhteAmEhp43DqNE8H7S+yIB4+gYVECCaSdmoYjNO
XU4/DJlzVZXdTynQZqqIdb5FBgwe4n6ZQEsEMrvbiQyOaQbGJ6QeDDBlHhbv1ugtMyhOCRTZNGRD
A0w27UYUxXe/gWwJ8ZtqGprLnfM09LLzQn5HmePLYU9iwd+JquSuWss3Dj7gBUCIR7M7a+m8Xiuk
f8k6nZuuSbPdtA2ZpXaRzas6W6lGHdRmEJxFF2hNgvUKx0Qpi6QeGEYzAlRvqgHbQiJMWPeNxVVO
ptNuGKkze3n5A4cOMVwmADAtiLaISyzwd5MPvqEiza56kpw21dQCnllc1cNaSKG6EW+adMiR5r86
a0cGb76QCU4DMGHMzJq8plJ3LLIqpCv+x7clbmtVTiNN2kDf4qNbcy7HETyC32EDkTuJ5cCwumdv
EhW0FL8wuS/t9vCd9OxoXPlH+p8H4Qx7xObfOnikEQcAhTUq2GaSrzJjMqUTGy2CbePVWXJY+MdI
LB9qYKW+0p8dW/tAB6Ftx0wam1I32enH9m1N07iKLXRZsBXhgUl9h+q/mIpOkIhWfTDXStLrGUti
owciTWew4Dt11q02hbmJgRMm8tn8ymhCaIRvRr6PUUKw7GoZOV7BBqerjGGxgqcL88uWFAMrslpn
xjrGInMzaSFLedYRUOJzZwbKMct+vtPSnw0Hwjd8kFnTb7dLwnm+fnnMfvaeEcMLd8/1jowj5YNq
8kgnUZBVtZ9EUihCFbe/Yw5ORtSnoQCQ91E1/+F+NznbEDPv61RboXMzKwa0bTuzDmXgBJ2PLbYk
DdI5p/MTjV+AjC9XjnHUOKPD41V63WnFyHduxjxKHoGedcv2wd62Q3XgqRaYtQKfDECd0nphDRel
G5o5yJrFxx9i2WWBz4gg08c4qAgg7Cp2u220rOCE5Iz74XUUGlRnAM+cVCojSTv28WnrikvPxf7u
yRqXDLDT4MH2rYJb+8pjVCbL7Xilta4T0OlrxQZMBGE8gsKxlr8lf+rr9ChAxZaA3Xvkk4fjxIbp
tb9cPcpwc3ZnPq+zctLMgkMj1LE8lQ15eiTibN+iqZtHFBt+sIBRgV8bNG8mX9rPLeBYFPCyX212
7dWbTr6c42xzjdzXz27+IZ9M1RYQtCrjk3VQdEohX/gA6qYIySuQ6rhE8/5VDhd6qCTuzTDglf+6
6DEPvXJZpPIMR8w/EjF9fKse81FYQoZzkdlT+xv8Ac9ZxcnodxiUoOy8zbY0dWWeBhJ0G6rJscqd
1WUs6hjrt0+iVlR2BOG2A4RpfQSV4Xu4oFvG15NK9RIEUWAJyR/mhL3f/3dObMiHYumDJiavzN3t
QMcUUq8kzssozr7/KO6+3qTVjdc+fgXBUtlqmqt3Uq2/mkYrs3l4RnIUPcXqtKPyYgjzybkLW5i0
ZP7purRYsdE3ef5FzjsjnMsdVf6XMQkup1v+subq9urYs8mJiC/yRXexpfNEtElE43vl1RF9Xe9b
swf9vB9N4yJtHfV2O79iyfdNPuaLl+Fq7xkiBssMrJkZqN6mWyXNMxEt9QOGUnFMjt/kjk+fm3JH
XyX6xiVQ7jilyAzqVUxcxfiDnI6V+qonvGFee77OBF+H60LEUQVKxQKpOgIhqhczFmnKe15Js3g3
FaTj2lh2bTV8Xx8AxgOd7e6USR+I9cZjJS8enWxv5CNN3Dpt7Whekxplw8XuInRS7jqEGCsjC6PW
U2HYtX+UH+pSDZnU1ZUhsJI3d0onp3udZUKXjgowvFXKCS+7PNytpDNs5ZA5SNsHTNlXc3bPTzj2
r+z+Dy8MK3k/XmfOfcIfwNSbLz1GVQKn2N6N2CI5DmApx8ihQG/WH0Ck0Wrpir9iRxWNGfUw6oXJ
uD0PPcOhGHSXbUCrBuYcxeU8Ju1muoWgCzIho2sQJZLFVy5t7x4GgNqXYAQ3vNHuOgBTAFQRqXuP
PWaM0jDBz31dZprGlqseToEmg+DtU/Oi/51n7GHh65MvxT6aJB2YnPU9muVhuq3m938kHcGg1viP
jewNmyObhL8ASSEd5pkqOvzUsc5Hl1WXqLIK0ExRKZHxrtouFvMap3wkfCa9PxUBD8g5BJOtVjt5
kTMeOJooOAO+VBD9z8gY/C6u+1uvoANykQi6qkeeilwuPJpVfD+X2WcT8Tql1DUcuAz5U29cI/wT
Dzt+ChY2WlWRoXXXtluL9TstYiecqMZ1wURV+QgAFO+anqhbVEt8jHzIFXV/56OTu3QfjeOXcuQS
Pksyy9BPlCTsMwmmAptfsNE3wbLQYF4LAYR1FTQz94qZRHxbk5CqJO8uHZeSM19gyKUVOsMoSiaY
WUKH4Fd3ltJs+u4STA9pAM8/GgoiqTsOk/HwbhlhhwVLnVWbWgE4W9JLikE9raAokQLeqyvqTx5c
TyaQJB2lWdpeYNWCF0ED3cGTwGU71fQppplvURZa7yPWCST64JfcSRk1SCWlgiT2eoatjUSp6zt9
oPmyG0jyx8fnIjbTgTUnqIPx33rLxRQFirjvUCkP4GKKNx6ut5HohNaUjVsB5lHFAXJjvIF4LpQ8
0QERZPosYIXDdJeo7Lr8j6peFB+Uu0yyJQloIUs+bFwEllgeW+xoPO6m0cxTP0wFkeBI6UBL/87K
hRzb9MtVFChAU+IfCSNlERz4NNfnzHrmNGVD7+TWNL/2wYpkxcKRbpkPYbNVLePjgSaa3taBbYLa
WjWi12h2ce0VN0uASDBy+TrrA8iChe5MKPm3bnJIWKWx0F3v5Rbr3vz2IBzgt1KTglRAO5w4sWje
rks/h9pea4ZRyVzMNrmMRlrtpM1aCQjoXoGYwpoKc3GZATtAQir5Vwr0GAoplIImpv2jBhQMRyH0
A3jRWUEN7QqGeYRlG/TLgVHDA6f5We/Ls0DNqg9Rwe9ALRa8psi9S4mGwPYNTnbNQQ4PwKtVkwmv
Deg77UrxNVR46paOYSbrwqTvDln3k/CUw12P0kVgviBGhZ+0+2SLbAZx3Eq5oOHMnR97pjJtpX//
RsnT8vQHlPUu3um9zZxWc5JhZcC0/d7nkSZIMA8hhol6trJhIKY/vIw623bWRzda4PN2DB/u1zok
FQuhVOBRUoDLCY7ddCzb5IB01lrxXBNUo3m5vVZz+IvDNiQqvyM61LeJxy44HM6nuFyFGlHYWNMe
lnSTrF0nuPDrfrp/DbD7JBtDqeNkyOAh9Wj/1y1D/uFbU/bglxbFw0yYPqwoa8HQjHL/7VuNITvA
hwBZEdPQfdb1BZR9wGov+nC9wlrnzZv7G/slP7B4ZQKGwb2BrkdL39qeAFZIwo7QnywiewWe/KPa
oX6u8BJQv8El/iqmtfLxmu5BiIdUlRiOIHPZsYsEHp2TIkBBaOyXTz1hvHs39dWurOv5QkhL0FWm
zMlUwfAD5dLdLux9um+ozpHrfGWY/We0Yl6daGWcI3nGutwjH2sbTcYX0stw5cGuoSw8hzOmRobg
YxDULBo8Jwvx8EneADK5KgExxnGvWFTX2bRvLZrpUJoSqfTDNSVkZuMDhDOluEORYQNIWGoDajjs
1698Lgy2pLWg381KDpcv1wmSbZzAVoYiRDQ2P5aIsthjuUm8aOKdVRTDg/xAPPjwpazTAAMoN9B9
Xb4lLsdwrN1Qdw9lOZuXHwmdonKLXlxKHquALjfN6daGtuiRqm7XtGXwM6r46sv/3wA0hLLJByhO
dWU4BhPDwHxhjC/a5vfmn2w5HMPqznv3M57RHcZy14l/8tpb8b9DozvpbDA+w9PKwAz6vYfTKJUh
GFiwZQ2cXAgcWXVQiQ8HBLPJpuKeZJx9UYGZmR0tRsCG92tbi5rSjgY4LPkWczxIbCrBPcBjUZZR
zHVqiIK6VUuhhQFGwQeDXmRgKG0IROxepNMVNeidtn/1rWH6SPCGDFOsF3p7nAeGd73SbaGk+hTh
M3oFOJ3kfDWQwFVaJf8nSvbvsWYSyY06ry21tB/cfCP2jSnNtGFYjv3uvNQy7A7HuwHcwG/e0e2d
53WjVARurxgapF/hJg3urLvUU7M8wjihn44sOEa9+NfUxV+2QL1l8gbWLQ+smhBNGmYXe62A4gAJ
lOghVqVjPo63nprB9v9rR3uQSjY76xwtpQPy+E98o3D8FWaf3/yryOuiHT5+DY1NzJtyOtCddeE3
mGSxpfm+g3UueWs94njrtmVbzOu4f6p5ID2W3hIU+x1vmd3TsGfAGFbopp88I+cWLPbtbn76C7vx
TvmYMpzXWMJGLN8X4ARGFV0ekeVl3993RTSpG9K6Og4NG9zn+H+Tdad0OzkuL7+gkGN1UNOW8Huf
EyAI/VU84KMC1cOu4wOL33sEEzCV3Bh94hWK2GfFVLEV1IOhb/U2DsA0j2gjlXD/AMbgAPp+YtJQ
QlJFj9YR31d+5HRIa+g7Akk7YMusVSIRiP+5mbo+y3/D5J35mfU/DlLhdF2/muBztSxP5tzr2+dP
QMBap/DLdmfF4bA8Ga3W5TwVAtKoG7D/sSbtmLpa+VACa0gMSndcyMgU9glFuYOPq1g7vAyVWLe/
UiZ5L29EHAMOq0hTCI+V8zP9xdgATVhdddvIwCa//0BK0wgUkKf8afi59+3QNP0D2pJClbVV2stj
OEX4DWIxNzZRgkHXozrlT1xiJL2K5zZF3LesyjeDPJe/sbRqAz/KcMEqamIlHah6/iwpD4TDl9Vy
HNqEg/zRa8B9fpS1kXdwYGwDjIafoLPUb5WRlHko7nSyg73lgvFM7dLmsPFUIcQA1WF508Kp6hPV
e771MUaCoXOP+2eOTyRjfA22n349vMoH9uXCYLUibj8N0F0MSRCD7vb3ONPsDjQjPk/DT7UZ9K53
fIcL6m9QI7a+RjOEZQQbUFWhJrrJk2nk0pL8aL8QVOsVk+/LR/CLwEcqImJkuOFFPKrMW4vcbNyL
U9g6sOYwHLZ0kpmoCk/+0aSIEmyH1rDVjoYvWpvOqyqnCEfxZUJ3tC+FlhUUpF9H98UHu91ptMh2
03x4OcFZofIdi3z5E9Cwxg2uCPy5cg3FgGWa2rE5H2Tbmhq+OKJpEykl9wEJNGVfjbIlzi0S/AI9
wa73JD6OcMrExqYHB3zT6TXGkPQh5OkzLDC+xAXbDm1ail83JizOc+jF63VterF9AlfOuz4MkSHp
ec4cyI/LhKaxfX34Pl6hKWLlQO0nW4MW3aD7OXC39eQIu0WuYQjKRk6mPR5hqrHjloF39h1p+89F
Mya3ZqHVVdQNPP3gILEJUzO1fntObk+D8+cHecQS6yUTt2Liu5THYyRNNhoRsqZoOocg1YiTfsUL
dSPCCiIzjaB3hWlpFk6sX/DXAwae7ihRB2OnSo7PLiVZji1eMpYnAG28qHgnKoDoRZN0Xi6oQXYi
gvrjaZt0U+AtbkPnjXpNYSNc28X5N326VcDsC+moaHO8JfEQMXS2vaooro4Xi9ubqWy6LDzgfu9X
3hNE7hXqVcAfxL5+TK8GEs91nx7TzKI89DzJXteE1ongQ7vVcBZBq3tEYW1mmp9j5TAfp9BHggrQ
jAbO6wZr7LR3VO/7cic7dJCQrP0zsjlU0TyRa+CVBqCA36L7DHBB04RK6ZlF5hW0x9pVInuTJq+h
PIrgWChF8wWXEHC0CVcwryt0H8BloHssaFqGRAX1u5JIil/tHjaF/0WRX9v/U/uCckpi9Su1RqAl
/uCRIbB4lGqrJThCv9GnqE94eG50whECaxVT8ona7DpeF5zmx0u0CynfA/cjjBcfp/reLmA7nTJ+
NlJDvECxBLyvZecB8hRvo6bl4knCeEvlUDqNv4QOiHWy2Gqh08IL4HiSYaXm0sp3ux95qk9sMWek
oufHzckz0Hf2HfAH/m4Cwge3G/fdJwvuCZcNs4i8yqq/68VtgCzmfnlYno+jGU+2t6Xlbe2cb1l3
zAnQPH2l8OQgbp/sP/3z0OzAm2Rl7gGOeHoGCtkERgl6IR9CHYrP/1+4l1vXg0KZelmUWKCThp9d
ROd/BzLc9RqmoOBMWO8O9hCiCL+Juj6iqA5IRE1irKdsR7q8cU3IdM3qNXmuehkkUZ5cnUxJPvC9
lEELs9p6axuMnkHPAjz20ICFOpIQIOblGIKspNIBOMW3dpDj5ewR/xZsPDTEK4AMdh5iORLkmEDg
NzTIX6i5Eok3jbaflQYANyHnAM2KxCaQ24hrHPg6BGh9Z7q0Lri3G1QEhVaF8cYFwD5auk84awxf
hAfQrvPz8qZzLQ+f++GIiHrRL5gZjqpVSxmWLPn6sCNeoBXAb9u6G0cJ1PRCkb9MkyVDZJiCw3yY
EuOYDPwrlB8oVbIMwQJbFyS3a/emcpZ56GsBMQP7a5B4vdqk/kbTxFv2qUrmphvHtQFQ3FKOXFVU
k5fIxjW2QzljG8WYRgx1b8UGZCUUMoYALcNaN8Pi5QNu4RLGpOITirtIYR2XiS8S5pfm9QPYyj13
Dy3LECl5TrYKZ0ZCgSQMbgBqiAzqC724yiF2xHwCaiemV2TPPmYkJlpVaUJOznNaj+OACdIcVq5e
uXuNel+X7vfSNOWH+rbxXdNjdmW4OtA5JpGNohUndeYD2+iRsl3E0xyZWCL/mi/04i5d48tmGjya
NSlOhwt6WP/p24dXB0SWlJSsKQs/KnWu4HmKPeSI8MCFnN9bGdlOCE4C/OUbbn43JzhQ0Co0VPoO
x1N5uwTYpo78/gjgssNoq1ud0ZL7ZqqG8c9QxKwG2XhihIGF+wvy1P+wncXTytVQDaJUBwQ39SXV
8vFHV7TMvUiclSU5Ocjt/X+dp/TFGh5LZ0uD5gl574FuEuiVKv32fw5hcHLZODhZwQNsiIUfPmWI
tFG4BvuLKTVgZlAh8Nnv0wOoP6f6IzEzgrlV7FlDI7rBxu6IRB2aEt7hu31nRIsAje/w7BkonCP3
Tc0aRbZ4/RX5H3lVi6RCI62NdWdA2VzD0hnAgg8HHC+28uPx6W/R5Q8gbJK340rkVOUg0ONEkpng
LyRAxUr/EK3iy6d+LDQW1lFnoQiz2resJvI9Grgatb5oQXVDShJZLXsjPKr1hLoojIKH6LvwkuM6
/gzxSE0RYqo5Bvxc8G4KC/NRRdzuIjhFTi5MsEZP/cuS+fHRjb454472HdMw9Lu4D3I/2zRdh8LY
RiGLTQXc4TP54HZ9c+PcCESl28y3nzgUTvUmKoTub6GkcwiXf2/do5G6ybVHMihymIHIHBzrxFfM
JPKbm/peeLfDnpGTlOwd3AX6lmLaREsXEb8bSG2T0un/4dWSMexSTvtWldWulJPsIomkOFi6/yHd
MOd5Ohl4Df1n3muZ744oA0/MJcTeWZJiGkPMjaAFTN5vftORAOiVm0eq+72B3g7QQCRbxLsqtNb5
oL7ac1C5aqZJmvVG8iZbkkTc/CTVmMUi5Yi41i2akgGy4UpQUOzK0lMbDpziFVBI0ehBNmttftue
4Srfm/TeVHIKqTqIMhra+2baVFlrXUfnXPxMo+JASoqGpwjzQjeZ63kOOMWXZs+2BR+8YVxgvfFI
X/SQOd/rPHJARe/r+SHOSFTKiJ/3te7UVePjSfKtXfqORN/0mco9JI64q0s5vv0B4PGG1eM6N0aD
0/V3nlm5SkYlae8CXKhBvH6TGZyrtCOIThUmb9pMLgYeTHcvLdIMA+JR6ecM8jD1FAll2QroVyEO
dj2OpL/jQBOQ8UFIEqsPcvmxjkwjX2hrB/ikzVaOSF9HQCOe/0X8er5QhZLvh0tsYl3oyQhwgSu7
gcncmhO1UxD8hsHzgt4fr0anzu/5GIcPIm9Hb+LhUpReUMDLaP8uqv35N5HNWp2LiAA9cMGUNy4/
T+Vvj2XGIUd7C9/OgTuWdfLIBwRmuMSxdHD6qTrihviWeAmPTR1XMh9yaEXCriQO6MPYfSx6V+NN
erzczXBxjfgMQbv0dpLcGq6QSJlaP50Nm4cCElMYYyV2JBT2qnWbUR91GYEBadXZZ+cCA+IB1xiL
uZ9WTKmNOwoYapTzUg8WpN4hqc/ymREHlaLRhCogPlDACXLTqHQFcdzFpBxHSUbD2WHU4IlyARbm
uDCZ4yiWI1+uraOUVuKpYrKdbayOn9Whc5tsZqipp+hcSZoiHDuuT4QqqOtXTUeJ6LrGCLbHAiAz
Iz6vJgNHO6hY7OpIy4xhAJAl0/LTFRhEQmC+QICAsFPekfF0FBae57YYFbHM0uOkLn+4oBxEIS6n
7Fu97aOfop4LMqqCAUqWMqoG+4gy45rIs0fLVx5qn2srNAVDQ9l8lKAUtWI8oW+7AokmNpWle2Fn
cwdNsRqhtBxeIJmNCNfRTQw3nccV2NSzpUh62qd6kiqLhWmGJNkwJ84zKeu5xs6GoqJljihBRflZ
vOmn4C9mUd3eIIER8ZabbMm0Wh0xSBS/WVZu+XD1hPHgZumNjUQEHszSYtXFgiTYwQGetkOIzvVh
6V5ZA85InANVary9qXeUYJSfBAJ314vglH27+dNs3JuaKk6ScJKDt9l8WaPXrNhKCqOoBWjoU4RU
oszZhV75gySSZi4b5O6Pmrye6K43uuU7sSMd8yIAhl41x84qK4yAEVv1ThJxYxCm2T399bDzSN3U
r2LGuXQqKfU0q1voBEaN1lGwCUj2xlWltDRSf8bjQLlu609eV49MfW63p8g0L5eGSDI6yagqs4Us
BToFuNE7V3WXEl2Gryp7qxPABjx58o4zP7tnwa4ekaqT0Zf7o7kzA4CJNkgYnDv2GHZeiITawgb0
MHcnbnGPr6+tAtrdIdF0zAWlK1kPe7njlcUjL9nfBdRyd8QWFYJdlYIgO4r6SOaBkx4fjJsWsR39
9ermdNDjxJMKyyuu4a7FsX8g5HroBcSmpP46knax9oWGfn+Y6XgohZ2NwUDRpgB+c9JTPvfnlmUx
VBYys3cEW7K3XZPuEFKapjD6n04evTi6m7fC7aCJh9Fz68v3IXaFQOsY2XKoOAMCZy/g2RyrCH51
bTZ2OS1bElGUrOivw09al7CBV4TopTxTd9/m/KvMHBE4vKC8VY7KZkT77Mwfj1UsPCK+U1/md0mL
BMgR7cKXJqste5ssZ6z+e8rTyjqJxEv7i3YJzWiDCoO3bY8PLheL3LTleX9uaJXmyUNPimvoMulb
OcNI86Zcw1rOwYX4TGT03f7MzpGPAu5a7tZl2NP3VzFTAiB/deRuP7W39wCwJKr2kUh4iYbS40ab
LAf4esKaxlUHUg3nONrfK3Qnv3yH4SRD+FkTPC/GDHID7wzwXAo/Xh1tfjxJTigAWQKaLwCmDgIr
aWicU3yjrifr8395u5pl6cYWCLKdARH5XjG1e3teizyOuKQQBAGl9Kbf8fAZSMncVmI53d7MvOzS
nYRkkyWvvb279QeaAT68IW0gmGhEPrycRo9TDuiJiWhT7MljbSWfK/IhDRHaGk3O7lUvzhb/4TLM
zHvvY3J9qU/JIC/ZkPK/zU8mhVafkVOJqPhqt+NGHrIzh5jBqfwrQ9enzLMl+f8dIlhqb4msF6eF
4Bn9qOR9ouldI6SriXtlOaK9h8ihCFT55wEomuyzW6Nj7rRP+zpRt9LcSbuSFeweP4WuROjFNmbv
LJLpwbhMbwnfTawxmQn+h0CLYUhN6hqAzN0nKu06y2LrcMDrS8w2hTl2u8kJA0IbqPPXg6qXbFds
e43BKS35NHNdFGH8opkC9m2YTva5GVAqBlaDJhwWZGGWNI/iWDsCvV596XftFKTMU5VEXG2kugl9
7r0a3/ssnnxmruVRqVnf6Ymza+SRBsIzVVZzjjsMBPDJYJ5FEXBOFGirJrfHbTDK9Q6uNcCIiheM
mNu+CUOxc7KZrWwPnLTx5rZQn8cAQZ559wUIdzcnjwoO6FRIfnWDkX7ESSegFD/tTuFJ5lQyVWm+
xy4CA29aRgETCs1pP7rprfBHV34wSeiasoZuAhuc/vBg7xnxS8SnlL0fEJAqAbxYPrfLc4tIhTrT
Z54muLw3+OyQuvnJJlePw258RjsZ474v4PqAgeA9rjCuu1guRvOEW6KQqYgcLGpWnfjMIvIvoqe2
wK/+RIqt4sxZhZOVKLezcYdu+hod75s441ARLHSX+zIEdZO5mRWkW6fu+HGD8/sNvsM7vFSBNIzM
Z1gsLiMlAYShHhLWOr0X63QDw6p1VLwtRyWtHrqdpol+OOyQu+GylYB0WwDObawDFXymRlraf3pi
EWJRNcUEryp/7MDRJrdWGHxzupN1Q0H+Sl2qp9+2Rxya9eDHkFOumK+IurTEwAOrpwlaE1Aa6NXA
kkUE8EG/qYh+bBPXuQfEMe4MRVtdHlodeKKj5XGVs395MmKB4pfVlFjm5cAM8f5/zmOwYaIUHtvV
WPx+jMpShBytU/waCT8HWFWjd6hehoqCKdkZq2uKg7Qy3RcG5ip/jy4gozZexvhhkvDfJ2AWAZZH
ASqNyq1CpRwV8oGgLPmvqktpbZbQf7Hq2ipAqWKGcQHvK/UXrDRuLwXlC7chQ9/vyBuymfP55Gd8
jUcEfTQ=
`protect end_protected

