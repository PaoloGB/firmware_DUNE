

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
sQ9+7UcnCl0zgHeRYHA8r5bwMZLo4n9NZkOhFz/txxF9wvEgtq145kQQS4uZnO/qxvCA9MewS5pT
27ngyZK2GcOgqQdNIWHdiB0IL9Ko24C+i5e+wVLXaUk+SoaJT3eAeNL74bbQbNY3bzdK7QXDXMr3
zIE3MqWRHBY2DBt8lXECaGfZxnmIlua+lpQecfSQ7Fnc3C3gcMuqv6PBlkv2Fykbm93nOIaaUwf6
dRwMaIwW4zcoJ+tTGrJbc5LslpkH1qVEax5IAqa+syjYLLYmt6nN7Xl4bIUarU9tW6ed7mbx53FO
A6DFMWplD8SmPDECMXggYMlKRWoEGm6bSy3ipsi2QrgKFIPdNk2zCX+0a2YgzdJtJSW1iXJtoYfJ
8yJBB1RD7I19aSTzhdpBKuu9A4DF1v1fm5dRjpnsBLXrFuDhxVyITSGYPv2ttB69+OB8WWhuVFJf
12r0YBDFtsMVGFnsSln997zlFgSOFCW6RPElxUE4hiGd7n2Jjkfqee+jdkdbZypmqKYJLZFfs61P
IlpAmfj/+zvfDXYqk/bQgU/qY9WQtcuPIULICXYY8t5w8TzS5zM/vInSDJL6mEHsu8ncJQzaqcDl
OIhIHU16tD3jn6sQQnwTlCOGETiNVgO1oHKE7a5TnPFtJnYs6YkJqPH0vzaU00vJs+JA5KnhSn5G
qHRXOiR+vP5FHHphkikzSppHUys1r+8orlz9PL6I5WzxKLI4+fxEWAj8nZDqGaCEiLIBDOXLsxSV
/Ya9JiM7ACIbQN3Jd6MY3Miz9Ge4DvpvoJ6OZe3jHbG1yweG5afrzpASxS7LQJLXLYKJVT8jClmP
ICkdbqTWZ1AIVQDDJh/qT3ar0V5zdUhdrlzLaBDd2ascS10sTYt2S0bdPtMccb0CdqcwOJeBKETS
S1XUqtb1bWwSacKKaKD8VoaMdB/JkGPLrNbJQZApVIgAec0COf+g7xJ9Yn8HCtogNZ4IVLvgEUe8
jWlxlAK8o/5aGyl22FyNiZ4B6pRAN69cdFoTP0oIbpV6uugBHmf6VFkYd+doEd0NM61thxb9LUjh
CsqOZFBhS74uTRzLbwmadwcH7CKIZIxGhMGiuqYMMEt7FcoD9Fl+UvBu2fl+9m31CcvZkc44k5ty
1SA3JRK9YeWmI5HpYC/i3tGISaB5fPr9pAgKdnXPTuY36C8EZ3xlbA3bhzfpm4vWIzNUDnMzg/2P
+yPwGHUq5l4frBfH51Gw4jyKlpRejBzoR8OW3pQDkk607Psl3WYk1L83eqoYJ5hJqQlS2IOrKrjK
ISbwMR/2GssRPEFxEaRyqNPjEiXjQ8bfWYXNQf/Hh1vfcwUuQUkswdWjWME462kgY0AlDgodR/Uq
S905m3hyNPQfSenbFCOAs6C/KmkB4ld59ckjfYZtK9pE0pWrSZtrUN/snP76ifJXKjOyDPOQcWGY
r2WiMsNGTnTua1pHYWAKdyuPD0nJLiywvpdrm6Go9akgyatMs62+Pn/dIIb1CY/Fx9iCUY4fBu2u
vrroyes5pKBYVG7n+mAOFTU+jK0B4ek+2QtSj9xmQTSpy9ZIcEPnnQR62soL5zV3g0qam2gTin/E
FL+LBnnQfpTTS6Uq1Rmb8th/Fnewdxu+wYJa4W7kktPWHMrfHTb2o1a3KsvPmxXU5x94S/u8zP9x
NrZZ2VUzZlUGuvnI1oVyimH5uXaoW3UxK+Th2pUBuk3XLM1cosAQMX1VydaPtaFPZRxykvCZAAWI
Df1Kju7sEGbV1JNfxb6MRZX3H7xk7cg1Z2rUQd8h/JZaRs+WnEmNnXxdm13S2Vk6DPAWmi976irY
ioRy8dHYC/+hd3PCSi6CQVuQBpHfXx0V1S5PMzxvwKSICDr4TR/1c/eCDntvJkqv2Te8JYBCgkuo
zUbKRsPAUUTLXPvemgYTQgkzSB1kqashK8iusBWJ3ECNPb1mUwhZGjkxOs1qU8GN7QWNvNAqTIjq
LEBf915NaLfL69G7PLgqkL+6N++4ryQWefKCRtl3wAA8xImGCSMgcYSIqMszmeWISWQQZLgSUTIJ
bFFzLIvVPRWF/pCjcwG1knzZybvW3bI+Z9kG6wpyxUd9HrZWgITm7xndtyFd+VOQJ7rLUGhCTF7a
C+ZwcpocRYjG++5CyY4Q1v5dV+Br17aejGkw+iq1EhtQrBZzWaSo893G5cSRsoWI2YuEAal9ggdQ
OwItkjklOlhhmiaCvpa1ETrZbOmWgnOijw5lrwg60wxQhlQRtaXKm3LFvWajxNU41NWxQdIrMTac
etI0syOQIqAO2FzFLWC/0GK0P9wDR/8Ms6Di1UJmtJyqix/mFtLTeAqsuz+oXeki0AA/N7yRj8Ge
I8o5OQzylZtPe+Hsh2j5fd4dziUKWj1kqQEJSvMWyseqQC3Bt3f/V4mvSGM+eMRCskZ/Q8v1bisJ
i+rh61WA46ApEr/jz6p4tE6C5pJnE71NsShmEL8watnffvJ6WD/gakvh4kT6jYev1IdoBhMn8P9V
ENrPrZqr221S8HekCziGrWAlSoR2Jq+KxBMyR8Jvft3RSueQM2ECgZneKeNJA5UbiUjlo4g2YAcK
ZRkE5wCuxZ0ulXEgktZng9rAi/XY+C6qe73XVRJfRGcMhjenpO0ZcTbrtri43UYP8T7R0DTchboW
H1HFykS+FGm+XIhwcvLf5TqCqbFNtoZxzuiBPZDDGiZFN9RCVO1xemMTvq+y/PDKncM15AREP9a1
A5HWYrQA7lFk4PVEldyXLggnN7YrbCeUGnte0QF043E4Kjt1yn7la0SwzT3f2hW7AS4/2k/BXxHq
J59Eei+IrKQFK1tZ50DHVDcafdPAoMCk8oVJh4LJvG6XQRKiHaZuccJbicoNV2LBcC/t/VOQxi97
u1Jm93HZHUuuiqQHwCCeIvYxuPkApypPQbz5MzQa8rMSgJDcYRbiqC8KfAWL0T4ab8ntS3wzlQ+c
SvAv2vlemRqeycAO82KlkbT+JnlWzHYIVhzGVs9c+6WxYmVV8uHhS9f2sF+dabVuVPmv6S/6TC2L
ziF1DHdkXJjOF1/m8caahtwYioQAGBGKXvF1+M1KmYUd8LhIxYfd5/G3Its9048tDAab80urxZqm
oOVbsw9wUoXuqBdxhLCd4e4gl51HUN2+SW7aXsKlXgGJQ4MIdV5mSysshPOJl+EA9fY8z/tmbgfS
LFZ4Cpj+4dVUT4FdvQWrPK3iIwf3InnFqF4gsMNeYriElPHsBIGFCZTXk3T16Ig4SVOBaJRYsASn
i+5bn+REdVguhoSkWzQfAmdCrowZhMd4YCIXvAS0ZXlxIFCNJnbWMODXJ2noMOVUvgmOix+rgVf0
V9n9mjroIPrEUo3Q8eDR/bCEImEKr8DO5zhBpGMnTkdKZg58jl2cLT8k1bGI+26uk/JYYZHyoeOG
ZABn2F1+zp3GyrP+J4K2IhqdITlypa2aYA2hcRHDOpm4mratwnYi4d4EXI9ZdetN65pcRSekHTZL
cV4NseBETZ755X7FFoc7NR1FGEDKyHWOufXof4aDP9RIx6TqULv6Zzt/ejwCazvnYKjLCcTxclVw
hMOOdVZRkCJXESVbUbPUZifZr1BJtPw2sdU4VgevsAbPFcakMjTnK1LDyuFv4hrOx6zv3E/0bTT+
gVDcXad5j6kjLSYI+ZSMGR2UFy5NIGvRQpqSFLpBhLnPhY/PZet/YiE6CQ56uV52apQ0eY5LmSOt
et3hQNx42nXAdriUaw3NTPcjYD83ImCK8eGiREi9DkPpCfMzbU0dCKLH8vDs6sq53T7DtwvQNfjx
LURnNiXmr7G4FAQQceFyDAZrI/8Q7wMbHOQTTUXqZDZGe+qjZ0qG7xoh1x5XvRagb4rwfTf7c2f5
QHH8ycX7hHVPDRWWJn1FEsM+F1mbQmjULjaIJoD2D30coQo2uM0qMBil3MxWyM6mdOhYRDZMLBmg
pIFiMIhKppsiIMATKkElF+67+/rqmCnavb24l+TSpTDux3ZhR2JfSe+6Fd57fKWDpAzKznABCumO
6hKBx1Bt2yfommcv6PPd0b4dTzpOmSuMLBPzFMi4JyOU5ZDaCFELBQ7Xn5tYYgGV/9SO0JBu8TZp
BYnqoqq7IVx9UPuIDeTZtzslcuHEdg/RyE4unB50WlxDXI7bnYdQ61q79SCGhDrcbxhvWr9D7t3k
g6KjFVdx0A1ilBi4p16Hyp8edR8klP8KBTEILjHgxBMWaS3oLC4YfmIISCE/PiBoLMNxHiuZT2lv
0+myJYx/qBFktQfISJeWnXtynGj9xevGrzJloXWJ0iC5Z9lAYxXsJoFzuRkpFxVIYY3wVXeSVqHZ
3jF2eEs370AAKwi0y1MtoJhDiWMhbpfMD7JNTvwAOGUzwf8DrcHaLdXKRAkemrUtnE27ns8eYf9p
+fHgIRzprKRD2T2Alkb+WnAB1diR6da/+z1Jv1kjCnbfxZOSOD+AWHg6y3tjI55e0aWioOKi0mGr
Iccn38iGy/NY+QIMxFn090xue5sydDhqyH4GrlW8awemjB+Sp3if9ipQH9hlfK+P4PD2uoTKCw0X
zFJWyCYq53CRnsd5ADZMJ1UXWGA7eEjHVtHzn2V9t/1eYdEheAPoueRSXpm43beFZzyzYiPeZJba
qLwyrGJuGfHft7ttCBYpfEK2dRttq0S/Cplz8YlriP7pbOfMapsAklZahYLz3NgVX4MI0IXMxRAt
j94VAfuM3npMp9SJmpI648gW01WjhcNw5QiLd7+bkx1WPNFo5mmWrHfAWnD9UlfvDlsNAeV8kVFk
UferfuSF6gwoA6JGI0rhUsFqyFiBIeaHGYhQ4ra9uobib4SsDASXEC4wif3ew4TBeE3uydmt3tWo
JwCEGfvOp5TB4MCZ7WajBidISW9FuzILXTylsy8M65Bmdu7dWm4i9wnGPtl48WSs/jnIPxD3jNGh
JH7uURPYgr8CoMfrAeBKf4bSN68eLlMUi/wvpqRAZB6U6kRlMEVWA9ZqvOERr9T3lIkSmr56aOAS
Qn4uEqJC3mFdKoilTNRfijXN/kHwM+nGVv3k/WgvCTZIKJo1kBpDcPIHJzrFVRlHnxNZwYADzHkX
wsfXQMRiXUV5Z32HxKDXNo6tJIItcsRBt2asYUeH/e8EvqDWif9lXUM3BrAhcVpRY3Hsd4BE/e5C
IHjfpr8Ovqi6CcA/wWz/UlvzYoa4imTpEvjKj4lYQgJTBb7gj2LWi/q4vZI1rhuH21i1hxcXITWQ
RorJ+IVbrZNI3h3vMQ8XDb5RiPHGZfR1wt+5Xfwzac9mlsbTFfum3LVCEQzfLLj/1Cqw3qTATs1o
15raObRBILbHK46Yv+5oUzA3RWjgmRaji7737sFyYS0+SlGlWG2xoipY/Oj9ywhwNwsDlJqijCpy
8etx/VDnVEMhydv0WRXWyfiLjUmJZty2xJPQuwxdu5x0qTDPWrlohChfRz1bmF5UZFN3E30Ui1oC
iBpbSaBrBKraXtqHUdDj3ca0tBhdLrvNAb+nWcq0njVGb6NI1arEexg14+wbnScP+mGstasT5j9F
88/p5J2K2E/hpuVbhg/N/jBfaqwPs4wlhghPzugOo4vPk3V/RRUPQabs8n9NmOCp2bw5OskGk5Zq
3fVBYvDulr1JYWjoDUUE8IJacmpaEeTyOMZ8xlPwmXVO4abFPn52pZ0fUjUyLqoVu+Qb4ZYI3a3X
1pHv05e9kw1cdT8d3uiSwP8DNUOpOEBrrW09wjYxTcNL4VAy+U8y8ktIw8aiRG2V2U5wBOKRrKY/
349nGVCagI2BoV31zAfcUnAeoNeO0mGUJ6u7Emla30xQrcZ3ptwmDQmPWZa1mXv9Av6mAkV3rdQo
tfwHALaVe0m8Q+Bm/C3lsTqCSxJWTr+62+BKq3WPcAxpFd71BD2TpQGEsvahkIek0ddxLxD66aZR
VKEwUVOTbtA72pgojLTkc5KEaSID1yj3tkZ014/kIRbgRaqtf/MKoTuSPcg6CCNTgoxJ6+uMxiSi
0HrjBUr7jYNszPIr9LUqtub4694UbSK8ndge0QlUypu7ky9FgX+0+FauJcApGSWpIyP+uwiYhaYX
b84J6BkY+mzD392sQh/S24bUrIbCNHFe2KtfSAjLBwnAkHmHJEKjpF7+VJ94evRHohj6OSVf7g38
K8PvU6YzLQPfjRMLSxgQs2tg0pwM6h3ZAghoaw6kch18Na5bdq2wFotWQtsP8xW7iqA0HRGEpGXn
4yByfCndvJiF8wunGREjC/oanVilIVmzsis3dpKKVqtxeOJWMePlafUGkQkGqOxYPeCnuhfwTQtw
AD6V8Nyvxv9dGixu7HI6Q6QMilH+vGXmdmAqnMp/ytLn5uIWnn0WGd1DoQRvDYnQkGh9Y6Z85Ybh
rDqNTKcLHnAY1vbuoQur/CcsMQkpANcEEnLfMMeWs27oXsQI0AUJNMyoD+bBGNi99tyfS6kPytq2
CrEnXOuQu8c+M9QGs6sz40eoU2zM5ALsJjwJ2z+WspKYRGoxT5X2sU8E6k9Sowrsi9URGPOvDH2a
lykE72rSvaNRMZ4TKjQy0jDF9DSMhNEdER6pRRNg8ztpAi8NNNHiKgmQzH51rAtCNezxUPJkNfMd
+nf8VbDhRPKFzj2GiAZQaf7324GWGXvJHdO9aqOWbgJYTSmDXBiR4LylsvE9M9/5byfq7VTcmCnL
4jmPxUOANqLBvdTMVAkRTGtD5Nh5xLbQAzBgvhxAVBFX6kcUt8aUkIHVz58Wutwmg8sIzaZUcEkl
ytdPfUpQL3ZtGje4ngku3TTxRXg/HYuz5TJbQPIROJZo2De6KI4UIUIkHDwCw64tUg13yY8ayZu7
yjtCkCPvIWQsfiIryQzLPU40bI3ZVmhkTcgYmCfVagOAcTl+IrzWKqVR1kdaTx/KwjvOP35ntCTH
Px66M/Y54rk3WThxqBHPeju77PGx5v5UX/8MXFXXCPPn1pjtqYUfR6LDM59w4BzzS1BjzwYvPB7X
QMi2LzoYz16Yo+TJpilzibwzj3jOJUVD3V9bilFpi/8fZyeMB5NJjfmv3E0ivYmDSb+5Y/1/FzI7
TS8f/nnIgy/0WcAnziUSgp1/1VQHWcIKlHftqg6dkTJJuyQxQjQGKDzhJWOU6XwtYIHPPqtR87ME
BfIzM/7I/RnBvb6JmFsNd0hUw0H88w/Ew8uBDR/G7BJGU7fmET0/PsldpRqr3qa4lJZPy6l3eB5L
lKoowUNyKXKsR4Xs2IKRpv7Tp80Z21TOvKjJzc6nrbyl24S67K/eIanXj8ZWZAsnO7ewdzyzpzaO
9PCYSKufafEcriz94IlI9MlWvVda/qQ2P7H4MwkEqSjvrvxPAqNXKff1Xv7pC5Lem4cLCPpYQ1YM
KzV/mbLuwvffPs1N+MrGZm4m4u1YMbgGqQowSKoWAgjdiXv318GXgefTqa3EvCOf/6M8SVfNw/fd
IfjvXf6r6uihr2YunAC+9FfBYUjW6XQJyb6v/ko/GqPypTwI4HEx3LV71rDAsVq0WsE+xu8TDR1x
d+UZfjOe6TiraMlxCvtjz8byG1Q6/jTcmp/tSfxUgm+vltdKqw9I5+JYSorSpTnOZxoDi5c0Pa4s
OL5HsIJppDSZbgU7vTk5cUrqlK9698/klYzytpienD9HMuKLBadhKrwyBmM7mkGGZF4wYdrASKDk
q32WEUnVYoZyhv8bug655+GcwPCD9jXjBD0/rUTQZr9fQmleDt8DGNDV9rzogZtZfGfGDPs7ON+t
NKV8fL+s0cKQ6lTP/+EKuWVHfQ7La1b+IqRoGquI9E5e2ectkBpQwX3DCPwYjTNxQKxK00wrCXGX
2lTFz7S7Q7dJIeCyokyLvQpdyz8FiPoirkCrtaMfIUgFcdgmgBV1HxNkWu8ACOhgdQBbu/yGuXtG
BMTT2TQhWcuvUZmsC+x+C9dcDaelTgO+up1rAmRithCBzUAc4DXmY33lqQngaILhXL6gazqWh+ai
S374ybfo+t5KP4lXYUemRARZMkI8bhbdfsXSGxVkwuZU22rm9bBrHj0gjErdtC/ZS/PD6/cfwpZP
oTSAV+LOyb5ai3utM8eBObbWjHrjXZoMGsGn0BgW8OM6rwkVXOSz4XTii2AMc+jQs6h812T+GrNj
xAqfRCUEtocXeJM29WOf8Z1O+uCTd1UlKeA7A0yzKqBUp7GH7HsdfTsNxAcbUwSW/hMz8IHD+kxy
66Lg42BSUtVThwOtoL4xmEs2db9rbo71uEI87U+WzBqf1fD5aXMSZFk143xxEYWu2seWrx7RGjn0
2huxbqsi/Ysf46UV3GX/4Vcdi6vhxDDbZrU45DiM66x7dvjHObiB2Tda0TICVkix7fKVdieHcFy3
I1mUuxznBPmlzkkni54JGIdzu6VYX1hQS92domkG2tj1k7fL6/DamKBwZBv0kKZQ6f1d4mME26B6
gt1IvVwNKFcvb/6OBZVKrKksFNUIYVIKaL6jE5MhPTq+mKy2Ttt98ndH9YrL+Z4lU6GPLreiz1ww
RFP8eXCog3w4azamq5WvH1piOkfVCKGsyMs+lHLxX0CLWztbmU6sdNcXyE6lRkYeMv6s0AbDjgap
b1SUCSanEZUPKRTFRd77I//tv/f3V5KMQ1TXaDYpMNuZLlP0WC6MGQz7nCVZRuO3LiR1nmxrcdg6
zkbuMUM/btuIDpwtf9bd29e0xQQlsPleFxgZkGJ4TQUBYT5B12ZWGZsO6xOYOBxlLSfcJpBorVas
6DPbZrVhohGT7MjjVcJGdpjGu5NBTjaVpL1hFBfOOUlVwNT7zVut26OcVxo+aJ3TSZK1As197Wrv
/WFSdRE/rvvdoZfi8n1ixQdfMUsFuwfl9D6p5z5w414bQPab9w9t3detBsDYECPi+4JXTX9C9vE8
EvWnoLq5WqXBM0IoT2GmxgVgtNDYdH0BmUjS8faQzXY9/LsKcZgc4DNzWjKM/ehMiI5O0SBstBnS
tbrYAa6ITexLxXFTlgqsVLJirasexOnuqIGjbGb96XF4O1Xhm9jEx6Tcy4T8kqmlYAUY2YwnqxeZ
pOUNwzYYX1B7fXxWLkJ0WFvq5gDtFFb7GfaCgkpd8zH+sBq2alIwajS/VvNmHJ/tR491XWXctrkw
2K8nXzUSadCol/OR5rbqzqSgfQCzXcR/wlMeUgKNzxamDeZ2mS1m4yV3V0x3ATOWkfv/av67Q1/F
kaoTjQElDt+73jXbBHMs0qtP5zxTkfnA7Q1YlH2iE2h3l+6piICDPOCQE7NabNLaX5Fo6l+2rS27
uBOJOASCRi+2gIhVc9E5E29H+jKgfcdnuRAvrc8eZX4WEvGFoOqIcR4kc55uxil3ijSP1Z8XmRor
Iya/h+butMxc2CqC/nxBOw5D4oKFL7JIWtWTB8aFNGHzDs3CRHMB32UoX9PwkLLxIPMWxTzTeit3
RgdeVu5D6fi8Yh6fknisyKhd2UI81/SXeFmC6e6wbxwkzny2S7WpWmaMmnCxOwvtFYzPY2ElK3X0
TWmkLiJebxN7dz7ohiHreKWCkW4URuBdSWRTzCmRpwxQjLU1xlOVLvtecmYtC2HCChyuGCu+gPud
oNOTx93X+eKEb7dWFDoVmuir8gy+9sszq/RJWa0zj6QpvhlxS3GTfo3ePknqv2t2cX/F8Jr9nVef
qSyCPFmCd5I2sOXfmvN7rOwxXORRqV6XucAGyVq8eVRiPdcEgSBNM0ATkEK2R3tqIo5no8J3dbpd
49xLkf5HvI/zGukyiLmgyCogvVwFKgL15CbMHhTim6klOOJ96yrumMij00jmxs0cVWmBm9OeE2OY
Dub7Y2cLa+OOVeneHfp3BBsTdtq4jSld49tLyAkoRq5VUXXMlghaqjyxewPhU9/xTrwQAm/iJLMZ
pyFuyEJ0I+jn4IQMJqFfnjl53u94eNimN89rBzBUg3z94oKKht/NXxbUG7cvqMtfOYZrDEIRS2aA
Hgl1f6eTCrPSAQ6tCQ/IAGl0bKGQnJ8wd/jgGAUHB85ZTNAzIPbPUEclZ6O+Wr+Xw9BJLBgrTbH1
zWpFGQUxXyVNMY2NoyE9JvGdp+YkSMKV+JxnPwb6EX0L94MbcQQOIT2hXSzQm69xxXIvC4ETQn91
9pxuhAOZ/FqEpgNd9k6PUBe2TURYsRYlpSYoJEmGFW0Pwn+9ZiXOfIKXxAvq4QFIwH3TWvHT0N/t
0QkvEY3ZLgt0VprBSOHcPv8RJHZxB4Q8Io4BnOgPFnmYy4lOBl33NE3k5zNXr1yl1ZOiovTcGS4L
Ze3HRZFbcb7AJOYuI8oNKmePCB+MihR/2tzMkc9zqRDo3/PALfqjF688X/kYaHGp5oB+pbzmU6VW
nwkBz62RLfBjabPLLwXiD62VIsJFC8v2ax2Cjh+GfMTwpssRqSV0GaElKVMrDcX/jWOsr7uf0/6D
XQgcGjA9jvGJdSpE+5i4GazDWsKFhAbeBv8Kx1AZsyUQC6383kKKFJYz7QSKAmsxvTynliZ1tSv4
A39Q5RsPtt0z443HFSgwWQkCCcDsyzEQIILWBsiozmMRcRkI3JHio1XlAb5fUlJiyqYtQ33waBM4
9rfESFEbsdz7kCwDHbAHpoO5veS+kUrtuGMLi7pdnAg372cxDJSyCE8OM4Tj0JuB/rmQuMqkHhhj
Ojn88MV/JCMNF1BXC6gtXtut68VTGkvUDmp0Jk5cn+obN+3q1RMYpiLdBVfVFXDV9WI0H4RlCJP1
PJEnrTw/v/afuN1QoNkgpuDGiJLXVatEnGnfZbYvqeEwAYq8DewqG5F5pQjY04tNYJlHMYXh45lt
41IiEgyafPrKvyzlDzS8S7kleWnHYCyU1oLpb/YYl3fx91iqnQUB22cCP4evDY7Da2MP9mQMBqdg
KpxSb9VZJhjP9j7TD6DkGsMiicv45So6uzO/W7XrTqbMyLszCfNET2cPlIx1B8Bkju8nT19gMSAO
vszml87MEhhXWZGGMUPFcXHu+Qzb8/g9LEOI0R488AxtgM1+0Y+w9m3RTuPF1uhoB2kVAxo02QgU
0ZXM8j0SfC+hlSCitkGOuzQPLKBbnNEA3DTZ2SBWIRw2eGlYRu5s7wXebG/xN3AdWWkAVPj0yC53
3e9cAwF1ikfLHQHFgEr0Lls0RtxodoPi5fC1h4ujjPJXq7FQclBFfX/9Apz/eTUk9i6MkxRSp8HS
6gc/pfH4U1qCYXqsucBVO43y9oCwfkFlmgOUtpmZYUCBnEIHnvW73lvQdhWLkzHWfS06Zf6itM0W
rNwjs3/02Baat2NtjV8Si4Z2DOmVvmck6JKrBDQTdKrSOl6NxCDmYNt5+pWQcWNIjdM5niVFMXlJ
fMhJRdkWzcAIE5bnGa66CAmw5gheGCJQus8L5SazBg3RY/cWChNlK/KJwBPfKKYH8mamgoPRgZr4
+BbxaPkpBtYhPMg2qpGC01NcmX0KCht8ayncuXpnaQUYvtu53APW6Ze+6+QKInPJfQTpEtnOOyzm
UcvHru0p20CjcGAxytxC020Ox8IIMe6Wc6BAw8t0hj6YhdF+9Oviapf2y3GI+uKGkehaBDWJzZS9
yXuQQ7O2871YywXb/PajMU8d/akde559uk+mjLHwpt1MTAVnEWhz+a34BNpE7ePAZX0V7zpVMX+t
QtIvMxZcEfQ43b3Ro8tC6vzvPMyIvtaZXyoQBTuCUjaYKt+6KSpQ0ptvKW5SpypZFYNjVM0Xq3j6
nSksBaVzIflq3UvZeHGaDEuPgIWH+HzYSyyMAmYsCFmgqR4KqlnyoZ0j6s+X8I9nxAaqMtuOuqo2
CHCzhgGpmn+UU2EaYx0x64lRhWx/s2joKTZMdESqRF2vwL3SR7vilJmKUrj4LFSZw0y9NoaneUvc
lp/DetJqPSXVGaCQ71TdYzdvPxjhu5oeAuAZS40aU2drnwudPTfZyxEZnanwx/cHuUt2bZWlQ5y+
i43Vmfo9PhVMtNn8L/AFsjDiXQDNansaLKJkowIJ+hq0m5U0Z0ytVONL0Nm1In3hJ+RGRjt90Euf
F6UZVEoe11hktddOQjOVuLumW7QnrVOVy5g33guZZeNbabLflZCbqzha1xa/1Y+g0jl2Wj19G2sY
AmNqBK4kOg7t8rO04ZOl2TkNRpEAFglu89kFYO7j4IO612hsAU+4ww2Xq1zfNYg7gVd/JEUuxfmH
92urjouFAK/6kDtFGs0yQta3ELJIqpvLSICEzbpPxo0g0eRjB5eMTUYUq9LWjVxoLG1PHtKqABQN
K9LgCltWUljZvyfJqlVenV3F5becfnNuE9EbVjH/ttXmH0PtsvfJluwjnkZJiVzIqQ5s6csrk6Kp
tDRK0weGOlhHVVtKl3XJDch4fWdSgO0e+osUCa/0ncOFtfDqKhkguokuACId9WaIBdvXV0tVGaVO
Z1fxNnkrXx+1N6Odoy/oBdjW6NGIzIEnKIcqt4wpYxruKMrew2KUk1Gne6iApZP726hHqDMLwJK1
KosgVIdNYpwlpS6bqk35PFF3/zYjdVi/D/B4u5OAs02LBdFUuyrKPFc4pi20zx3Q8Ktm2so9yZwR
0zgbcezclY3TKkZgrJ5n9xJ+ppw0ohbKyPjwUz8c/HbNNDc7Oy+9QZhQbZkniiii+lDs0SDuOLeP
agttG+c6Kx9BIdp8Kr15E90u8KDEZ7hkvpttd0ujo3qWMLZpRsufRfRcmbryVyUXjgCRR2eK5oxW
kqfO+37Pc3lTPENinJEUaQVOgfRS4IxYjWFxfQ+LbrUrjZfitpl4ubwDTUg2z++70jgJ48+H52ta
bDHuGJBlAEt3xIM8Mkd+e+L1I7teA3R3Aeuk9OPW+/KBnJ9HjV7NVnPXWZ4DOo1KcsuO0/ECNGrM
qRmU5dc6LAmslw4gZh1U5sGNE3ssN9sy+VWoNBPKOeW2UGC9cyY7PR12XALVYJzd+wEqGG0Axfak
QhyUn5JRLY4ngwwkoSzlQgFfYYt6XeMhu/etdK6RtTg4D8mSF3/8XRxXLVWgaBVBL4lxXaZz7vrP
X5DEP2EnKfK+PFD4dsFDrtyVkeYXe8iTx7J/6GnXHuiMURNkzf1SXosw51bi5nySkzOIun5W9dGp
CAtRRXMIy9nBrBJgCnIhiBZxj2KUKjoSYe8yjWae0SfWQoc3y4FKIJzGmg9TuN+gUMhqBMPpKJ6b
WbEtHfZvSy93jZ/7c0RS1KJ35Uws2BfxE7pt1/r4DVFvvlrxqXsI/gOiZubvIYKJ6Ya2zFGXyfiJ
NlH+EbTLHjlaV6R8m6fEHZZ7fPW5VP79L+VQ9Mlf995OAf55RbdL9sTy/3cFeWy7Q4T4bEe+qRWq
BdOBwZAMhP3UB5T7LrFlwdXdd9eeSjAneVbi/EP8r3jQ0XL9xW/IcbrC2//MVDk/wdYPCnhOsHjn
LRbElC/5m6Yfu7qj/WJO3NOwJBb4+Lkllbp0K5n9P4fKcrPfv0V9hi+FmtyQ0TaVFf5fJNJlYFYW
vg4b7DETe+6GMcnrMFyVR21x+g7l3hKUpP9ja568v5JpGrIZSgur8OX513/uvdIYnDXCEUUS4y79
m9Ns2Fs+XeOUQvfk2WFebVTdhy85Y/QKFo66gQkqNh+T7xxAiUO7M9WYwJwrh66jSq19PplyRrBa
c5jacEai7EFZobGMqY/rBk78hT0S3X9C1KFhr7tNZNeZWJ7aoXIBBhyL1e+UH0ZS7jZhs/VabxrY
OIXlkFfgG6deVodlNkR9dhZnBbhiOdOLounZVkodrRgNXQ/LXBLm+ImwvS33SKjOZoJWOBmawFIz
m86//65uJIRT6XJmHi63J92Pazws8DJXM2SCCHPl8L2cDuZ5S8Oi+xahgXfuzNPSNQRYD6Tun+qQ
omN1cm0l8CjKIREt6PfJJRxAvS0Sm8h4A9XfREpaj0FV6hM68CTQAgt4MICv8QeKR2SzZRy9vsxF
UAfpENg0JoILbcSzhENlBQaRGr/DaJGQTm0UeARwdpI9brublZGGRcMndgHt6BAzRAHBTDXsqx1O
UJoxrXRejZG5kWkKkB7wIvkxzEBXG0CZS+8ucPOiNyiCwp7VjIjmogarZ+Pkl5PRw+ABivwWOazr
wee1e83qJW+wmg8Sn7dCA5JYOXT1ZXhJGekUEQrbaN0Nqdu3ZlWe3WWX6EYHHE32+nKv41SvuASa
Ao1p/a6E8hpC9PYZaXuoS1P+bkA51yX8n1XtO3xxKbjv/08NpXwHGKc3GT7gZczDKTJcqWWx9FfS
/mYVCG5iF9iA4eXrKBdqMxiNLzgHQWNWJ/58nKiOFSMXXRR22+Wtz4Pl1jDzaZpvqBYtUyemOSh1
xEEDrTtsS51vcDbbnw3XrQ4eZlnxjZkOBVCV0Lm6E6H+GuUCEWoOYDzWfaqD4GcvwK9fb3suAXHY
WYi8k3Vs0n/uRjnSt9Kjw+5OstqgDLm/vpvFdaS/6D+z6UKc376ubrIcymJbngn6UVMEIYB6rcYn
BozveKbwcit8COVHKkCGO0vjjGBG/17c/5YSmuLpFx4cd40hSndh1Kbmk16awu16++BcY9F0/3CH
CMe4L25sbnmWzVqLhUB08FE9Z/LnBtCMc8gWgg0VgOUTqwdABWPRlxrOsug4X7/12lsCvtnxlVcz
wVaflx2OQNbJIDn3SBaFuO/j4DKHppZDyaZYX3PX4BGo43CRak81q8Anjey93tG15jCEz+hdb+He
vq4ovrIp/+DPP1tWJIVoIejVVOnySLhNRO0IPj5WHHtNdpLjtRiDB8hb1AR9m+Hldc7dT1wf4m+1
rscv4TqqIlbuX5bWHy7yOrRHPsaXBZkC9KeTu6r+1THeN11Nhs53SH+1yF75ucE0OmG/xI3YhwRb
LUqrox9EHUg0iJbu2crp+sPCGxuzSfWMdRs0X12o4XFrxBxzTgl9dFTnkD9aq1W1OexbaMzuQUP+
YHieHzgrmeAJ84rCmgl7ST7mGqju/j0XLbP5wrosKVr0ZJO5Q6xCVn54V/EWpilf5dLD3cm8/7XW
8ZJNof60jSejAaF7rKqPztfW44HSUIX60Rstl5peeyxBGLgbjXchNMS6BfPh0YGCsfcfYkQorSmE
Dx/UXOCE4KnnzU/aqYSGLygPexu9gTxft29ZUrKat/oKfYeY8q/Vr/q5f8bfAm2mnIRHHfNNvzHo
okBNIdkdor1jJ9VEIobHezrIyNOynQCNk+2re+zA/sVkZLmlm6YqNnBKpKY18AxIygazy66hAh4r
kbbgb1R0PV6t9MYmxhlMdkzOgIpVxVsjm7f5068+PZRi5yS+LiwNyb4p8CYw+dmuFv3xpZr5Nxt0
yeNNf9Fd8a4XQ087kg80AKEL33q1YPr2MarQQDbKu34PytIKwhd4f0/n6MlnyfXi5SESJ+8o79FU
4GOpJVkBArd2VPr8+UsTAIHxjY9mbYoPHbZi3RVjqCXkJfH3PNsRhpwXI8SQFcy+Tc02llmvbrXq
L+Dtok3AjRXTKl2nE3+XW0ph66t8jAvCejUfFbShM1XdgD2sdkCkGt7WeuULXgY8f+LNHT7YfY2l
JHj/XgEzsFoa9Mrylvh2ujkZ8iyoHt+6OPtH7gL3M4qXblxvo/yL6n5cOmnaBhVNRvj72OTmbN+h
nSxLrazF7lU0yqpisykVtVwKa8KelX6ywPRhCPTxzwXK3oTqMPbepwg6e+QyviHcQHmMsrhRR0/c
h6j/Tro08rvdkDln9dg50OYFkzWYgiAuxj+TbCweizTcSObssIDWr7Pf1QneNofPirtmwlHSigMR
eNcji/ZWx+q3jryCwXXqsE+vEwwpUOEyaGsuGfHKggTMhkHbn0jJBai652Hl0Gy1/QpQakv9MNl8
vp2KlpI8OFwE0Lhtru9cconJUE3/O/9KExanf0Chrp2iL7rEDnEJeuPLkvlcZ1uxbDrPz2A+6lhD
w90kr0nDl/Id/Ys15ynxCFl4eLrG+PZg3orSn206VbPCByvPKE+tBcrMynBp2dqW4q/RilXG+PKG
6JvCndJBBV6JlDouqljdot2QzEMhydvVhdydLisp53ykaIXzSPzH+ZmJqCbkoqSKFQEiiLxQVIXc
0rGHhgAYY+gUEEkR5IZ64Bxuon0IcEdbykYwe+jmFD4H8JBpTwPFG+kv01KEdGTQstLT75t8fDYd
PSlxJLSXmitplEB5D/d+QOdSIN8I3/dOWWH3FDS6O3iJRI187G4h+P3HR1yuRvdxRC2MtEujQYTp
Pqyb2SZ6fdgCAsbJqaqPT8Efxi+Jb3r6gudk9Za3BxwUkY1UnNHXYwSJO2Upi7b1xeV0RGaw/+/b
4gn9yAb7wAVatS3g92t+gXTfEmcnnrKz+B+Cy8Yp0JOfjirlnu3Q16gLpVGeFzFHI1RiXMRV/699
SdmCCZOzPDNyb78qecbsFQv0tbudU9F/7azRXtGZPersxgqS3hMXy7eOivvp/IJmMX4vgvg5JPh8
VkieXbCt5ZNUdNVbVkYLu7ZQkVExTYM+7ZH9ezHzS9QfjMoKdgLtYymC/b8HBXQYk51UfYf047Nu
tiGsNqVpQ9hqtLvqMHdxxV61DkgKF8qVdJz5haI4T5x3vt2Pa3rl5/njdHt/tdDjX3JQXyjG8uSz
WX8HNGbd0ndqFqKzDmnVYd4448eHaHOKEP5S/klexxVeNF0SjKQqfKo6zaBWPDGCKnvE16XJfkLh
Xr6WUjaPlOo+0PxBR9Dz3Mi7FLtduorDqxut0ol+vuVwIAElKA57cWSKxyuyGpJ6mwqosFf8lfMp
aVDw7uz4z8ALTTfEV5gYvIC91l/j+R4oHN9yvlRuom8DCdK1O1yVxw9IVi/PPVsT9oZfswMUzcqp
uc2c74ABtQep68Y8XBvp1+4EtmhDWbT4O4OVtxmPkMQjh4M9RfN2Wg3unOCPohcbSliSxALHuLFY
J7vPJn1q4mMEWfHKpLl5EYqRv5vY7U244h0MiXUouL9/EF6IR85y7s2y8IOIex3NMKrPnYq5ZwCx
+9A/nVThdnXKjn1PXdNaZwD69J417Uzb6lU35Gt+/1kvFgB/EeS5puDNBoJR/ne2qU126L6SnduW
bYWbPUnHJk1/N1iKDUxx6LSk34uWllJrwTGmYpqLZqmP17BakBwIi/tCEDkQvsdRnZz8Wo5jgS34
iLuPglV+W+gIqG9JhCqK0FrOOVdquthLfbZbUTXvvz9QSb3QuocDmaSwKc8gRqi6HCWOKz8w4jtK
1R77UaZxSL9DVioFArh8Z4ES22oTL/x3iq9woHLNIiIoYxhYrD1VhMFo+7Xf2o9gCZuskZ17bSHH
hOr+Zw7xq1AfK6HICEIqeK5x60NtXmbDicpLNpW03G098EhNeZdYPgvhg1KIWwLuvlS7zWD9gFG4
1ahQNoHZpMZHjH38UIon2VsbXfazd+sjtugtoPj6++cZDjeRlXFKiH5hcdAddnIlCht8a/ozfu1A
fwqE276fM45CJCv3bwgDRoTsW1/+N10dtlDsxD29ww68sdzzrTX1+r36kbmCX+7ro+ZjxSPbZfu6
H/qsVcJeIa2X/+rOxVmmLt6QiXDQ9wWaidc/CkDHewNwsrWJlsoRfvvs3JcieN9BYoMbzi16Zf7T
Ryz9NUbC2ucOrTs2s27F2uBJmKH3OQ1oq6CpM8PE3AdSfg7/kouUdhiVQrEmi8RElvIDHRfKS4GT
Oqjrho7BJzcudCGdu9NlYp+/JTIlqQPjmW+4165gS80q+L8U1q/EFldkn+cYbi8XwBba6Z/KtT7/
ChmtsCfcpOnfmtUp0MEriDqYgt4y7SVyGpBjfYe2RYn8hntNZkXjjaR1L+0gAjyY59oo09T4TUUQ
iqKNKu/Y/YIi/O7dz1htoB+4NvY04uQwZ4HXJbLy491GWEcHcQYY2HeIT1NC5VIKm52ONvN26Ci7
XsISmLt/DoNwj8Q8ip9Fq+pA5vHhB4hTu1yrnvAFO/yZg7mAunyItzfv5sTNgVEr8yI6kYICULsv
XH+BVJ/TbihlOfQTMW0txcA1B15fftEqWqrpEu9ZlbF7WD4rJqBa6nYIB31rdj0ISeF2D1A+EeqR
CAMfJ6sW6K38J3LvNl/8eyG4bz+J7z6S4cZIKV6q7aJx3ODmuBFM9p3OV2DQq+t1aWqCYdRPkmjM
AnUJijYFP9wmv2bRwLz53cWTwO/8+w36RMSmluKdJMhxB7dfjDZ+CTgrqfESehgPnt8ub3nkzgKO
jTBRFNhGYQoemaUWry3CGI/4+xwR/CsX7RaSv6KkRUJlIwuuzXeANqFOoyMQgM30F8rv0DFlh+Am
4dToz6zSqadE1s54eBX6hwrSdkG8wKfjEzE26UWD809jJbQs9H2f2qvgBvgEA5S92yvH2O3GjL35
4F24lAs4siiFR5ArXgBwNop/Qn4IMM5xQt3D1WLxrSeE8S2XVwCpYhY0eqNIutaZsGe+lJNNvXxC
avDMIehJ7mH971If11kUoqEvikcfZXpGdaKADGdFlNVun7QYg7CraZ80NdwrhD6glBj1GNJi9TMV
jevsVQmwCYg88V7JNvN7nUckcwZTlwhlSlxDrmFWO1SkHSf3B3Puk0jUA5++yAktfyiXcCX+YaqE
+ZzQ1rt6f8k2EzS5jLgJbE1sDee0AOmAVmOddrLoQrKwG/Q7iHclCJpWQw9H6mZqyyZBsKJ5FPLe
gVP5hl828vZzsrFS9UeRo9PDr+nvkNofzpk6NyJatucH32zXwHgcQnTax2WliLaXdEjSJJXNvljl
PmD2oDVoq5a7Rle1+WAOTNzc4ENoTsxxNeg2GFkGjQ2THwtYVQ2wzahXhHpgs/FiYuFznxKzC6fG
BziHA1I3fLO1mxbYWzQ4oZ1xXo8v5SaleAXalLhQH+gaDdCRsmS+GAXfFuhKmkGr4dDiA0HziTQ1
NbaqpxS/px3MciyeyoR2TdFaYUh0Ndqml1nIg0QgZ7W1dipTFyRk55fKFjcrz8Ee+XyFx/lNwbje
nD92en8oBQx9WT4VjXcAJqvW+fOuK8NkusLQk8Jv0MoajjNWQ/qCgl5fkiUmHaIsqPLjeng1Rxhp
RIAqWZ9c284H0ZODD8Ski6zglOm5wUZJ78EXK+anzkX7wl+de+YTyEBnjbPcERp7UGtpCSjAluD9
EWC9kGQQfU/xmcK+8yVH47C8OgSB+HcuI2Np0j41y69ffDrGinseTYQVtW6HWjmgOgvsPGk0i6Q3
Li8aat4dHgNPJfaZSujkVOVHIpYpE1fnq4U45H+3pWpJE//0yggTAJRzmpmTVDdxGAFb5zu6QSMx
wktZqvGSRTXCjWbizB7+WVGThQ1TgG/k3B5ro4f5vgissj+JG/jgNYSt1Uq0slE4e+nwfMYsvAZ2
YPul0IKyrq5FowHR5YitTrbSlPQB2Lq8hvhvLNysrnm1RlPfdXjmW1012ByOMB7fe0OWh6w/SbIR
ixnpLJvBOk+bXeFp64kygqRyicen5B1k3cVfyIMTxzUnCD4T1+iMfXfNSG2JJQgYhdqBX2HkorwA
HkLqwMZlv4O8RaFOpnZl28gwiBWd/EvxwD+uQt9/336bPgA728X8Slgeu7qf4Yp+6FgHXAvfiC25
D/ka5USoudjbnxSwgdvmd5mS7s5/U9NIA+EKlVynKASd+tWl1cCk83d64dPcL5RFQqg8dJF2ztAm
Q50TZKy3+EUSr057Hps+PpCDIlHYlGQTFI6cBicXhXBS/ZmejCFmMm3+m0tjQ1oliFK6MRwP2XQs
dElcDryK2naUplnTYrMAggSW1jNGih3Yb3VYf1JczbelOrpcGF+nP9XfFZBIoxQNtYKrBKVVv+Vg
noEhpsG5Qcr4Kcae80T2wbTzvLPTyvYro/Is7YX0lEXP5OxS1gZZqLje4RDEyxUr0MMwiCVK4B8p
o7gSHuHWkfaF7zi7ScEv0nszGfdjNuyC42viSc40ryk/l9IW8GV0rb46k4umJ5LCCV2hjZIcmfXw
K12ETNRqsRoLJAMTKJKz6ngoMcTqbalu7nIiVzgL7ghSyWvB0QyFDADnL1AT0N5r18FuW+bIiGBu
tWA+cWoEaG2AJbm4pOeAcnaNe3Xsj+i3Cf4o9c5cAiWFZZ+NhbXF3ASOyyf/YgKsJD3uSQRTudl+
06JqRdcgylfoOF9f1YG8Wve6w7phO11NQP+RECLrdyHr9PZXMX7n4+zmzkA3c73xE9SkYfhLD9WQ
8DxXz0h+Bw+5TERLxo6njpGF3fLsZfA6COb26BdhdYxl4qlfabmzQsaWQmdfnTvyyhe8QJveLi2f
CIAB4UYi1Dqv9P/EQucubVBxrOGFGm+XRIYd8iSMv+PNdsXGAbRnfUSHyKgzFMzS7s/VGWuc2Y2g
MF3k35V/y7YYSAohp3c+Gt0euNOIlGd4G3/xmqpgbPbX+2xYLvF5/No/Pg6Y5Tnk3oo+IIj+I8ho
0vk7MlaXRIDcZKmIgVMy0w+hj2AJCc3xn57fJ3YqhPpGUMgNtMoDWSNhtXs4aQogFgOWp8lt4y4r
0IamS7Qj19Zwk3V4SqzJNgA14KCSzbMriE/6ukH+cEQ6S9TMINx9TMB9TAXgBaQQjYosLhHsMKoc
M2nyzui1TLBTZutBlb9uaMByhqaUzLLUwxLUa09VRV4P/4fjkKivRc4nlL1dnLlrpDjmFh3zrKN7
IFC0vR+gonTaYyYXsQVpUeQrXgyGbYFKN+cWZLhd46/VIqcZSrfXvPhoO3tGijDhU7EUCIrvbTXE
JaMlQWFtdwkUwHj337wTFv6eU2X6W/Y2qY3NquhuiboTbDjZa/4yOx2UdUg5x2fcrdr2PbiG0aHI
62jkk5X1dWW2bOyQ+v3AsKV3PJ7Ws5NGtQPo9VYKk0vkv1g4mKVm6HtWotSIezdex1JsuTwzYqcR
Mq7WUmNTfVzH+RL4e308p4WjB/LWzyAnHUu93QK7c4i738MSA2pgKS5S68TMzKfpn9s5l81XuSeq
NahoCigigij9MqsbvyXORDQrm7giwjYwfLsjSynuvievoeBcRRydgIK/CvnF6lvnP2H4EnG8aQlR
Mv6I4xc/H76aDfMpTcUUZ4Pwhu4iD67beu1W9dnHgJ0OzFYWVz77yt20g1s1bZAIy87e5CLKCcYw
u/gn8mxtRc6dk8DSZoWqIN4ZsGRMdmriR5B/Yj8GM3KlRfkVPZR0ZQ5vMZhZwegQGsFzumDzPAAN
kfm49d5pi+TdH/KGLC16MNhS4I/kBhSdDhPWaOB7g3V771Dc2d4taI8+pbkXH2te3/eN8Ut1+FFc
9j4ZH0rAsbVXsZ3LPLq0/g6zMm6zRtmXinBLQRXB55zMj4lTh7YJD8S2frAFh0EP50Fqr+zgqAcA
C2h73ig4e8kHVt3ivH4HCmjXnTL9bmxrALV+K2GmY5LT/QAIl5HTgmEexoNrz/5JG9qgzVTC4lz1
Mu4uNKoSjidyAq90cLpTgC38Pmqb0AzlU9+sWM/HjIHX5fv21pHrbTzk3+udLY8brvdhhghCSPQv
9k7LsvxSX5SCFbiCwYPODDRbSF0fwPtgXWe5Oy+0FQ3qZN1XjAslWQjLpZOWzCPzrf2ePmzQU8Y9
I2AfeIMdWJuw3IOAPF2a83OMhIIaWxRwKI8vmN3FrK0fxuEIqfXLyu6FW+UKiFkUsBLOX0ImqRm0
AGsMeXe3EfXtAlECFbJUR91uO/vcEkuXm/fnmU7cr3Xmp+7I1IQ9Ih70vrxpGX0Imo6QmITKIIKe
1YTKc4mU3COUJA1lVnkc9aGXHuPkXzM2TwOX1QttluEZaSss+/Tv1llox2QhopxC8qz+SvX1FkmN
o1yfNh1uxMMN9AEL67Psl91LqWPPRBMsxz6yGcb/nJwn/o4Qmxycg4Y1DTiNFQBFRFJ/FHiSb/5x
Jx1TPMGau38+KsnXeKyU/24aOFMcKEfci+hA7EM52VI1PQaHjV5FRVAZyfW3BNJLeoAmJDwgofV2
jW+JoJ+4LqBWRibKlxmVnHCnDU3n+DjTDDpnLxba1H/QPpEUeAohB7SLLYx1eTS+1cxBpGmoO3hr
qggVmiGlI9X6+UjrAUfks4vwW1HGCRO4uDUiU4IGJw6xbLXuBRjTcJZmXkWqz+coCpO+nElGtOKH
y+16S7otxRMpjOIfH7Afd3bZXe3mTV1q3dxSHBQZZhq8BRHe3NMiikO2rQ9D3EpkboaOnriqo0Mi
eO8L3MNQcpPO+lzJwEBhdol9wA6lfHZHgppRPBeA/BXzQxZBDBBUIfHSlUFHRNeq+a72tgrRyGTq
zs+3JHodgbZTandDpu336t5LrZb1uERh616CR/y0qkF5H5HrzHLiASJt1dTF0tS51mFogghp5Ihk
RICd/3Ze2Z1Z531gIDbjg+PCKhvnbs0G7EiM8jnyOlBXEk9YVgKfJHGYyTNJN2NlGJxJWwGJHQbA
1C4hMlor1jaYW9d8f8shfaq4KbgaidMiZGFVqPyyBTr/HXkc7OH3wtev1rRyFVsAqUkWPL489Jtb
JfXD3xJfIDZYhrVSNl1h0J2vFfbKDpZrYtzr5I6ArjtDKxhklL7R3112UN+zFURarF3o6839s3T3
p5vPwo84qgmjZv2bFiEdUyFMPvGwjQtI4sD98V1Vsmt+oKPTx8eAjEk8m5dtCON2P/K1CZE2uaqp
ooDa1Eur0larcL4lcuptzQnsQnNJUDriLr04ETdqsddjOSwzmCtN4sFVEZoP/SUCY5aWDsiUi+Pj
+7kRWgYc8omaVXnvWLz0+8gWHX5C9OPWKB7a4/k6XpnyGIXusilUusRx5/jhyP0sIohKqyoSUt6i
NI0mX7iM1LFnKkkqCAY6QvqDcAcfdaUhKyyCOAgVyq9wHxfdotwKLcBid8BEDz3hIyidTRo+Q+jq
wB9w9m0LibQje+q/KhqQVZJYx8iNK/EK38AzkLbSdkYvZEAYGKmaCEdIa2kLY5t06LheHkn+tKqF
8+9E3DNrrb3Gkv5G1LD/M/ftt9eecSt2rfKKFhYteHX2434FEyd6dcsyltqjCW646cy0wScINmhK
voan208dAWXqM+ENXmdmvCnUNCAVwHrPGuLbawzDAfF8y4Lc/XmULHW3NhN2sFJrSLfVcfw8azw9
e4O3NPgQ1+KZqcJZk+zlrfyc7OY83aNtc6uJg5Ty9VdveXL2yi1knSEcu3oOzAOHwcPqp/zlKd4g
27nvDAaWX/SlyaSve2mbO8ZM9v09NuNsDuck91KOE+GwqIMjSOaqXY+d4iKC0YBatZG1VRjYYjZg
G4vOsgdq4Lrz6WGTP4A9hdZf7jwaGOnNBBIuOwISFA+AxrK6osL0ISqnor6QGq57CvBQG0g+o5qM
i9ZGPKXQeFE39K1sLCU1jI1WegZaXCDpqZs/rq3TJYMPRx6+y82RV5OZTidEIBQpdlTcCUJxOj6W
EQdfF1fK4UDlJY4ahe3eczdVRnIJzqFf4fn2zo4H53HlWu1yKanqLyfVICd2j05SnYm1Cw7dJT1K
nSUpWPsHmjXbndvb2SEZZjKKJ4FVhEPY/gqejIf+QZ2f3pit/ZmujtgFGsisOv1w/G/lv8cY3jAc
TAMoy5M4XU3iKEuwUbAkCJDsss0RjlKLRSuy25JfTbPbvpiaUio6lG4OytNrmlsVcQVxzZe5B3L2
HbQE+xCw/6mwFbb2TfM/nyLhWnqiGY1GaTcZm2cpQnVbHoIuskL5kmlTHPtl4tn0Sl8hv/zzpfow
BrqcswM3FfrCpyqHK8S1oCfH271Pcqung57h0AEPIbtHz4m0R4galrewIrkAVvofUDxk69Mr/4H9
58LJM4388y8v3RCCMpM9xsoOh7utIJ7c1EtG54LQCxwW+qN1pt8CiiScoth1vJh5OwP59sFrzX9W
Ce7juqei0/BNoRzoMWxIPrAgcpn6YJwevGcXt/6ov0UUGIDRrYvzMBkBhv9Bhdt9Z3y2osgpiRMm
hBXGL+xlGoJ6BsU3A+Ps5w0x8c5Yu2e78nPBcYSacAJXhZTm2j0SG2nRRrQVwb8OU0EUf7nz6tWa
xs6x2n1C8vY0NEd5/zUyRcQrH2qW7E49wvRaHnP0KZy/eVUKcB55x79fcgdI5OQPFWcyJA4H6pwN
MG+sIPRGO0ozZL+4P8QCf9rg7mCRTsgDeADHk2i3HwevFbUndfJVq3CirxMcTyQP2kM6PHEzpeJg
yHAhVuqE6GP6b8pxXAVxIuTXL76uMyZWjt1Y0fJw9g3oJMbVN2e34cuPTgiT52jGYnUAaOlgMzpf
OEVfLysZkLqCS65inptcLZZIfgLkFh78b20tu0VlfbU9fmepIP2r7C4lpG5GhZEOmpneNGDOto3L
Q2Fz2Sg/L0Ho494zvXRAoliYASc5yZkD1QvBO0A+HCVK2r9FjIlsIB0+xACbKUVHTf5xZ6bToj7M
G+1mTISuCjatgKXVvLH+6XcpnKxqXXzEPWTg2oGNzUBnt7LUI+JoBVoszI84n8yivNjw5/gQ/YIZ
AMcOmRVxp3WiHkgKOCkmXcQ9cHLYsY7qlYIQM3RFF3c4P1NTKs5PHxptHCuaXHDfPca7WAYsGG/7
yi9EhCeUumLStMXFEYwy02tbA/dq07nWKyok3YFIReO3dwwOHA9wIrsz5UxKfaVPH3nmIKhZkTD+
rTqTVhnns37q1d9akThYOrFTxeqRCb+CPCzoAjLu6JMG9RCk3wi2EEgCiRl4jOt2Tz33GgJ0BsRU
gzKhvIMkC36uWKNjUSlOq1AOCF9HcI1BY6bG2AAzCFyppTvMi1LRNPy4p/EF+mndCKn8OR8sKGQq
vMpV+SVCH7pM4C0ZCreEqi6dSWn/8LFZzplfeySfP1huYcqQ0Qi3OANwe5aB4Luk3HjakdCK02Tp
zPcCrn3mXOYy/Ttb7ssui6hetXOCO6GdmTOj3CT5Mu0Cec0GDVtxi4dPe62eDmlQ8JN6tUXh1kZf
qGW5o12Z0SgNoVFvijEs1mAfKYVL7aYtIbaxWy7ROrpqyf1fls8ATk9omGLcchjtuMKKbAPdu2OR
40DH8tqseE9p9ipjG7pzXl9ZatG4GAmneiwtAK/ftiiBnFofC7KWgBn4WJKAdS826b702GKYoa+p
HEsexaPupItVN/sI2rm26aM5Si7Kyg4Huj5+Ex4Pu/TW/1kQbNLR9wZgvPe5ctixtEf5MvEAQ1mi
9iMFlXIQ9BS8LvqbOl2xb1Lku8xD1pBLkhquDXWcG1HcirFt3aYZD8d0RX1fskjkVlPWGobHnSLH
9BgVxi9h8unAzZQ59o0SZZXSie2EhgvQRCrzMFyS8fri1lIDF3088LtZkrXs5FngJrUHV/H7bhCy
GZWPX2PSQkYcr095eF7remDZCg+IK/QMVkAR35AzZz73dpRTCYUdyJRMxbbN0WZerIe/TFB9c3OZ
niZIbt3Orc/WHaOaGfpuN6kzmsQfzm7BNDCEgZf/8LEPUU8jb9z1boKepDbn/N2P9znbiZNqMgo9
p+sfRXyRBVX4deaZ9sR2hCncWDn7nb4MmMB+lftTVdTEvispaTqlCkIVtg3T/YWf34Xvl6OWN50w
L5JxofUqX6/W2EoQ1WRQlyOC6I+lgWFxtE64VPobJku8b8516mkbsQMzuVCDd7A7tJeqUfLSuJvT
g+wAjorLjcY1DzaxauAzxtyt5az9gyCpJZ3LJ1p/Uk+Tz23i9Ty3F1BkYaixa10EP54idCmXmZit
zjjCFHouQL7DWCGU1230Evo53gMl2PMevVDHIXn5QAKSviQpcH4Oah+5YMmGKcK57YAOqh0bL9PT
rsxsdZ8FCr5mzMDPMYyKlaI+dkkm2wgZUabkMBqIQlPV4dzIvVM9weOYnMZgJxL1dZD7Pv5XgxGA
Jg//mD1Rqh3GD9oqg2MSofVjS02x+/dQtZsHIX+4m7l8bp/QTpwsU+1atAdp5SrxIAhjzoN08CAR
x9L6qqXzGf+8phxzWcCniaut8IjMZKbdH3ioyq8F3h3bfRo2jcIeYgTC/7D7hk/phXIkK1tLuqIS
0mtZr8X1zhYuQx98Zw9tqXAoHzLltn3gLw7Z8MZg0bZdIHEVfXNhYDxvKlYNOyYgAlFFEqjRuBOB
x53aIVka3QW4ie3NA6FSW70AAkiWbTkRlNE2TjK40u2kz+m8gFIdLc6k1dMGKd/3fJx/USSp/EIz
s8T0AEFLXNzvgoA3zJy+YHyAjYIkXciXNOB9MHnY1xzYm13VbvXbP626/LaFewY1Zgk1iAKtle60
cxHzGPvNtvfugb0szkypSrzVwXw+K6tGYByGsGQ3lJPeF1xCmuGgyPo0xIYiTq1N92qvjCgvxMWZ
nyuQ+jvlg+/gnjQQxDeL6cURzA+iqYknQxJjnVB6dt290vxhRVRE4snzyhN4dG8wOXcFDqke+bDR
zvljvQ+JhDXHMY5IlW/iqmEBNKIYXh3NOZGyL7uOJGX9o3BMPYPoRp56IXaqsAasLTPFyOGg99EL
moVUUI2HhX3lFA2EJ2ePyiJWPKFMQ40tuXNm7iZ3KOeDnu+dzcDnSTGOroRXhCkJR86kmS4zJyJY
dd6GOdNrtWY01NEW108VLVr0bbAYeS2OQE+IvCkn+HappEZEPn5vujx0B4SmDc59kHNAEDoEVJTv
xcQ298dN3Hi/MSWkyX6z4+rB3oCt/BO13Vr39XomLAefZwyf53nsYajlJ92uPZdLZtqQ0iShHMC+
MOJqzQf10jy0N7rBpqOQZxlw24hFqLXxSZgb/TtaofLQzPqdSW9Jjn1GS/V6eQJiFTKMChrkm3fX
V+ctFn95xd7zw4X/VecnlcnzLA7jRXL1eDz6sXYk0U2C1wIBnxUgluDkxN/Gyc0aHOkSua6GVd5+
VwEpbwQW0qwvYQ3W4iDK/DKzR9Rs78feuWL2FAO3iFgeDaluWDjY1PpPGKB8F6H51kw2zHn7oTuB
/peL7vqb6YhNNC1U6U6hz8VWGLglNgCrsxVz+Syt1EZeXc4knoMDfostE+ddhnbKrcHhNZrEDSdd
B3HWm7MCnlEALY4z+nAL/cEbUOPgye92FkPzMAN/u//UUugLI6yPizUI+HRvugWeQL3DZ8uv+sKQ
Av2+A4nY4D5FIaJJETefi+JMLknIs51RBX3U/Lw6yz9TS0drWO+KTf5/3mtrvDKCmJkVeVL9pIb+
WezCLI0jyNhP2z9lwpSgRt38kTqkcA19OxPP3XITCP2hH9JqKJzRqLG1aiY3cBipzHJkObKmhYyM
E4c5hXa2ImQTTwCj9ya+FE8uweSLpGMhV6dxukuGwt7KvgE1LlMHhjy+ukecQhSrwG0G6B7czgnn
kGqk0pZEskS/nvuC1jiJnnrehd0tGo9yYzhyZS90eFgagfgtRgDAIoa1/mKqZkcQJV3akx9ux9WM
Xcli0HcGVnCQLcONHUntGtKvowyyysDL5a0hSzuYrVj9D/OAhI7n102GMPmJIgRyNCeDoApCstLI
WlN9h/yEIx6rU/CcyJ0SJSCbM0bz5X1bI/tnGwrOmKydWFhtFRBUpf7BMIOQG8BJWG4whgs1MDqn
ktOR2Vhz5+qxLkx1yjwpdZh2LmsX0iQUL8E0bHSLsGoP9V/ePfrgz4IURG3CV561Svtr8IRdBI1h
Tl/SzfphFzVT6k7VmDZ8iOQC8b45wBP2IOmq77WNbHmfwwvZ6UOG6EH6PcDKREGTN2xras0ExNUE
wlmAtYx5yyZ/c3yjf7clVgxr6ScS+F2rChh2j7xtQCzrwcCTIYS9/33lnTf3Dbf6rsn83y6N/XbQ
4XKiNo++Wue64UHahFtOKM9EfSQ94K0AdXWcy/rlPN8qJTNonD6EJOBHOrKZVDxLKeydlANu6Vpg
mX4/oHdO670JzOQYPfwNZPNrjyRYdYhcTmX5zbyRWIBzNCXU2FsPWxckSYFr+F/HSdpbzIl2sNXH
r6ndCeCmt/m2UkeQn3Y/NcYRqozKB/rADVPup96D9aonjV8NCcjOOjq3oMgbBBVqPwJqsMtbjz5l
E2FjUiKr9+IU0kpZSbbMv6v73IH9x9tQ/EanXmfpxHJgA1q272oXfl5l5bvxoy2kX713oEHFtt2H
3i7eDMkDXRQEDNaTEIVxCK65FV1rf5Lm7Ooq7F+QA22ABuPI81MRC7d5PnFwydgVjk1sqk7mPHpI
iZlzH35C7pxxdGN05XhV2I6274TlirXf4iA5ykMvE+L2FuhipmeitLaLFXNTjFEASzeuqfF+wiKJ
+WPxKS0POGXTXLSIza1qXlzrBRa71FF02K3tUxLesZLL+/nFhYr+OS4WnC8yPAhjDqFtEubtgmCC
CQc1LQq+/9XbfmZvOe5TviiRhZatwDYhu0iB7PcRC7NRBB3yUMRHwk1N/wpiyfSG/+3zIqQ+3tUT
M9DA5RQLjiPy5T5KZQJepgRvcdxRxzSuSYfkZztB6Yu1gAkI3kcEpWNA36VAsBifXFhjh6I8TeWo
LXYw3TUmv7I8MXzOPgYsUivuofOaSiegEi2t5LeQM67hGk5tM64/7opWSF2TfTeO7AgEluDhXjAM
dMwTc/h3RcrBITXFQzsimddFaMQXbBmFMKUWpU8ldKqOY6PNV6ru4AmTufasBxf0u942w190nm+2
qv0U1CtYPmR/s3npJlaqaWsH2aZyl2qni4PyJP24ntIwJGwFoNoOLMrx1lo1JrkE54FFsUitCjpj
DbcrMturDuUjh15NVCdayCu9KKGtRcn8x26vc9jJFm3gTHEBhc3aw14Z1/+jqkyv881FVhdDj2hY
+ebPXqeAqtGD5gUf+JKnCDmA/euDuNj94945qUVj/t/P8lY/keZosB0Bal6tp6HGXr1CJOrdHnV7
5v0ZULfO7cI3WDcgPi8kZ0Q3j+BDgXIJ1I2/R2Ghu/2Xja5tNmxKfXcQbw9i0X2/ROJQGKo5zj0r
tTeN2fYCHYEBo1BBtP1sL6Jq05rjDrYfEYpXJpKHk3qyBM6Dy5CAFVO8Hx7T3WXcKuo+K9nE+wup
CVMYLoVmFVPSQClEL/5SkukuAcFWiAL+IcuZ3jF1bJK7OE5Gi33DJlXYADj+kEEIOCpfKB0hrURA
DE/AYuBFIFEbJnN40ykqsSOzd5Xhb5+f0KmdgHXA7bOGvctuKct2ZOe43KldwnlqvN9n6Wvp+UUE
QMxL6vjQJ/Fl9hPWjRTE9th3gJ5mq+ZTYs2sfjot3bbCOEm1OL9DZf57Rsi0BSkLOTLy+A268E+w
BdV42gtx6E64dEQxRdx+nr9lPyLRlg4Ai8i88SqGshDqIHQMCZYlc8BI4ilCATwLWL4m9aB0c3jm
iGIM+aI80ebdIrnJx5Yy5v2deLPeLJZ7bgETXI4JUvQecQ8AY7plng/rtvwLqsxSMua1NL6WK7Dn
HTmsccU/T0p3thKCxIzDT1OepRUZAFP/FUshQd14q0GAoLv+BIrn3v5sRVK2Z/0p0gKL7m30/mX+
+vHA1nvKq9XfqUDF6lI1oBfQDL020cfnc48g/vZvlzW4rXBlYDvDPgsNmifatFtZUeDdkzfCry6R
DQ73L0jyCK0kaDdqjTzoXTVzPVervJmjgkxCnShUP8WXoSfXa5fCLjEfPDs9sRysP+F6+OqczUum
I8TzF85103wSIlWkGUOzjM1+KPZMVQyRTHyYxQSCvXXmrfcAasXxHeHkQjEjTKMGv1MVP9IU6+tQ
WYV3R6zLQeo5jdgCDtjirTIkGeIKaW5toBk71Z2kItHyKSLIzekIZdPjvvLsRCSz5X8mDKwzJusi
YNCIYNaWxncw5lb15cCjhSKiIOHje6qCSNvZuZ0zX3LCLx+lf1LJxq9fHkCIDgLHPWbZMZHbPRX/
V1RDATyb0gtZ48K1JuVSbwp5xtQmRDnrl06c0HrAmWBHecdTQzZ8zkYixA6EgytGNNhy3LU9gb0L
Hu0VPBbQLo6tcDfNUXezEUBT9uv8AG+h0rA51VWZv5coNsr3/kfx3wRp21f9WVxqdBDRtv+VzbWs
hGAuJNc+MJS+uRUrg7Y+njHWcqUibFSm2UfjCNi3UgisVtTW921+e0YmpGgPwa5Jeo6nq4WzO8gd
c7TX4pMTOf82oT+7zcnAWecww5AxmzYsU/VC6j2e1LqOgbx8GYy/hG14LpYkIcuIEaa/U+q4giQw
pLMYK6K15HCVYnaW1Ai2Qkt+bq9ZXObDaH2E4rk5ZNQcwZjeLBYAoxT05bgwK0ytGH3I747pKcgz
ZZTzkhqs5TcZ2UYjWZinlnxyixWVh3y/PQ2cjd86LDhjAYhDtNsvTokggObW//xRI1Am8aAja5bG
vLcxyH3bGL3ptivnsLf1RsTZ4Q9XrPo2nOeHy49nWdASnUR8WXacGTgeOqU3SLObiR4mVnx+K4mL
wROJRi/cWdGGb18OfeZJlou9ynU03OP4SPWdud2POOzBnulcCyfgxyYhaYthR8pjitk9wLP0ploY
rTIzPr8KuoTqjhlQY97xC5168Y/0U1zy1O1i7PkSA8negGj57wOcacvIsMpfiFDkhYWl/xspdIBX
IwGGa9Blbw3V/sp6gI6VRGFcl8XceYncLTsMyoEInYfFoNje2rWsKI2XBGdHnJXF/S2ZDnDW3o7Z
+9l0Z2lgg2PrfZA0z7JsGwmgf8B8rps8wq/azE2g0FcywiTMe3dgKBpgAGhuyN8LvooxWevbuIFA
WJZ10ce+cdJtoiVFY1faVhhr4aLodGOIrg7tXyvdr4PkBArRbyz4tp4ICBFD58CQiW6wkioPXcSV
n2l6/9GCT7Nt/i8SJKzbQxqJZtP/zZUA6aC8HcR17BE9RNOaFLfRKeK5DuvoHPcH1sdyBo0Rn1bS
YJokm5CL4K82YaeIVbniS4jf0DtzKBDigRVzGsjw/gH2dRw+nAW5sqgE+18dVTXulUryiWXIXDIv
eiMe0ns7uRi/+V3m61YZKeIwTyMJUmZrWxlUBoX2XOTFBEetfAYfdE3Q3ynPLSciaBa5w0LizArV
oCnObrdrHaedSCHyqZKwUhUAezbNiLWuW5UPA8wiWUGNRlw1UGaYBqwqApdbD7clZEFBlGbpvnQX
4EQMsM4OpBeDq2fBkP+GOEWAB5PkP9Nr72BbnK17K8XxNJ/Lb35Kbd9lpIH4n7AVW0WF3EE/GECQ
PvSP7eM1Wt8Z+O3T/eO3wCeT8yfF17zYcAJNr3ldnTfcNfmiFdxkiyh663sFzN/tHekwEH8rH+6x
CwXttj7lbiGVlmHgqeVfEfgljp1vJ2UmybrYQPtlOnyZthndyx1ocdDMJosGpz30atNKupDGd1yN
SH41S5tScb4g5k2bjAQuFnv0RkWtHn77m1/Wax/cQaP83Aw2m5LWQYxQonkrBP3i9fc1fqEDTZi6
7Ozbcj4qYGRyDMCw/fPeWtdSlDpNxhS1iQC6bSvYRK9KHVARKYCGoD6x9fjXMbDBljlPOsoLTyri
eO2sGj4fjHBEscwen9OrijRVH4LUHj9HIQD1xcDLH6tst7RUjqzUHn6sBuJod1nz1+IryvkJhqe5
qzD3qUwV2LnUeF3mpiApy0UlCtZ+rfUw8eMX5lSp24OriISUsn9bw614EZNknNILX0MhayFkXki0
CTa/tr9rMl78YigZTxbb+lSjwK6GA80+vEw/SOBxibsV9J56fTvWFoiqC7rVXuyH3wFUWDeU738D
jcsjxyoQhFUT4vvQb2EdTG0XE3kWXNlJRxAccChHtE+ZfGtzuoMezSS0hoEZqg4Y+iB89HKHZttY
HaUVQhiexyY8NTntsahM42KALUfUpU+dzEV0Mz4I6icAoyk0NN+SjwzqtFvmgaknEje7oylPO6gz
n+FXT34BjxVNmzOy1wJvNNwAoGwG4KYVRO8scQGtt6mp6ZphkGBGYhDxabSzNLl78ekUkvHGAZUn
QNf3uLZmG3gmkB7q0+Ct8W+f6ju9cIy0zWQKhHEdn+zwUuE0OtJkim4p4bVdQeAC25FywvZ+Q+ir
n+cR+anLE11kpU+P5XWd/aHmwgZok9oQJqoYs619W1MyVCpDJH9tOtlxo6Bg1njEpge9JKh3gjAc
5ogyoPaCfu55C4xdGQOmvhtffEunRAwNLW349ZXo7suApT2Fmz2lBFz2mzmpRopdPciujr+wx99N
xhc6hO9YRHmXu9xLss7anNQLMSUTV4gFQYzGO7hbUimJy7KfYP1H75S/zV8fSvjcwVkmtpNILmew
2JSMaqFLvY2n7GswnWmxAYX6GJ9yDvv8hjIcz48/XiPwXeMcJrBqkpaFWQNlyJAUt25vYj+KRz8l
GRZYnv4wXmJtwvJq9OoqGnTUgCp4mJMzRhd5SxOt+bLrSVnXi0Zofyb6xXRog0tYfMvvIUD0xqqx
hpwcf6ysQtLCPE3VW5bLKr6qzSQRK0IkcDu4DXIFNWW6mM3tTIFI5uCquKKLcIcAIOwoXP3vIapb
cL99geF9DDvk8yVsy4HrsMGuSDePZqhIR5t3gxzCjNF4zmtvmMdMY4TOKpKHNXerHim0oWhEHiKP
I/U9ZtAr4EkrJxLVsDJvbiO7jbBqCrVo9sDV8noWfDfnbqGKrbyPEyE5daAu46iCoTHvnfrs9uMm
lM/71D0nUzmH+3mJr51NUhtrlF7zIwIbV9mXGltoA6khDO0hw33ltlnWyEo+/oUghGljXRZHYYRf
ivGws8auEYoZCRmPFmDkUWGGICjO2TcTWeg32UEWxV3fmCHxximir9xu7QJPqMrZDJQWpyhCf5sS
j4wfoxrrH0YV76DjCOm55DgrDi4Czjn1X65c1STNti2bRsG0R/S/h/4c3E6yw9rqrUhyzzWthqze
zvvap4Q0u8ykQUgoQ1nnsVgs7M0blbC1Z774xsOUJIQi9Hh4eplRAxW2L4aLG/aliDR+87AvbIjk
SfPYYStdl3gC4/YOI72ZpNFJCzPkG8Alpl1g6j+fO9Z2LniU0c5aVCb2yckKJ51F9PVyna9bc7uk
81aiGatXbMD5Ir3rHWkMHlu1Oa7h8/tu4k41ApS/zNgChuodUCWnnmvTMWRkIp301h9odNn1EMug
X+HkHVz5boT6aoCeNmKyTp7V0JUkYD5fsotOrbaZprqTynCWwdHWhc09KsZV3p5W6BXnZkB5EiOZ
rJ+d7GwnIYlIK8+a1p+zviv2UxuiqU/ZXX0Zb5iPVTyWsNdZBXit1AzaSNvi5L0YIq/hXkyBHHIU
MVdfUbDLLUSJiJBagQbPIS7bLwz/pDzTMqU/ymjgo8Oe9fUEeYUM/LJqhYZEFwUuLgqbrepsH4Ds
jCIIwGZI7kgERHlnhKzpa5NBpwuW6rMtiEb41uk6VIQLjmLe3/kFVRJI3oyD28zLj9VmVphiXidE
DEzkb/i2RAjAOFgKVuwu0zfC+9dD7lAliirLrA3f8oNbx3raBR/o+Axbr2TpcY6CMdJDOKQPojCh
P/c1WxoJbP+gn5KyCZTtz5fBZQNuy/Dt8Qr1Ukv29WZOELCsDnbzBPSl9P+QUW64zycHe6VAA8Ik
5Q+ysmvOTVDsvW8M6HTVMPAJgncDSxirU6vsw25HreVSBgG632QEo7ousw7xtS83ddWHLr9Xk0+k
BPUALf1Y6CB9xDprt1jsnETK1LRywPTyQhDr1ngFlX5j4LUO4cBXk+xCvbC/gVDCx9SAbZnOy0ay
s91Naa4jo1opOL6Ft/IQVnsoyBiApDTvEMU6NzhMMHzgAtfREbfjWXTdej1seXWbf5h7ezsM2JA2
6eNtMhdgNh4KZTG7bWTqRu50wgdDsdacpBNkHyDXz10W1XopWGC+Xugz6C8LPG2atNqtZSeiiZob
ghmePphVg13JoeKgZMZUrNQt2NaKmYh3GVrmWe+gVe4Y72hRb90prhi2jMRmZHVKYiOQTxQqPuyc
4Z71nRqwdD9UQ45BzEkMFtJw54B/6RuFZb+AIOFerUR6yBrdxCtW+kuGLfe52MymMRtyFRi7atAX
pv5LWWxzyPG1YkYF1C/Rqd8ex9mezARpEJz6sA1Aaqq7FdjOb4zNv/IzgLOufSizUL0e1BUafUYa
6LVTdXS4dEK8QWYw2D1ukwN6sLNENnGh4Fu+LCovu7rPEmg6tduvGWN0C9aJxpedtzskKi+i+AyG
VSs0sf0J+XB9b7vR+GWDfeJ6ZmvzQ8t26Mjh7/IYtkrwSKduV0Q47e01ttzYiXDiL+Y896CSSIhR
284LJZdrcgEvZ3L/4+LpgEKqLxlyoL7x4ekDCZA2woTt0L824dYhTEGrdAY5sfa8LYGStijKOBkV
OO/qWxMuDmvMBpZIOn8yxqwuvqKKrImuMohsSD38iOQS2A0PZ1ChdisV1oLGEOsk+ZncsNmihdwy
Oekzk9eCfTju5dx1XodMHyuUe76w8ERaWau5DHvClcSg8uG5aHn/mr4zaNO11KgZuBzMfDD89J1O
aAJ7PfIbp41UWtAU0xMtZvECvyamPaU1pa8WscLw90zfKuoUC8zgBNesO+I/phFp4XHF/TqJL7Pm
6rgmC8AZOrWRi6//Dz0WsfKr0H5e5SsMoCgAPUMaWyyladFmt8A5j6zEX6IPCqn+DO6w0AkFMNYm
EeOjvh0BaUd1Myyg7NafYTljNAQaOoZFoYtXJwPym1e2iBIxUZpq98N9YJ09WN+CHafgVUxCIPu/
b/SvO6e2EoTuJwldhlBj4IFGrjzrBk/NGCw0wKbvGZgHVhJvBk4oUxx0bHXXeaGoQZv1zgtt7PQv
w6W2yUKxvsjf+5rDlnVv40K7LlTq2fSyL9IjEOR3daFRERxwUTIRvsWmTHTyXOYMeNNiUlSF4PjV
2HyswFpGF+Usr3duKnlm6GoMJRwtGmabVziNCfI3PDgxSEvVm6yBmk/qzKYU8QdLVVhW6IvYD/Gi
nzcEInsFSk7frOx6c+UzPnZ5oC79l9kHOr1sJR5suCB+iph9jiZfGGZPPOaN8GyHsRt7WAPhDfyz
PWC8FFlLICQla0gGfeuzXK4ZhgeaD0QbK3XMPmc73xkwAFRlPF0P6IJ7etN1W0iwPKR4DEWxb0NY
INPEeFZQyVDSw55/ens0/wX6+waR3LpKztVKHppuazzCq8f0zW/dy33+3Fz4/KMV/QSlK66nm4G5
uFFKhxr67JStl3t0MrL1UtUsHhibTRUuOsr/fEfGCHOK1MyownTd8gbK7cVPmEZ/m6XfDLBLZB9r
dAc44dSQ0+WxA2NE78lrBkXdrCGa5Yz+3hLvCfposLeldSCESwsqXTFR4fqaPzG45fCOshtOHs2a
Dqf/HTmlFtjLfVEDV68o8i9N9e6YQrmXDEd+jYht+8UqzlavvMXPwHZXPDLahJTY9zHFQFsSi68w
P2yTXOKBi7IAOeOMb8dE28sYugTjOvvu7Ec+pbQ5UEmPS/BsONk/nyLKZ8JV8C3G2ZDouc4boL30
JgwmB9kmc1at1btEaXsQ/03UtosH9FUUltkSM1TvoVDexxY3VCygVmAUldJ+d+udXNvTiGBZK1np
04wTS4iZMAC8ixkjJ2n2Y3pCMmGGhd8gB9gC1QvF9lB79/37br3XHphVRiYJC6MFkaSh4r6xj7Ll
yp7ETYYjHfNCZP69WTqJn0VnN3x2ZiyDUidXZqMdin41sSD2+7Fn4yW1NHjVxAnLtonGexppdSdq
5KbAqOH6vAL/D8Uf30ALXrxRK8Nb1kIY88DzFJZ0+1c5rig5vGm3S+Y79SRj6ixmB1rB6oNEwCNI
5lVBremuUtB1UQGc1VfL7IHlkIkeJzT9VVjMcCOP431iyvliq5Tde9Li+XGbzy33Uy+GEhn+n9Yz
RFZqxe+xBkOX/5cu/YM9o6K/QyN1q9X54h/l+NXWMb61ffZLFga7zkrnpTT3x/e+owu2gZXktNCJ
i0PfLgQsNQRhoPpsniC3Fmg7qBmCxZBr/2hHVOCj+976pqzF9aHWjv7yregNVab+ujq/Yeca3k/E
slYNrcgYWMbs4jraKp2Mxm2T633Cv3arIjIH4yw9tGobV2J0jjuvVbRyL3MifmuZDzZCoL1rDMLz
ImYx6bRdxJAOjlky6bBCvz86gWqRfu6VgPSguLkEPoxcnV9YZJTC/gF4uStASnp1OUDnqHSVWZ5x
YR49w/odWE1kgsrzYzO2gtig5/j9W6E+prZbb6Fn7MvZ+euP6+hze6xjdfeuH0sH4S1J3890CJ21
yvvIG9k6n1U7l3E6gXpLYrIpF3cAhCpahkoQXjBvbFSIc0vJBZJ33t2WsBqijuLtxxp/iNu8X25l
7eQrCUQs3kV5/kNRRNfiUo2PUYWnKKNfYwUl5I7tAmV1TwqbgVQX19pRPEt5O/tukzvrUzMj08+J
QVh4JdiWWuqVtuqNp2gRTHtlCeTNp2+IwMwowAXsmXcookBEFNaM0X3UhVMkdzO81PJffe/fBczw
YLDOUs8fV6nTMyOITbpfKejy+aEKvh/o/NLploNvDjlRPp7CUVKe6c0W/i74KVyV+YQHH9QvVXnY
w8AEuQW3Wu4F0aQvwAtmJgoA/+r5AszDfFA55I6eY/o7ohnOYzNAAVaZ5xU0NpprcljacHoC0hu6
JY+iuOlO9Vj4X2U0p7p/7iekVV1pUMv3TJZ/6ZRBBiyREe02F6xUb89461DYyCuB10eEqjeOPCAM
QSb5JjhFFPSYcN9jA4WIOLjFQ5tbaS4HvVrtJYlJSHLnXBB8vICFAhE6fVMfT0TCACcYsvYaOmzD
r5sFKo1KXLdKb3eu2FoWxtRLHYlNZ0/kuOGlzk9teFPB9fOgCIbRRt4Mk0vKtzysUxuSC1uKg6NP
ekOsZkQEbk47RGWn9kE48YtS89CtXjKBgRUFmQDWVzsZrks6N+EwztfTWnqpAV3uKeKqiI5VwI5w
fITeS3DhelEFgFpUfhfdwIJXfTyA14bjUhp6nxcR1MmdFfj+DhD4Mbk5TNppFdQ2BHXxvnnBNiSG
lItQ4EgUy7nQ73wsrW7HCBMS8h0sG6r/SrAN5Xw+ptffsCOC3xFf8nKICtZFQV1t8pl1ABXf/Z/g
WaWGehFZktzgSJSKtdbFHLbgfIw5N7qP0qAqIHfvatjUvvdcy9WFV4q0CiX4fnST0Ch2kMZu9bVy
agcC9B7w9nRYm+syn0fRnOLX0xBu8nNl6b4Jp7CSMNNetRZ7ysQgeBwKO2aVpLUdOMbgVGoUxz6O
ECwbnLhegvJjIHqD42pVgpmaDvcBqYY3A9iZqypUqD50QAwS9G5vjTKrg48skWb7IZ99zIhp6QRg
xPmMucBebD4rsLYzaGccNSZHYslcvfBf1GGEATb2Ajklatgl3Wzm1v5Ok2UBQmVdH4IZpc4CB1Lv
Ep/Ox7KNzG+47nN5xlsffGLCcrtCvsbrEx3FvFxYHhrmsxGl1M/xjXCOKHxbaZzAHYf9gHI78AMW
9FcjMNoNFEv0EkkPNlVMBI6iNnmqm9Mctln1knxBYKna4pVUyAZlFBIrVPSED2XNnGQ0WbONydZd
Vtm4EDWzbcM74botw8EyuMcCZSS6DWI8WjBYjJfFBcv4nigXMjr3uh/XciM0o3Vq5SGtY16lEizH
REX2At+DlYHHu+wYMCiR5LmpgVviK6JzpYSSDVdDOE22LqDktVMyUBBDJwz7F5sfYnYSiJLGCii3
0fmYsfut8GdOxxY+4fQojDAYLWuOds92J8bW2vDurj8rJlR+cSjFNV+Uh3ZBznRApQMgncmnxTju
Cnf2aj0Vo7mgKc4mSswMtfewm/d6Puq4L4/eMp9dNhc3nQuh1cWUmDSIXp6CdYUC8TEvvKF0qonD
lJqiCdX/Wux44+vN6i8sAzedkdrq5uhUNctSxBQha3hFiC4snbjxlcGCiapf6sWcVnuVuyChSOYY
LK+sMbKf7QuEcGQc6Qmex3ZBEboTqjouztxrw5Al/bHs1hGRukH3Y7dYU9VaYILasgyW2XAFPXBM
2cN2iFMKZSz2MWQ9x+7GH2eIY3ZwCQc2r/wXHhO52BtYQJHCeKe6Iosi71DIIJEXCInJE5leSSyx
wlO3BucADe0TjzD3K60qiQXrruOrCetIc1bzSWhNfMXbp7HjbWGSYFhJizn2f1XOwAsfqOxF9bn1
wGvGyBxZUYPK8KG33bPI1a/Qthm0787mwZonULzDCxl66nbBEdsSdOabygTDUdhJimU7aEVf2iR3
dqsQRhQZV4a8DiW7cSa+IofejK7r2/EBOnh5h6XT0Ar+kMzeFWtV5v3kqDUpM2Rhn374N+2t0eV3
jrLtmu6RvYrESLrT3xE0hQP7b3/hIP6hW86NE82Ogq4hmQdzX7pWvR6/PDXtxN6C4gOAe7N72dKJ
bgfj40/uh3YWftvqepvOT+tMUM9Ve7UzLD+HB/Mn1VeEXaxTiejHlL431zsw/uZvLl4FDrczWq3e
pbCkJ41hpOGaY66G8twCli04T0IZHLLh5xwdow4uroU+brvUaUKDf8B8sI8FyziBzAaL2/QLhnRH
NXkFDV/3N0ZHC7rVv0faI7Bbrdw4Xg3ylfAR1HIHx5f0/9Moc8Cax8m7j30fQA2OovLzV/rOU+/4
VAaIRnH6O0z5LUhTF8BwvArLq2APg0a4mqfmmv1CQSJEjnpJeL+lE7J/5ELXUR06RgqySu0FHT4Q
XfiIQShTbJkA3/TQSRAGaHPWpBpe6MZpG6cTetWSGkhwUuSRMkoQxNvd4W17fzbLlyypdl8+OMUa
bi5Tqqm1pnrQG9bxJ1L/W4dcGSyxP6cj8csFGD1UrwoG7HgktxDRrOrNbR76tsPl4+OpTTNBTG58
KrND9oUgnMMTj7EW7BqKi8FnBDSS58enJ5qoD24+tfcGJGdEflOAPTb26WOZta+AQjVWg1T2m8Eh
Ypmfrd53FqDZXsba7jc++rjS0yp6hTvtbs1yY90cd7ac0yN5T7Xk+dWZfEnpKoiyQIkgUVtH6nuR
RZhGct6sljyimqJCj3wNusm1WV+8Hadz5UzlD/TrG3xdCw14hA9NcQCDH3YK52qmt3cpU/A1K5tB
w2YYUVWSK8BqPOzV9qe1KO8IeFQV3vIGTjTNqo6H7BMXFchnFyAcW1Y5L72FDmdaIaNix0pFqahK
qi35IdkOQEiLpruhVHPoKMH3sbhvXlbQFyYhp1WxVW7P5150WXtUQzp9YjEYVh1uGDm71IxEjGQh
S9CBaQwcbA9LzH0FlPs0yKtM+BpsStAmZYpWvVYxz/Dc3I72PDKwMTCLPM7lLO+mStHocwXDENdL
WX3GNJMBVlbkTR2GCvP9BdRQt8eg+ptK3xbs2pJdHKT+KyKaFF39B7qSRt82iUxbpmt7vLsC/b90
vlBAKq4RoDEfYMHju9MN2AybEQtfdZ6GX4XI8pBo2HorNDhltwHWVhYTXbyYRcwpADc6yehWBLhz
dgL6M8D54IaZYL6xG1KpNaKjf/2rLhW1BJ+YC/1vEJ2YyLX5/aCNjxeE6h4PK7/aznqGGVkS2J+H
WpmqD0tabXDcpX0ITNH83ytBaoAm2mvROHqYmR/6D3kGjWNTwkrtwdd5w8fWFvMyJunpJW/d4vVZ
JhN5Q57ftLbbQk5bJSmxQqW5UV+3jPFKjJVXJLbC5df8FukuLxeZ0CbYm7tydacDTK+6/EfhjhwB
3gop3wsWoBmPzsozuCBvP9FcLA0WPVVbAhaw0OxzS02m0lx2iuEM8o+H+R05gD8NUF7thvtBRS/I
gFcRUqcZnreHylCRY5koZsmURhv3K15rkCfY4LZFF9+1ucyHdr47u94y2jDlAYalRInfmFnnd0Qh
YA0sJn49PLxqnrGBiTry+gW4CIPfa2gT8xTmShzDsYtHoXwKjKQc1TqkQblknHUSIPzv8Kz5uvvE
wufdk+b+JxxiZBjDAxVJwklPqLNsDl4j3MoVkl0dER0EnB8RWohPrkrkFdXnk7pizQKMtnWVRLv8
+MutyHTt0A0vxSpCR32YmMAX9Jv5maixhLxSKT0S52u2H2iMLucWXaWGsI3IKisb5o3/1n2zEwZk
3qoCmyoZknteJt7Q39vjfNTmOz+8Voro1uQVzO34mSeV9u3FwFwiSproyqZT+EKQIs3/yfgBisDy
QxKb9zomVNp4SSLSzXiY0y8VdyPpZtaFcbITOJNWD/gKMTPC0KsLhgfDaMCQ8+Sq2V5ESc2YrNI0
Ts9RV5h88iHBY442V7bwECLydYKg+CXm0Or+EffHJPFK8PBEU0Xc0dqvj2bEQUZ6Ag2Ia9lgtHmQ
XgdFy4YwMr8uO9WTJNK4jdYZhRROv9YMMeogMmbTEgf7LQDxhg/FpFBRgEsdxZSdOTHfdKxrr9Fy
XsuXx+WseIPJ+aYYjGv+wqaHj81GBuQRU5EenPkl/yIcNmifejZlNVEqHDgtOdGjXCnoJXCzd57O
lyz53lkSfVcN4H5K0QMnB8TW+cgGPPCJ3u2Jzfs6MSXA1jHWMZs4ESBH/ohhEB7NsgCQu+WPXvKR
14fc9FKAqVK7F5Lf2QkAG/H5vBSLkHlBLGa6hs3olDBmqFhivACr5XqStWvlS/tH5mlx4IcKsgjF
Ghx8LuRHTZB8nnrw0QZlH3IKZHTKflLurHIaB3tb/g7wEy3zrBE61Y1gaxiOcWpKuw7S8N9afYi/
a85ZQVfhu1SifcTFlHbL0/sKRJZt1jm5PFxWo84/YK90Y1hpCGlKVplbNtQG1o67qjNQDZaZZrlx
H1s2Lm6h5djXgqZi/KjARNguSaEHWgnCYUYiFVzguRJzZi4Fnc86FgUYOscRMoawymSmtn4A5p1N
punuo6J3lj5Y6/A35BcXoHqN1XtdX6X7f/xNWxwIj/qMhAwQeaBN7a24r8J4ZNBP4bcIeoNac/pU
qgsZPehIl3d9BcIk/aXZl2Fo7dXT+2rZqlKAGgsvySKf82wyP31psvSvsrobpc9KE4WA7+nZuQwj
A35aErccoAxy4WuHEi/Me8szP07TRzwW/qYQNeDVDTokPuVLT/NAyQS+bHpwV9gMK7YZWGZbJ+Cr
29EJjEqaDpohI7aKyN71PVnO+WkJQlQ9OTaCeGDzTbbYAkty+IZfRBJIrTOn5mKTMjLjLk5oCFnX
GnQfa7mDC4yCBpW0l+YPGKzUf7uZbOEF1LzeWsuw1j8PTN0zo/6mPoiMiLm2fnO2DijSSYxv0nPD
awWhrj/DDotr3uPfOknQRdaOkmVUejmz1qvcQuh1AC39DibGwD/OnNeTEDCTEsY7uPQ+iYSjeC5n
fWwXKfWDmSGAMPcCtODNXPy87IOUPJVjTPttgUxGELBnZqbYlVNdiRUuCFmcRyzUupfl4CQVk56+
iUoxtkHoPxXIQ5RxkGnEZ8dEV1/xoNVaETP1NH03k7o9JcYwO3irIhX722JYgFQzVR3YwL/d7ux9
W/wmIKf7xuWKQkT5duPR3kWxZdQkNI1Nz02BId0yB9tVmbM2LjTSSvSR+4uf2zYaeGM4xkkqVYJv
zwLT5BgvmNwQOv+nxULWHi+lZWP+ardjAFmVzV2UKD46iFyAWcLGtBQHEupqYGP+Uwxpzll/69wd
mfGa7jXjYblmaMz0NnFPMB+KulN50uL3PZ2JfPKF73dSK5I7qdQDoIOiEzFB9lF1yAFyMJMFuFQd
SZx7zENdEF9HXzYCJAgQjrsL7LMoDE3EAVvK52O0XCHjVl2NFzRwQ+jAqT2lIhV/Su60BNMI7n+R
Yg0vLju7/s5B/FFSLydWZ4YjCB6fUjC0tnI5KHxSlNvUQkbNqhXATzGw/hp3CofId/auhdYXjSuB
Et5MsjW6D4/dNU7ng5CkgUgXKCKh3tDF2RApy1yfPlKGdseQYAc5kqdKuvjBXfCf3Ju4NzRwvQzG
XvNM6l0JnussAApyXFJo6VDF1C3/3aWzZ0NiT+R8O3ig+0ofIdv11P4/jzjyVNENacTGQ2rE9+Z9
4JJRVJyVXZ2oTGQEbBMi7kgV0td59QSc30Se4UC/lvZg45fWdnp6WbjNQQag0zMvb5cvzJej1WE1
qKo5OTaZpQVWk9hDy1qsBeFnHZKAJGsxoS4wPPIfpJpEHzJlPgChHvObx263CJxzOGrxlVOTuOLw
G3tEMYxY3IXxgLDtK4JFZVINUVsPqG7Vgg+R8wMuxBuG5IpZiDU3nl7BWcN6J8p+OiAA0YMC7bxO
zup0F35CEk+QSJKEczIX+9/CIiSQkHWT3u5HecyonI9OtF5T4sFh6InJhDi6h3rVtdIS6Htv2J8j
hKl5AesOxwFbYFc4YW+pV/uBVmrETBCe+ep+jpKQG0bES1Qagz5COqbH+9H0MH2ZUgG09b/awpUJ
2UtSkLQFZPQyEHa7g497oGf7en0JPp0/xFQSz65OWftmtPeArV6UXc3AicCPgfmyJNsEPVkTmywy
iJJX6VcqfV0p/TkF9+wE/ZhmksQ7S5aPp/je00Zo0vEKZVafclqNXqeUga3RPUyq0QLsP2b/k5M4
qnNFcAsCodFbs7upK01llY8HViObXwBitoHRc1vfadYbSpZCNg3PrXn+Y244q4LgvVTZJLtDW1CY
aMI9WGr0Fs3DkzrghxiRZnir2eUeyu7IrNJ9ho9GERT+d+ZmIU7HMgPBzyeJaGe5q24dNfKOfTSs
S8eH4DWvJcaYSJxzgGqm7YxsNDiq+0KVniRI2PnDErlBcx/8SoUQf2eNAxKe0RAhGzunCiRtDcRk
iUDZHto8wlrHDy/ZWEQa56l2zu+B60zTk4H1CeGVfzbPrCkGekMSU+XM+94zWaFq2sCaEDhT4kW0
2f43d9xfmCmGbwu0khDMwBKwiHL7lIrjgKAuDWwUet05DuFsSMzvNzZH9MW4NLZHsqcnaaxuJb6n
HVhzVyJZGvYTLsFoVsSxzh+dx4WP9SLpQ0ugmlZq6auGLZBDBPWQUSvcUytwML4ZWdyFtt3kaNGk
bRHCZx7Eq7vGrYIK7mrwnW/CwAS0QSKfX40Eb4UeQAhtSe5aYazw08SVPRZOBqiRiLB+KLametzy
N6jb68ofwOf2iz/QHpHh90JhZy3PccpQocLFg8vbIIKDcEXM9OGQQc1lIzsVjgZeDbaPpDUtVGMO
PBtOGTBH9YYY97jpUP1TNOovL+ZEgIJN5ScbG2fStvI5dE5YxkEN6lzaxJapTXYRxFTLiJmmBpEQ
L99CpnHf0ip4kNnI0g+A1YM1xqlKhyjzppNHA76hnyZbU22YrsNxq5xTu+aDnDFxOQPSvBmy2ejO
FX4HarGT/ygwCQX8EMrEgdHI7w3ZUQpjcUIjxnq0utoIxKcLF4p7QVU69h39Idnenxt4SEznAV0i
vzfk0NAZShXLD/OIUHhlcws/Qz/zPr4AEDYz9L4gIGbo+KN0pseKW6UN8YZri8UC6Lt6iTEbfEwx
nfbqWqRfgpl/OQfTr8UyU8sO++Fm1bOYQ0Dd3wTttEsdUzkhNxBA0CvN+eCrFFb+WLu0wwxD+Bot
YdwpMvApNzyQ4+1TISfyVV80f6eZm8Jy+AAigeAVkQDR2PZhUU3dpXcCX29CpUVZGvsrYtUjwwbu
mmGDcYJcy2y4dS78N8zDTKXlk7nwRnTq51V8kF2Oe0bSQrt1SAVbQb+dUGezVdFJA6/Ny+7BYFC1
LmU6PDVaU5cLcRfgaPQv3Lrl4cayso2sNMnVpgh4RR2K8sbzL4gIlYz1MnW0dNxQFKhxJbep2ABS
wR7agiklkw09XMi4xhSk6pmhtT12Xe0tLvDitMpuWeoaZffs/r1ArGTMkeYLvtAxXVvv4BKXlC8W
69UR0EqfCWEXJjVn8OD63Y5Te2JIjAj1ySMnB5cZZ30GSZ8htKjH62/Z4KbCCGA+NRQR0cQUPwcU
NevJPtx+84V3nGSwGaDK5WRjX6nDemMDX8LSJ4p8/NicTIoQpMXGO+A/4W8SGcnJ3PLfkzKoxS85
+47j+S4PyQ+RooQEeN+nhQETHHu1WKJeRqtKhzVfZ2vzwEOiKczuLZhCyx/jdsmQ2ojbuVdKcvV3
0iN8aeuwmVgj3Wlklo+d1Mu4tsIqal7f6uOKhnDRBY5IP57jX0LAhiExCAIAuq4ItGTDUA16lZIV
v63qEqIwHB+PNoG/wKSOgzEH3La7c6gP+O7QL+WQ+UZEh++fAWVn/LpW2A5odXUMgmOE/9jYkUFV
cXXXJ3Crz/dLaTy697L8ZJGyA/lzDgu6HDLPuDZ5xQpcZw/M/1SxP0nUJ4XmMANEhuSA9a2QAkth
ajoK9cF4tiCw68gaF8vBcUK7V9WQHcuhvipotAraSt7PDjnx2I0R5PuJ7h+E4KJVQhpy6R4LXMCm
m5BwnNuQfttKFiJHGioWok85RxqwzwMJDvLWXJ9HPJCNjjomd3pIaIwdN3RoghdBSmwpLdrwI53L
xCYU25abkiDWMa1wla3aEYXO4J/AaqDd+tSLe9JQYahKp6kKXWHrEXLkQJlOc6zFmBtuzEHUi0XQ
duNVGZ+i5DVrU0Q9QgpPebpsqh4MDfcNAWFUS9lcuWBVm9bdqR0yDXXs53jRd3USjGDD2TEgm3k3
EHe/Kt9r3w8NHrzKRkknqayR8/95kPZzPdrScLqBXUSk5E5zR6aAdoDeLXv8bv3t+SZ++SlzWGz0
eAd/8XTmFMMVxMoAP1Ids1XjmNIng1fOtGsFp3v06Dqyzj03kZVdsrk7prieqY4w3aEbGh/H0btN
CVwWx8MOYMsklkCckdB7gs0q98nKU25oGcmEBrt7tZ8t0i4r2B/+B5tUuN+//DI1zHKsNce1IIAD
w3rT+PrlgNYesDJ7f4Hb3vuKwRXl3+CaDWwRdHgiGypGs96TVwkx4UleUts2m5g+1Wo8QeuuE6bw
c3SvDOciyo2fzLwk5kqx4i28V5854me8qaqGfLv1BfhKacR27hQcXTZKz6MY1p+pU6yVMNvTN51W
pelVly8At+PE9ArXBhFiAM9o40VdsIaUDjU03ElXF0Lz2thBnaEMfkUrp71n56ZHC+tSVV+v8Bsm
PCQbfvi2++n91QONh086ROfLf7ajgrl7SuTZ46EUtD+XZLv1Qrifa4NEIIgZbLIwhW8a+3eGHKO/
tu7lznY2+20IJUIwoCjjBMGhvrZ9FX3MUmvUq0j6hnQ8cbfRTV5pi038/N8GHUBeygtdZ7mOLAVH
8j3UU5zIXzlQe4cWieR6fUhhyV1BmUatGjc8RkXjrFmk2/kTMKVBQhZdIelh2enqRXfz/tC4GOOW
Al+05LvdpS3OOhM9FlLNWg44gZL2vJ+/cD102xq+DQu2cQZeio45mdygGF0N9IIuXK19kh4IBWSU
+zklY4Jjr1Y0B6eqkwAj5SUnL0KObkI2v7q5YCcxl1SYoUONxgDElmDpUSkHCEhrZuyqrmh2AoTK
zscTxo+65hPclUi7XOwI3ZwlX94/Yo5uQmUpYqXlmZ9IczieSX0k+EdlpYYGC08VizM78FhsPmhj
dr/eEii+z4IxWAQoNOohD5uRh00oTJjmZhxVG3r++f3DQvO/SZIsXXWaVf7FadD4ZRmkterfgf6h
U/Sa5Bj/X/gifNh2OGIGYk1QrLy3Qbe+rMmV00KgLR1uFOevZ0XI4cB2JmCK3j7QiV811PuneqTL
hhEpAmic8jipfAgoSqv5zIQD6l4U2qYG1b198w4c9hHCZGS5oNeZpQgn4t1LiHTkechRgU32gAOw
2ZH03x2xxu4TX+LsadF8aRq0FFtQ/hw4xocEzClHUvFQhjbMT8TYhXE5tliciatD1OaI8u19sfeO
2kfE/aJgkWieILHnckDyhQtesjxb0KKTG7kdBL0r+KXB/w+AvbF6IdtuRt5X9cUtusiYndPhMMLi
J61MMz6kykCICm/hbx4+c8iK93BPmHnpNooAwNUx9XWC5aNVB4NbDKGQ/gTf9zYlgekbnRyWJCvV
00yPvTAjicU/K/IQ4KmopujLzuYL/CXrZQ6Qi2HTMCXC8rfJQT7e4HRcsbI1mkxbua+smtnhtyRA
mArJiOFrH6NWu1ETmh9K788kjHvMFckw0k0LDC9pkK2BvgOeem05L7yGpgTn5SjLymERSQC0QIm/
3bTPAsfUEYAKkDTIJVJY94GW+QabPByueprjgPRgPROLa7b8sqBCTGC8M3qCn/oriI2pYBLFoupx
Eq1sN4Fm6zDsz/52u/HKUyQeHhXEQTDgojdG5mF2igipWDwU4KkyI/s26dExU6XhLepkjFehPWKd
2B63Lri2Jn0QEGjqpAZ8ZvAk9UTVWsUS17xz7GCh0ufWJTt+SK0pJNz5rUgM4+RuJk4zamtJUeY2
wq1uEaCMexD59Mi7PSpDIsPBurlxYA+M2jao5C1hT0O2WX12VvQoySOYlqJi0R/Jsjl3HCrmtWta
ZHCxqJdF3eFXJc7WG/ckldOo81erR8zNLzE+IblRHCsbdCJwcRwJ3kScUuGq7ec9kBwxogWJdsBk
WmUbrgoc0KrgdsupF/goT+GXgLSZtTpBbPT98Ow8GEZ0VgqeMPx5yoQojL4Ze+aKJQIcXS4WelEH
fEtj4whXSkVWrapngwe0fSmM7/K9iUn4CiT0ZW8Ey2kDUyTjCrBwvWo01sATmBhd7scrVG6p6rF6
mIaZmz9BiQymdS0dOj/tQcgyQVYH55qZx8WcS23Z543c2RrNbNe4snlU5rDSrKDTArxvfBb9PUul
2BDF/1AXhXZUyZ9cBfF4Eb9iiTELcZ0AVpNLlx2PUoUi8QeUKskXFtnH5EXRv7Ue8+ZVD7Mq3BIt
d+x99ZL2FQ3pivot70xHEngwpKpBh+iX3KMjgZgXMd5i1GzTtUUYXE66tiVBS7z+1OmDiALYEJk6
CwBghnlLEvx+CEAL2k93CKw5uSND1VE5LwyG4Kg7NQFirZQhb3KomdCWnLdJ4aOIp/L8a4aKun5g
w6Of8IrYV147TOw0cih4YAUbay8hFFNuZsHPOYn+N+bfc25xEuknURRzpf4zJeW4gWrUFODqRzZQ
qvS1GvzeMHPRPGAFFHLk/yGeUZ28AAKFrpPs8H28j1NfRI5rxl9q3PUf2AbmZl5a6aC6Jtj68QrH
Er8ibsi7VgfbBMOKcosZ9DhOFir0v136LS2nA4nye898Ssc3NkuNpRbmU0Sf3cmdFBkAj0IfjlxE
FFmZ/6+JqWk+SZHP+7iHmL3lXrIKbky03eH2BwZajmrCdf+A4Sjty/+mcb+c3TWmqE0z3xGYNNkg
1cZ3Em5PINL4UWUZ3ZscPY8wNLn/CidzyVB7WU6krFAa9RA6ydMeUaBKyfQAELMbBFJ7DQwQgXMg
X376xwZiUbSRya8ihXvmfr9qFUd4o0YXIbdOUWdqMn+cDwx4GmBGrZzV+0xdB1WGOvfstV5++694
M1+B22oFrV7+NGzFUfDvR17xM8e9FLcEOW5p31MJ2cj8tlzPEa86gruOPsGW2HHNPdoAF/NEfbU2
ZGrRjxMUGYGKmy0Nq5Vr6C070aB+yR9je9/gP+8JIMEUH7J3yBbDYFwNHcAaSmOaKOY3TV/mnbGz
5wZEhOegTawcMjIZIIQKHHI1qeJCKvSIMcWo3Scsi9t5paMJgGksIbdksOBm/K8Kn/qrIzu5fJ0Q
A2sVNUsPTWxpIBNxSY3yAX7g2Qb4omWSD6cqI+kX85nOgYdQ5BH5R50qKsPBJo4sksbMnQe1Aiao
4ce6q4Gw6VqnjEI7JdFHsDhTK/0p3pdBqJZblIQq9wum3nsnU4EvfcBnWFMIoiq2e5ZCBuVGRYnu
3XN2l1i8hgv0Er63znvkxUmSe062SWBfLkePyJO/HozB2cw92ip/1eZNvU76tDrYA/C6gDzi23YG
PLittPOlC8vFksx4ztMGZsiGoKrDC9UQBzYRQtTIsI9zsYKFB4XVNwH/awcaxOGKu0ivz6fxdyVD
RqN6Ru5A40tjyfB3e6aWz03pyhtYfdKIcqRGs7KU5XBGCPiMMJpTPiSMXQKF8cccd1Pce41lEKfx
OKb0H0y3yn1V7XWwZCwmZYrG69ZGFslC1tgSuRrBoHYNcwbLRwXqX1Sq5bQ8+6kQQLffGkyQB5Oj
ft1Hs2CU0IuNyy+i2WOgW2bKfbiIMcJHh0bxh4sFlPbNt06yfIztQwfyTd9X1IgCVt1aZc76WHXT
5x3oEKeaLfmagVpZQ/GLzy2yv2lF4vIGIuYqvBg8gqm00sJlGFJjYLtgnLJdt44uczKuhYCVkHbV
zrUfUYC4KNq5YhiYkOzmVt4I5nD34y2SFHjkyzuRNYH6bZ0pv2Nvw0lrwaPcJxWZRNwtJ3g0lsFg
8BmtJPo61FK0xOAn+w1CMF0o2iHzd6c+9n5O3Vjap4VN3bGIZtVqwYd/d6gYx7k1Y68yG3lfwOK3
f0Pt1JvxvzMVHvzA3ebk0YVon85lT33aK+1AanXt3GJxit4dTNT2tF+/E/KXkrCtRFfcZd7zzjE2
hT0QmPqGdz5wAUliEohj/IOnmH/+TzU4svsEQg7znR6bisFs75qVnWvv1/VPLyThzhaSILu9gTPU
0tJ1jUNAgi++7ET/rlVmap91epx/BYhCVvY/HEr8nJx0DHjKUOKaTOuJqp9hhfU4NAi+8ciTbcHY
/h5Z68b2uwIkM2sZLBKEE9f5NsN+tEELNJaRu5q0jC0Po+QBtJjOEKy1zhwHMFbFLCOZZ2IfWbxO
9f64Ca2LBVa0wDv0jHiJNDlFSqxx93fpBMgmRf/38B1n0HiG76omjkaH9ImY+5q+1g5nuklgUIt8
hlJj5KZtSExEdTdBcTRIMit2+SUDINv9ABijPj0nQXcyPLPtseVb1uiy9CPXHQdJ0vDgLZvouPb+
RYWGBF9+fhrF6qbBbz+oIAQEY5FmKNkYo51qr/ClFpHtOLZ7drMzr4vXmSSTeau4WYIzN3IHRyqV
rhLeUGyfgAuIaEv/rQCZUILRQu6YGO4vzdXc654E9JpgaGhHMji3mz6Hs0mGsIJ7UG3JewWHs/FS
MSP2iBKFDSgpIj52T5zze7DY1ZmZ12TBsjdJXLjK0WHW7JXKsuAUR+1etxVPeLpXBWfnl4ym7VHO
K0eo7WF/r1MF23bX3I3ciFeGOiyUD+zkKbtV/7OjAGMOjqeK1sITtTr40NSRRjOQQgmPGqkTYmRW
S7n4Ss4qJjOlkcRYxRMOIlxRiNLjIkc158Sw8jBauDS3MKbhycCHLP90cB+khA9u2fC0VmqybvbA
rf53g9ZgMjmdqsQKmd59DY7V4HmVpbzpChcmG03oPAMuHTZDOEmAC5tHyPGDPDzbSLbHjwor5zTL
YVVLKULpG1OmysH8GTaN69N/Y0EqS6UJFHNCU/NEzCd11aP/EhDWGTinugrMllhGmKQtHayHaOWM
bG8FVx4O6cHraOA1AwsGsitzwEHHsjDSLe7luemCNnLKRbevZPEKujmmhq3pGyKyZQfkLj0L0Ocx
8ZYY2Nz6xNBG+hNjh/L3GHpWRtwBz0YPRHCqAixhmehwfUk5m3t56OBlY80yNcVtGSiV3MITT7Ta
RpLev9g27ZRTfwcWA2jQWgCU3nBZC7UBz0ZiG1XVzCFOqn8xGZK+wKVq0KEQEdR46j4O6igswRHD
QpfAqhKNOSqMwkthugidiI6R0zmnQl0BkY72C4iaM6mIVdQ3BghOhXiyOn3ZLR+g015rmeavdv2F
Gn15eN/tIp4wst245Cgv66G+XSZgVW1+iVvu4FIL/xcPbBJ8G54h1dueTiF6K8kBhzYq3/ZUY6ec
DjSi2JA1wugmObmldLo1w9KEWSkZT0a1Ln8l1Fo+Ofjq5vi49XKhzGI1WZieYoDVypMzk5Pn/XOo
Z6fmjvu27qQ1COzW/HPdglL9NNzA8HvI+/4LVWdcZisEGXwdySo1GZcexL7MENHliZyAhnwjgdu4
KoWzpCZycRUQc7SmBSJUGiFpr52mtjjMn8wH4fzcvlTcHIzMef9w0V2y03aj0HOoSkRgGnEzNq6F
QfpP4VkksklmxqBxJ8SyoogPILuE9L8D/SdPd2ihrBvrPcpxrTXqbdVM1EDfCiStRtVbKt4T33IY
TJSc1MlCGZae0SOQTkFgQQDVhCAxg/OGeGYjN7o1u5t1+lLYydscQR97mE6o8E0CD9/M8aVs269p
/ExEwRnBs5PqRH7xFlc2eZFpKxK+9K9Qpq+t4BPKJYTwiepC92y/vbJxhlMwjh9+L68xwPCxBbis
9Q5//G5iAc8FuA+7mBSqML1liPcL0HLrS3xaVPx2lJmibcguAxm8ooBrNEBc1O18cvLxw9w/1hmC
3w7Nx6JhZlu1C0L0OEojPQb9RhCgkS1IpAjKdpzrXbV+I079dOk8gfT9exyi8Lcok6otMDpQzp2N
A8lCiOAQXkn2qoewSclwqYdSraeOur7POdadCLhPZ8h+wWy761ZPdA8wDPIJRvP8UAGDlnjK5rYe
cIdHvbJo+g0bxegA7v2xA4bz8wU7pnyFKNg0TiFY3lvMSEFh/bV5RvvdwwnycszvWgUTQ/bs6nJA
zkZ/sytQ1oCszTtE7A2B9ARLCxha186fP0gJztbVHpsgcvVYp/rzwBMVgZxCG4ex6T5YH7fHGdZF
/xtMhc2r3OG24Ac9EWpIzDfFjetJVfXC/+vEd7cEP2HV3MfAbXGdQDpsR/1ZyP3QnBkKCDJYDJUb
3XChNVJoH1HwRjIkEqWHAtpQ1PQnNsJM5Owpjuma3/f6JtXsQ69moBeQCCDuxTRkoZ7tvdKxbJzO
surcQcP6cq9Atv2pfTZOnDPZ9TKLb3WRRKArlaQYeY8NYBAGY9IACbVA/6e48pZ3gRtG02Z97jD8
jGGdsGS/dVX1/2IMNtK3rrkcSKP4fL2b4/Z3jr7DeGlEWZn5MissDmHChh0jYXlvTit6qFqgiRA9
FCvzjkf+p0hDCzzYNy/6xi9rl+yzelwD1OWeoyojF/pSxQK5YiVc2RIuMIfX/5Pnyw7D+cfW8yRf
ARn7uZ344E0HToe3t9G+PBYXoEwQlRNdu46OFQBd18F90/ghdbmxm43c2QpDIQQLHqdzVDztpbiy
nxZBVCJrt5+Rur5fOW9Ky1f9a6tCsHtTV3FeFRpsBdbKy86cFlHCGsCgESRdC7SqX7fUmt2D0ihS
6LqMO2RYB9P3D3qzaJm5PXzMd9K83sx7Q34xPKs+4j3BqYsXP6pat91/7rwoOHS5uHQZ+GzRqzRB
xLTjP7QJmezXlkXvZgiTydWhlrK2TpLCY2C0NkozfrM5OsvWCSGEojEXg6j6Qx2qBMdIANo+F/FS
4cucqd1aepefLPt+Of//orMacKYgMkJrV2PqIwTTuD6URx+rrrvbTMiGy67oS+ge9t9Y5lczyyRX
adb3zLROx57Pkm74lAyZDo8rPU/BEhazNXctvoKI67sQww048tOJ4RXhjyf3U+gGfGAsGOzUfNc+
68on1VVsa1/4wCgysXusvkdMvAdaoafIEZmTu5QUpY5tkq8EmtS9LfhPvVBwmyMKvV5zNY7twSNH
Nzjfoo1e7Gy4cdq5gj+dW5uclKcMZheopY8wEIlLj9Km+zGgaO+QdEQTYn3LTK2ClGw1Encdt4nf
bYWanAS8RLokGNVS2064ZxEIEVp1f0HVKir2dakVLYBQsVoOvAQjgVeRz6R7ZFFVwX03hZTSan6D
AOVX0bD11C5B7lNBlAiHgwcHmeuWRrQGe9n2XXIXvBo71x+lSONzZ9ntal99vMaGL9hiE/14T4ii
PzD9R+08IrcwLrcj0ypXABg2A8ZeUSqy5w/oOKp7+h+gXkLGoH1dVkA4YMcq68GYyxJjtIHIFBzE
HtQk+8dghcIzgA1H1RBq9rwmAb8GO+N6LBMc+scSB8v7Hl/JL4ZT+xRCw0+VXR6C2A1A6f04mqDT
ivKNuru7W0JD+TZZqZ9o9ud6caKwu9TuXJSAPzlSQJUoNQMOm0KOQEzhH+Lt7ETp4a+MaB/i7XKI
q5Xj2GVEW+ReeKFcDFGeSM2hAMlbT/SuQEeSIVE0iZqbvLDOJhas+628ZSXuHzZZrG1s6I5FJla/
qN/+x8Sb7n6NOzZMTIoYAK9bA90mS9O1LCC5hYxbFHrJDcIpjhG58DLPV83UqdqnI3UAyVBbTREK
RbpobEL+NY4PcxmHEyzAk96dNLU5BKwTPVb/+MqOuzKQfamHDyP53FblKLgi1zQ24Qz247y18apJ
vFGOtI3UDdl9V2+1sarN+PWnwx0RS7vJQas4btS2WNg2VdMo0AdSzKKnRScMgFyAoNZXHyfJNAgA
5fpBwytQJOAvdtxXeMaCbch7jcSiIxyeEUpp9kDQZgBMnmEslAou3nGRGsjl6TdIfl4c9VKtq8yE
u+7Al51PF5LIuRRtXF/4KE+DFOXlrCMp7VgbYM4HpCQ+gYCy0v2H3qIlnBiJEsnfQiJoYam6jTdj
ORv6J6e20zINq7ApNoMohabNHvYyzHou2Om8KpwpA0zYdPZ1kQ8SV6WReml0FWbdQAAZiz1zHCoo
++xpx8sI4UWALdqcpkpEoyYHMLzCCyQi+61xxyJyNPd1QEqlr/6GNiB7bB14LJymAS+ho4pCQksy
eeMYga6Mm351uobFLxJh3LHOpDV/hTy5b+SGKGdvoh3//9kpBjWHq/E/eP2NPKGP7kBjbHKOvefz
hanJW49RfLL7BhG4EgEIfHUWLmNmXUjVFbDqFALnppQBoBX0ZLsXzNHPBfeX+aTlirPTCCmiE6BD
mfSlEEvFO7/5HWE/0vwbMdWjjLqVIDKtUO2WZy1EjZJ9cOqjtGgfr0gsAGl+yTifOIVqcyb+yOV3
87RUK5jYhY+v4l15MZotaZ0ZhdLPiQMmMBwE0S4nMk6QzFUjJhCjFHzngC9uUHI0lzIlmjl1DUL9
9+55YApFRVvIjzgPv3sCN6eKsJ/NGeoYMWgz0WWkrRrkZ1h/xEpbB03IqCZ03bvAUAtgDHgnSAMY
QTE4fWDsqiKlcnSBu23r3rXxGR+E4Ork/gKkzzb5Sxeu4O/mERycYzEXLBKbsFeCV3GmBU90zx9a
GCJQplePy0RMFbduyillS7+AajlXtp33OLezxuRY2D5oDrp15XGC9yWaILWSLB4+uPUaDeZyFkX+
cYNmxd3DH9Kh09QfqXUiuaLsC3cPzodm14ucyvCNG7yt6yx0bo3KCmAhw8JqVOC+iBV8AXFpRzYi
29HmYM9XY1zhw6iRTtdY3sEA6X9UIlvLQcuBf7EYrVfoLKc8t4wE6YSDKIIlCtEq14OyVqFNCrdc
1dNf9i6zxpsVz99RZLfn/ch889MMAlzbwugZSEGiFPPbHudy6WyM3d/tnvgIjvQ8NSffX9n0ZWLs
B/iH69vnYXcZz4tISkyMRTVeFYO4SLZOODQvsAW7OzRhyP1oWEC8ZYlk3u7P8CYCnh4OgIZL2XLj
TmGYbK4YvwdASnmmNUWqdLlnRpKkc6WXkaQjN3YZv9B5UsPoUv+OHlYNw3bhclcQGY8N53vmNhrO
G3skU24NCv4R0niBWBUl9kuS1aItBXigAyFVGU0iXTYr/kxeoJ5g2PTPjZ2AE7jBkWuuR6mRExHR
EP4d9Tt0MpJTi5cio0EGqM9rZAu44kurxS6TCmdwKa5XUoaXtrzLLe+4NAvOVyCOCi8X2G3Syh6W
ZPEkpSva5JSuUQWw/eqxipYQ7u69aERrGgjXmBBTaRnQ/RO0O8yuGVPzAXRuZtbDns+qfsOyp8ZX
IP37yiLMKXschvrhEue7D4vLf/bjSFWZzmGMmk0lFl34GV9CjXrBll5VJ3s5zF9mSs+cEIfu0GVw
8YgwoP8xGm6zZpVMep2UHn7/da+YXqWLp4MR1uLYqqcsRgxHkFLllsy8qPG3UbHfdyiuqLZpCdzS
xx3S6a5wkw4DgUhZxXUXO6cxHIgExwsdD+00TlcShQZutrS24BOKjW+GR57QkMhUCZNMIxOwqhzG
D++jdsRP1HMGe1K32Y6fv62F4soS5b+ntr7t2yszLbVX6IMD/3FxT+fFbOj8dGZ93vl4FmXrcdT0
lXL8jgq62CknsT56NDDcc+oY7wMv7BpjNT6+FhSfhJvGRpgkSaSTqPwYmIb4nL2aIMgD9nBr7t+R
Gh13WxiNM9g4nFAQzhCmL3dTp08pWB9CX2N7qJMDs6Q4JBnBOHaz7UBwSiYHgdDRTiJYotBRU523
fV2hsSiFSpJYS2u+sUnUGd4Mohfxsc9hy30nRY4r1mz2p8bWiUDvKY/PRMThf/WuSkkHJFAAj36r
lIAky3TAHDIF6/BUDA3ueMuB6wOetGsloxdyS9ZIJhzIBsXMNZtBCdjhWUiYJqAQBGwgHcCmOtYZ
s1YWdcxTrgvlE2F9LDKItv+YifevcYcdR09vCffLGxwFoTe7jROXAmezA/h6zISwfLTwGmcBmbbs
4bYKkBFYCY5SCwgAU2kxoA/9pjKG57aa/NN/aUZmN000JlEjGDIu0h1p1Y94z2somrsDHEXCYVXS
rXf9yQ9GyD1u8XxhJBOykv1p/blVtv8VZkz8fCrGahq8YWI822trMAg9cEz0YnRzWkmPJfJkNMDb
rYSJxFiaJRN0vQ/aW1JBg03DZ9N4Efty6O2CACTnXigKu+KloZofvmm7FDXXO2Q0DW33Y+MazVSs
6ivCI2J0KFENOyuOlW7fYoTlumHhHW53WA7bkMOo8CW4zlJfznFMT0V8NMVazrydlOWXEvLKWmtl
7HUDcbmuG8QYn4noFtzoTBZmmsJdXI0g7SNP6uE7XNnODgY5ta4L2YMn95tcT5RgfUw7H3/PXmdv
GtOVnWBB+FGHgXwmYa0KYptuj6bc4W2MXQzVuXssfJqkaaER9AcNjqO6frPGHoF7pXTlnd8bzcHV
QWb19sKEiLRHj/Klu3VjHCO8VwILe3bt2Erga3PQsBIS86FUUs/hq/wtUtXPt4KXNaQqAp0GoF7n
Ym1GbPjWokK9Nql4I4ZXmTWO6Vh4SvyHne1S4/SpZImNiZiMQ4NfA6E2LI9Vlg13fBbrJEXi2Tb1
XPXylUrzUEumAjc/c/OpcpLr77iIzx5z+wc6GDnL3deShVHnNB2Rracnt1jOLN8FAboZEqxNIvi/
yQQBfN+n7aMq5uJ7CrXsZU90m/BQQpfg/bt9+we0h6XFCEsXAvaJu2CmcBNxvM7oUPc9/lxLdOFh
3tcqdiV5F1qMHpJu/sq5SbwUw8/7gEfMAewWRKkDaVQe5rRT22C8SGZDvt6itBhEiJWqm+h8sjde
J5vikKp1Cnn8yWqtYxlwiAnSx5/6gfUNbmnyKLWkm005nv4dk8kBynwUBF5dZYAnqmN2yZ170ZGQ
OpeV30HHt0Oin7mTzPvpH58NjcsBApVfBXRklplPbVEwUSNOZYbmbEVqom2r+qs/SXzD3ONYq9D3
PWm6Ny42vZnuMiUN6MTfrIHWBnQa/FHJnt6MEAGVPqth3g+OqRS/Efw4qSsLfc/X/r4j7DqhzqIz
n5VOu5vQdjZCAuIPTx9nWoqYXtVkj2PqaDGNTS7SsFhKOim1VxVD1f5Bla2SgBDfEKjxkpwzq3bh
AAy22vSEs7Ahok4GniYJtsJfKJfRof+Cd5vh3I3KunkFmYavZ8aQmNWm29FGLDO/eVu/1SQGgmaP
FhdhHayfCUr83g47fS5AATqDv3Q/UzBRNL4S4YdKSeObpUFPg338W0ROesRcPblkfNG9E8U9tbzZ
+2XGWmnygzIR7+t31GoeW2OMaUw3QhB+jCAkfzUpSHhftp4fJevV6ByOTTPcxp2OHuwY5bsBmJNZ
j84KaIMbTB+bqAFVQVs5aO9mm1N6r8h+NdVatZobUex3facWi9HcC1fBR6iAMRj8N20KLcZc3J/K
1RndfD8/G7j3v2y08JYm/lD1TiuDM6kB+vE5hZ5Ce/+CCyYKFv+8y21Ex0X5wM7lDyYlR4HetATL
We774xxOg703dhbb1iPjTagMfGzMGlxqY+X8s9RuH3+TOxjww5UXqzTWBFW5yeprmItagu6dlkXP
0Xjv5yPvxgq8fDqzkbGOcAvHyk0B6n/ebNFshNeEaPOj6wNaEvlAZkOVMOMQknrckI2gwhwgSQ/9
ejYaWCjnduqqpWLhJKZChiWatzuC6neZp4vgGQ9iZMCsvKT1E3IR0oeIl7+9taAE/gRIKpowqfeG
W0jVDVlVemVK3iTrXg2qztp1dxk9BVoBDtPPDnjGDesCAwRWfsRCloid7kS4mzKs+sZgDNE9OJG5
cA11/XIJqeOL+OKtwrPOGer2/G+3k3/hpOaWXZArkH/quAk3uzx/l2idrdItSunSRNy+Li4papt5
BrD2N44sok8eLr5ex6GxP15NOxGhoAQnQNsvdY7QJjTh/C06cEAqpTIUnRwCJMAK0Bh3fMH/GX6b
P5MPbuMeJ92kWlqNT19IzhFWi5PwAXURnATjaqJN8Z1rebxgwLfuzyKomwcpoResfE/bg0pdQSp2
B2soZe2xvmZYLY0nZgNcYEK9ixB45lOOq+iNkbP0LjMz/de5uMsyrtfyA/Wp10MjMktgOYCqNo8h
+iACdriEJ5UuOiH6dUkdePT+k/KeDxbYfle1doT/RxPaHn5jrSW4UHhdtvIvxksac9jKP0xcC3gL
ifEtU105pnH41QO5QODhpn8rHfHrmLAq17mR6zN6FaUUXGlhhYagbnRV9nJumj6JX97E7Ex1ptEK
ieTI5LzMipdoFgK31qdae+jE33pB3GlrrEf1uZmid4Or/vIky5/a54Y4Xq+9eyCoSWL6Z/ACYi2/
okffIMpCt3GXud5rkeacEGd8Rj2iHijpe37u/LOKm7eBp2s8v02f4iO7LmHi30AI5KfGHeGWFDsN
XP0suiyjDWwqsDGEgU05+WDJXupU2/ii/nIUrL3qfApNOXtwzE+LPiALd2Cp0CMOw3j4XOu2UZNs
HsQLaNKJ2zRak3c+N13cOHGiwI/e8LDj/qhOASxHefZHAuyAxgG5fWMp0qbvGLPVqsP5mcgXcprM
ZihtyW5xopyZEnmuqotm34lVIqcmzcyQ2nmM5weRt15IGbhJmrXzptvY27lBkWE16pBMTKo56Ccm
wHMV6zbAtuQE2i0LyGu455E/Cf+Gy7QAxlUzH5STn6SBWTni4j/M41PWHeZZrleTO2DKTnTQwKQx
jn4vdVVJag1N4E1LMj7fhVIZ2xK7rKdNh6TWPIMi/IMRtO2KBUp2q0Or16wvd3XStr+7V92R0jgn
eQiCJ1Dx0S9RmWRhkErwEfuC5Evu78jsVrZ3MgJ+nyTrpdjS+uDZ+gGOSC2Y+LgcxsxnN6RzHKU/
uWOuusl5mj7jncR67SVEqWAc74w60HjDlsyf+VOa7r1CS1UQQbSm7PGUmd4edzCaWgWZhPmQSQgI
zJ5tkbZHlKGNZEU20M3uI6O2zb419m5OtQ4N+YKLOvjo3HqS97YM+tQhs8OtSyEOjli5+2Gdb9x+
SlpyZUuZvKH1sD9QMu+EyPoU1HeJp4qurGpGxhFadQL7Htq9tNBbDucIwfRiQ2DaqaQo9FM3guYA
9MF+ZjZLRIZ/CU+i8AA1ZxG2Lr2l6aI50Rcd6Vr3hiWxWS6k3ngreqPJG1xAUkPnKt0VfIYBw4QO
1dnzwQXJ1jUM9aEXKfQdubZWDirtQneXjTcdGH/u1asGyIe0tx61wiu21CNndgmWaiW4alrffFlY
NK/1Jb3WgqjxEU+MqmbnTjxcb8ZEcWMp5Hb+J3iHS7xUhueht7yk7lHZ/Y2hf/KIl0IzR228DRVW
S2eKkua3s57tdBC2zAR79L4GJUuAuQBM7cKMuUjx7RUDiRW8jyFUBXkfZujuTOgLv1w7qXGrG9Cm
+UXOyOUm9d5wrcsigTdS+bocfl9BE1om5J/p8v4t79dkxCRFgNh8BK52LrQoOaKh4ipkJYBWmj+f
ZANg3WrBWIM/9SZci4AcskuORAxlM/tHbLxMz/+6AmZl39Lwg4nvhoo9IxHVenqgkc2nJmTp1Ya8
EQAGk+XaPS8Z97WTS07mzDwUdOgfbhfqEKittTb3IzT6Z6LSGP5Pa2qN5DWd72AOyGF2uGGyEflI
pd3URDndKeYQ22PUXUt1If/O7Kagd5VexdjnIQyR9IIlrXjpNMWrrfVbQHJq2vXHFv5l6qcM6cVm
UNp74wzWWNRHLKRood+rpTFZQ/nxareTr051Xy9f8R+u+DAGo2ccLZ1s6ZD5wlWLMjHXkDqVsaR2
wRgNwpqSRaA1f525PQME+V/rrRN482J/MihFTrHqTBPOYBvxjWB5gbsTsRDP6OuMzKeypLEGet9A
pB9IT5FwXI/c7RqszTWV39PCaNJk21N2AIAK7gw7t9IbDdMt+puLLZXsk1tRq7wD73CRV3CpujR9
bBZJzE/9rmuFag7Wi332XEeZuca1ahWxjyqpYsJZJNUxdNnh117ntA82jpliHQ6x1lqy3IhlmQ5V
lLQinnSdJKj6u4D1UhtHP+wd9C/ESxEImIL+l6GaF2h4wCzbHmCqGBDhPnQX0+e/1Qg339ChpsbF
Ah7jzY9CqR5/yNL0XQlnQ9kTTxE5/1v8bauonH2Da5GSYZhjqmcBh8xeGxsjEVaG5pVDwnIsP1bG
LhUY0K9ILGpBEmrfjzATTA0YMDO7JYhkbD7shFUrVPwxVa42gYoNm84IF56llHTTvOJRa+zhtcmO
Txt2SsY8J9vfH9M1oJgbaZpxdtOqgqPI/fN1Rqjj+RDGYcnZP9LHGVy7t3WSzDc5BJ8YRF3DAVWh
2UJXeehtIU5bsnG0qRm1s57JvA+iREViDGvvd7bnjtINNwrP9UCuoxquzm/2U12EUPjMTRoY5ZVj
ftIdkr4oyFPiltmf/67aY4s29j+3g9jEAiyyOaMxRlHsdm6nctKT1vDkW3gXR82otm82LZU1LxYm
Az/jmYK5v9Kcq+MykqjKapiAj6w33b3cO/CZsVzve9nQ7ofrnnKqJea4jregX9CF66rPKYYpsurs
Q9t/tCpe8Hm1NxgIoIHNe1amemuyy0tJwJ4xKmYI6Z37q3cVjAjlIGCo8XG37OprNPjilK6xZ9p9
M4FLSGQ6CZduxTqAZpgR1Lv3bqSEiSRn0+1BZuQGayGBYqpKUMIU3nmZXPNgxS1EqV2oLND71Otw
RneNqRixVa3/P/JJEM4vQxF7uiV+5Dl0VBPCfudQihBlbjf9PXf7w8d4K1ra2ZnKNWaxJXelhgcV
ikG3DXZtoEQyxbKtR3K2Mmm/5Vx1MNDptcEUxluSKride7O0GKRXiMUvQAAxoAZJRABc+FT50H6E
VyYjYEd0XmWyGcs0W3XfRZhUP72dbOTGI0pez/UVBa216pIE4PY3Snnmq2s+Yp0fyJbCuPHmtAFE
2Zzyx1us2hAhCxzBeif5x35Y/8kVl1s/tMn+htYTc83PstdQM9gHSv94qD+BwmL4Zq4+q7sie8KC
x0rnB+2E42A55JoM/WRtOwIFsWvYZFwFiyb3ZiOvHBhxgpb5dvH7iPJr6M9pnaeEOURrbyqtfXFu
Ho+Kq53YN9Wt1Q4hh3/Ytdx60EL/oBOP/CNd2k6fqZNwIC6VJ87E+b4OJioWGW2W/HMhCyWMo5Cz
fSq21OeN2+yADbd3ZDuMFicLdNyAIgw16ksuhwg7hrNJ0yIIDclRAGt9Ql5yJrqoMusCwrJKFH4h
agX9YrTa535ZPvQJ8+PpZBOZ+fwekXIG7VvD1hSSyGvKng2iRYh/2xP5tsMJ28aygFexltGUpj8x
6cAofiu5QSy2MKCnyeOeocVnS8led/izhIwcDDOVC6Xvktky7JGGjCmJHutaP2mvYdniWvcXGLem
grV3zqj0oLSmmMkGhofIWUUzJ/ugcE6M65lyk7Nb+Zq6vGcRVMFLBehJpO3IuCyMOImL2VCAiVQQ
vhNcNS+B6B3XL/miaZLs+TH6oks6fa1CyIkwZvA/mwYIovSvRivXu/J2AISL3UbfyyspiQ1GtzTI
IMJ+c90i9dhpWHkMHKVfMTvOu4MjEmXYs82EBfWo7zaJGTbxzAPiVh9m/F2YWW6hOc7bHvc30fEC
0ouAaUSjxxvBPXk9DQ/7RQ79DXUMhqaBLl3olzJPX2EqJ5EIfByk+BJDBtIDH41H8V7ou1UaP0nT
CAepP3D61oLP5GqYhsIT8TLxBk44HV7G8lwhSbo4ok1te9syujtYG83gRdYrXFj0nztRb4C6CJ3r
zcTQWIHmnflQ+yGhXExIaOdWw5Yw5wr3bkebrGD8t5Grtvenhvsb3hu7DI+uyIjflOVUjbR+z8NK
pWWu13IFR/rHVvOsM650q3PPLvPJkxJCtHXfSq8fjyOdrEpMyYVthSm6mKjOyTT4CGzWrkESR+Jh
GEvZD0VRs0y0euoPCuprFb8l6+FiFOLZYCwosw70LSmvK1MUVKk/MO3xkoQYwdATEzX/L1HdeGet
wBfGMf05VoQ32bUy82QZ7i7/OYg4cUYP/DSYPRRytb35bmtwyuCKsDWNxWdR/NXBpZNTDxKnsTqd
aya0oc1WoP+hq/PJ3GxdbS4Yxse0rhWUgJnnspvxRaLiHLoGdBl87g2OIkJkpqS14KXfexa6y327
CuAAtxCH4zfpx+0Fp/Iua2SSymcaw9/f0wD/iu4DetSM3Z+eD53YD200/kOj2PXp4Ar9TcPzBxox
n4Fm7PO34LQl9kWCamzaOLmGbf8AeXyV8YtWKEnqmulrwV/09k0+zX6pqaJlSekQpU7BIVFTujh8
enDm+hEPzPhqdQGOMXriP4pmSwajgD3vzg8Z6lk0WmsbqqM53AMrAbLLofJcuTMD4rEjFiju1kWZ
8fKbQwy8M16QjAKv35qHdE+7FVXgRPjcZajl2GVJMOwglpTR0LMdebRGGUlqcrtMVAWRGIzKTsfA
7CFYCEUVp0Y0hF9RS2EYwSi+ioEiic8dFi7RHuU+aRgObij1sJS2Csos33tRnLvHLdkgGIdZrG0L
Usf7WP/WKTHXljk0p7C72WbAPM7Hh+N4bRs/Mhvf8A8xGOj7kQp3GVM/u4sF7bSPCBTQCDRfCrQs
JZHDg9DEef2h0PXxixa2jtUfkOYF6j+hJwXHTVR5T7sd3an/UjjRrwhaf2Jxk+6HFbqn9oe3Scz0
pAITTTFkU6pTclZ+9TwEu0D9Tw8Fe8RQCGOu9x+53qmPiK870nvbwsKdsHOMRHDa9CPoJecy6tSb
zuqM2Uc1SG8X5p/BLX/NsqhEPaxOEg4cn7KSDj3ajPDPYu/wrJ4MlEYtGgJgvPy5bagBuCTTgu56
SNaM136tUriBbuLXb525NYepOixAhFbv6E9BRi27FEz63Hz9B5paUee7/aN757f5kXZNJJO9/6Oq
CxCvd6EltwxE5vMH9wLaSIAWGLoxj0M42ayzamuGTvelgOUv245hanziKMTunxNz4LhJpXGxEnii
DkAuo3Uk65Le/wX0hFX/DkIOgnHK1QobBOBJtY2GM5yXonakelUUjp1q+wOyljvssOXPGNX1SbkM
5YvYlpA0ep6mvLe9yzsaH7tindS7M5OxECSL4cLl+h3XN1vIQcQkVuGU92YXM4SmIKH5I5Lvc80Y
DsMV5kElGGp3ZXz1H1iaJvdKWWKhBbbCegzwQZ2WXkFNuWl4YVPDXB0HCvK5TvSIeoprrjjX5NOP
hnRVgtFnpRax/c7HFMHLRQVSho0mRevrAwHw5F/ELUaVUa9Qg9a70oTZNRYS+FAnOBjYHaEGGa+/
iyiimwdmrGTyCy1hGdYQy3LNMztqv0SMoVO6OJz1LKyDt+z5ADpgUtf2kSOnaZQXgnwKVxMXOMSW
zVsQj82YBldub6GULoJ+HA1TWXNxstPyskh5iUjiOL4u8GO6G25P0mBLQNoLvgZlnI9MIC6cqG8j
8xjIPEZBwB9KIk9aiJOjiZbU+lApHYkudch9jQtp0p7wJ0K5N9f4l+wbdpM+axGSZ03bnrvLJJn1
VX8ekNSFq+oMx1wTyqlghvPtPvqL3g6bhvCkBtspTl3FMQDSFIqZ1eUCvd4L7CRcE7buoL/JQCMn
zOC+0K2YQ7H/Mnrib/7MjBscbE+tGlL1JUMmXyChyvkN9NHDsY7MyHoyqgYPWgKhwWuA8O7ie0HP
wByujumHnVvPwC2JY9DbbrKQOdvZzilBYeBIb82l+zKt3lWUQW4YcXL7x6kGvv5CMalLcCrARm94
7NHwfYketNVjfqWNpOtAtPvlPSH/SK7BihZPu8sOClKThsYkySSU4tWQzdjwKht98a9tlnXzfedN
ooD5I7B4+pG1VzpUs61H/Mi+AJRSW9JmX13Br/taXI4gS9ZjXmWgpY1hYTIX+CJM5oRfkJq/ZUxc
JROFIYiEpyiPKkr8ZCBiBGZlcn3YjlRXOqC9n6VCiAzt9XnzG2iWqXKQx8FA/WPNerFUIJVk0o6E
YpNR0JwOtoG9SRwKeaaviuXSYTBKXCNoluYhE0zkWdrFzeAM4Pai8emr1uuX5yPJInI9WaL8n0wp
WZuTQfAUxO4ya9LMILdmy9XIGjrrrHckd+E+7KV9Ob91KpTzTPY+UK8TojELO2K/MrBCFWNXHbs9
MxSPcX/L1rH10Z9vfV0vWrDqpH9Wha+ywFEVUM9Vr3lzn5N9hgOmIoJVSNRQEu/UVHTdgUaQMrnA
GGxlr3+hZ2lXggRj7pVuOL/NTXBy9KQbvAS0xHinaUG/JMaIxYWVYO4cTb7AzCsbGcEkGKmJ5Nf4
JrkchqrgdDpOnWmKlYhJw927tBBD4przHWwZjzgP1XrcJL3yxacxW/K1ngAfYx+dJi3iuu56vB71
PVN5X9X9o+bTMcDVMUcWBHVGu1q7QMbGrvrqfI3P4wGBst09bUP3xrhU5GIWaFu35hHLTksUt63c
whZG9nqw4cx3pkeN0F0RcdCWDsc3KZmQs2IXbV26xwNkxu9cSFBi+MrKO7kcWpJ5Gh1dkxYZP4GG
i+vMfX/cmAWcZyNonzjGJLKaEW5qvwnaGLKbpOt9G4MDok3cPuDjjxIXTHl6mtYCQ8cbuBZuoKmz
saS2Oxd6Zc1F58PjzoILa5GwNjC097ojdA2MI7kiSt9E8MeQKidiFaIYkEdeZj4ZI9BBkbKjrPrF
Z13s3TUuB7bWf+XwSA8D/P0fhglmVCwX9dPj60tiDq2RVP4hGzvU4nv3Qzh+yvfKRE+W2LRW4YBZ
KthJXwZg+1UHj/308xlLzNveY+AUFW7BY/vQsWQoqYNNCDFEk67AfxbzkSpSEn3k2YWIAODevRRX
B+eiJwbu8xcE9V/zKBpplYWw9bRpYS2T7DR5GPAGHqZWi69DPcdxdU3Be3W/uNwB9MlQiDuzObIB
1tADuV2HA3lqEapoVkHIG6BNPiQx+p+Q3s7U8Qzk4yvmaiNSKqIRbBIZE43NPVdD70ptXhFdon6a
ycFHt1z5VkdaHtO/IdE3/bJYg6Zb7uBU2EjbGDWzS2BDcGG/0YCM9dLYkdyhGOOMUhxBwBeMdrTu
A7kJdu0lNElxSA2gjGzJvMy5cv8r7o5kXWc0G9KMOJHaB5hcNjogP4FEYamsGF0vz54eUUKvaGvp
dBLidLvEimb7+PToRcJ98NFdhlyFhjyfUjdRc1eGyxSFGcOsvJKJ9yf0Bm9k1RVQfAKZl3xEAE8B
QVsiG4a1XHVh534hUaJBxXdM0UYVrTvKqGmkRSyy5lXwtOHPvRenU5f24TLViqwVZ5HprHaNOJI+
xVOQTUACFZdnAKOJTTyiNfCwWN8ZUlSzPOqHLrkQLzoofwqDLv/pG5T81/w9m/Sqbp+7P/Zv1Cju
qX0BCDJXbCGVRCMBVU7fPdgATmVhxSRI9LU0aYgvC8Qo2LGSmepJ12DyZbpA4HOVol7gHKl7irpr
t8h+6jT06vH6FyWxFc0tqpf+wqfButMM8KjOr6xyWwTcndyiQS6EWZUYtOW66TAZwe0j+PI+iuyp
YU5Vda+a4SsYpWlx1Ta57Xeb7Ga5d/WCaCVuVqw6g0f2SYmQ1wYLbR3cop/J1Zln3As1FSnvu1Fz
m8Cnis+S7c2JHMCcNMzVR8Q9q0bvaNNldyf6E9+iTMHZ+MXR5vi7VwUaPz+LCOCAtvnGJcjwrg67
4tJJXu+T+y3kMj3TCZzHkTYBQkESBXFxW0OyOsPSJdhUPkHUeRZIexdoQpBbsb6PpqZCgrhjHY12
Jd0Hh+RtnP+EWk1VeeEqSpA2/CdgdDjKsPztRJW4p+uKyfUlAIwWCqdU8oXEQENBxOz9X+TF8Cj2
tRBb2cFwctGWlxt4rUGr32SNyRzs0mX9dNgEIhdlQPHWCZdjW0JwrkjJrXPcy43SYcVxRHJweO4E
iaH5yHPyGkta6huPkY+f2/vqCm8+AdByg9h9iU9wHJtZLqFRTkKmT/nQycI28J9w2dIct2q6qO/f
y8g2s5mOLQyZIqwenLbIN0tNn76AZj9Uvrx9NLUNKNcV7ogfqBjLvbn2Ijb8zFHm6MmzAwBX7ymg
zR/y6TahewAwWlHsoHxYZV4ViQXSWlsYFwvw7VvpwSR6pdO0xPbffjc0KjeZTT7SLWRM63BElk8R
195rRvAAvrWZ5AI4Dm8cuWDUBuEKoRpkSpa59vYuGGRp2pnJHmtx5PErK+nnkzJYudes4ihDLAr6
rjrun5/Srx/4nWQavalXxlzQgOFN7XClAHCTDml7pAcpUzAOEjLEPj7pz4x8PMW1wSPStAnL+RL5
JaxQVafkejf0C3DIGuU7DpfhemlTS1FeEAQswMc7j9TnI959WHAhSfF8l5YobpuQGZmMj3a+UcTh
Qb3DhyAVo4bPD/BDmUdOiH1qFjgqbKQjXeZr0ynHSZWpGMlheIYilNIxmCt5fkrc7weEAuGHU5S3
iY+dRLFcjhK5PUMxYshLwvPWAhCQWMoBBmrhGklgxnrsu8yN6cMtvE3iXtSCqhXDrPG5En3N/aeI
r1Lt6UZ0B2+w2Qm4nietCLRukxBoLEweq2Zhfgpi8iCyF3+S2g3J9ajk12wJXjdmVvy4m+6WvDc9
nvGAoeFYyCHKv4zUTxwiWGCtp+q2ya8/oZZ4Qnq/TkiPVm9m1KAFwcCjFwrPU/QETtq4p9G3TumI
8sYkAt/Y1hoSSfuHApsEHo/8v0aQcCsrJZutYvyxG/oUO7Yqg2s7oh9nC4MeEEWpL0aKnV46FZrR
MyZAv737f73nk/tYpFx+51PyuVcKevxlaKrH1uD29MAPfM7i2cNDOqfiowuKlhlFtJfPoh94BGRN
D7VnXWqzfKzYYby8UDjfMjl+9orEj8QjJpN0MQF+gyPJfNP9IIDhwooaU7HoNe8y/p4VsnpJOb90
USQfheBfZW0p36WSDXun42UxW+VbvRLNkmk4fzemE+pLuhxUp6gZqe0uTSGSSZsLJv6prLK3PPFv
yvcejVfT9SfqGbXfsRn3YnEGu6HgMImOfwV1Iloc5NQabssIj1yHT5LgiXuAOdK8ZCQ7XfeniB6Y
mFV3E5uFeKyvn2r9iAvb1iuneP3G+OfaF+7c/IL8YTEFMkxQ+Lo4xLQsZBExxyjbVJQLNabSAk+k
khQQEm9xeQxDfhRbBpZU8VV1iYxrhYuRZTunqJ5PQrB9JY/KkXmC62f8YqC56zEDLqfTUOEBeOnn
QrlA5cvO9RrlbO0VRSs+uTsIww2bnCOpZnE4w3DPTcz6cdG/uI64fablW2FW02Kd7zYjQh2cX0E+
IL29EV7etbm5NAR/OHQlhFdjk7yZ51sk2MBcogY8INJP1z40NDUbE27woQZrmsWK9MuT9/UCo8YQ
Jr0mblHcF4SsZRBtmLiaQNSCBBLcqBKOoq+EgVGl2slMcfFNHv/I7l4EeLN2N8Q2MgnsXuSUmyEV
3KLsUktqykyKa5kTS0VnM8f3sWl2nDlN54qAYfdUbdBHWUgwkhnwbJiJu6rqwFiIoqxB23nMZVCQ
SMtseOws1gPizysrspCWem28Uinm8g95SVXMheV1ErBJmmpoZwzc0pROcsb52OFLAX/pYx2BxDDk
Uk0fEySwQtscuS4LaTQ2cFcuytknuc25NrXTYMFX/Bms9vwoeMNlIEpKe4Kz9tRUAUipPOW4O4Jw
o1vS2572CaAdPrXhXfquPWEmv4789ByUNwCTAPDUckOiKj9NnpSB5KKvbet9gDzLyk3skRRIz5P0
o4F56yCC2o2obtAI4OllV2pTOVU2pHkTFrImKSPDmFD9iexPiAh/vs7WYlALxSAcFfe9BTdknMOB
TOu3w9uHN7HaU7gapa5SbCSM1bjOZhkSt86+UlqX82W55+BTN4oqrJPPSZJXWzhmrT9KT4l3fc1Y
ek3yyxiFIK9ttnlChFTEXHEjtMIIbo+WdQk4iI95XP2feWFlXvge7OkZJaTg77H/FkNtIMyv1ChS
bEntRiBXMB5GzkiCHI9c5D86wtifn5hMBTrzo/A1xAds6nOXeAcmEH8JJ4FSiruCFgP4yPQEZkZ0
40Qtr/SxVyS14qYuab74mhUy5RFZyBerjnZPzQl64P0y7GRB10Bjn938fchgS6wkV762oWA7OHHH
7uxQb/+TARTWNwJNEOaXaDhuYqXe5HIBAoxHx8x3M8ZeNBN/d6Tbbb8v50/Idz/DvkcgrVJSxaQy
PlFO5ZIrHuxdrDoHj2Y8D3r51NkoGG07exNgerHYig0h+kpbKRd7/R/19Axb95evFCPYesiuRv8V
nQ0NTRgLiVRtBz+h9IWF9BxGNRj3EsVCKcuWHnamwbaw0QJV/dDeY7sTKAED8HMuxgotjP3rOfXk
I6u/bbuWqxDJ5vrAqGxxHY7kF3L56oHEdBU15Om8cM4Wg8He1TtgRhEctWtzl1GvWQP6tIYOJZ6x
wzZl34POYAm7PmJjKj3hyIzTQaUtGNshAeqJm7FvtGSGJoUEMyR+jl38vrpcFpJdEP4lk8xx3PMU
uqnaDoFxUEudd0QUlE16TrNcNBVj80WY1Zd1LuRDyWF1WGZ/PKze7tewIBp6uIrEuD+qTIOY5F0E
kvzz6x09eeQxfKQdCjFJtIEod7A2YhDHkb3tgxk0lXGDC2GEW/G0FjAzeUPUuUCE93A8EtNhj2OJ
sRqrwm9kqyM0ZYYBU7E/THtvqHK7emDOkWZqLAcmaqYOhBYfXuyLBxh5h2eIq/83xCEsZaiP5qtR
nCQNzh5MEFBydmNcZvivRJDRqhKMWuurvLuPcAj41P4cg+2Fz6+KjkXrpGkke448MkPo1dABL8uK
SJ8JxYlajOF0bvC3dV/rn/YfH2pat3b9e8pVqUI60yJkOinc0c1ehUU8jv5yOj4ilCVFG8+VWKKm
pcWNNwAlSojJyQ+g7Bsr1dlXwMkPclcOhpa+gEHijt9xDtImulyWRBZCUOmFEjnxOYWQvoWD8uYU
9HKln4JY79v0tHvsufVKke7Or0rQ72ujriGhHzBPaG6kb7LlXXYkxNkFiv6HWcwsxWf4L23zSMOM
L2u2UWBg2UVFsIT8+YyW94vFdo67jnHHY5QJ5HVDWoauXhlmaTqO9cE20yifznVVfQ4cNuBAWY4J
oLrlELO/26RjphTCFKYbvRa9GP/GLigeyG8myMEiq/BKyojjgbEm6DcPyaUmLN/Bx0/4xU8TC2gR
fgbsDAldcUQpO4A0vVx7Ed2J/aG5HCmw+ngzyWAx+GjwFhzGjRc4/W6w2zvBRNAMrLaYzJ7T8h/J
DbFTI5VoBmT5GIEjPEHZm1CmAerx/lHtI+n0Xsz9/6qHtVZhkQMoQnw6a8RiscDLeTGf8oLnky1s
ovs+nxFyiMf2KNlNkpjU9RRaYdRjQiybBipCPiD4kJwxqk2Uvuzkqqwch2nqZy+LnjfdVSvBxSma
IHmcts0xngXGDqDx2HvqeZQBDq3HxuZ7d+kYE/U1RW1p5x4s7yDOUYGqeVUFYP3/lnyPNsD+TdOk
0ag6BiDnz/0CngzY2AtGaY9+XJq8NKo/yxeD4h9U/iO2g9mP758TIJFMZ4DO7jYExtjFrlAiuMyn
sjYt1rgI2KId9yf6sx7OxpaVQbeyl4anqL3PGttmf4PjFKvCxG8oqOqC6yIdAoDUWsCbhGaBUbEC
OjG69kSP/itbQn+vS68sHlC+0cIwTDYdYj/UdMC5cjr7/ssMRUJKv8ChYvT4Kco4YJYMW97CofGT
y8Olua2aip0B2PcYln4mcKcxjOXH10A1jyfGfbC67tEHJEE8Hs7KZV7mifylNBBdG6d4cVLW5M9x
juzKPFbFX8nXIgdWFAwDM9DfiH9viG5ndK83zRnGbkmc6VJz6RUg45VwGKDNuQGZHmWBjTCxWQp4
CE211aEdvimjTTaLjc1yRD1zL70dzYYaNFnu9Pg44ahDyvsV4Am6UEJaLWRTwIzlYhg1pgu8+dTO
R1gdWKQTLs/t6cE+cztmzIr8cW1uhtdEMobIz3Flf8AqNL+EvwsGuupJc+voafcFMdhrx+RrAvgq
3oJN/VbaGiXjDYxw2V1A2haoOK1qDvVOPjaD+5in224Ax/NZdzrgCpNFwpA6puFlwGz1+v3Bikn7
nc9+owdplNP+IBGo+bE8ZrSfTV67tApQOPS3zDVHziwzoTgaq5OeGju/c8QPTCmBq53d6ka+Gk+B
J/895fJcANYQmrkAx1W7dfqwlrFnzkCsXKJIEA15ISuaLTcuF+/jeqFaTnzp1difsRUQe3o5csr1
GeTWRVIcblbw6NrRt3RUQbu7DjkWEaXO9pHPSDoWlsZ5slNt6hiDhsn0RQSpMJSr5fGScV1ax2Sn
yOxkP/jyOASra5iiV18dKkI66TmsehMVCB3ynMT6fXtt9f1usD0gXsRkuB+jxAe7iJBuBUz5LDJL
A2GuVjFbH4HIZFpbE2xWLIKdudBb2oUtQuppOgUTUZiflt5WZuyOuk3sj8/aDbnBB/mc8sHqaIwc
ujqaxZYj881WG8FWqpZJ6yJbJ/mONhT+fED/NQ4insY6vz4dE0M3QJ9nWf2JeEY9VP1ykBjqZvbx
9/SfQ0boorEdxQBcjiES3GNoj9MyWg0+cG1gfqWdxU6ViobVd/WUHbPUtGg6sUkkqG+PSBkZPLko
jmJIn8ajb1iGAu8aIpGMyF1E7v4pBLlBzpgDWEJx4zKL7TUvpJwQJnNPV/0uK9XoZygwdQrVqEBv
5OuK3xfzfWwRo4YdW/e9y1Eml3NASOe9nU9Ny9X9fx7MW98TwZ68wVnT3VYHADpeTfPiUK8pZc0J
8b8eE/Hh1RsSY9HAAYW5pDow9T2T4OXgqOQRz4Rk5w0Xgrp4lruxLhy/IiicZ2mtjWBVrAaNRMhQ
3jvGowf8Y21VO9ZH7WorgmvqYNlKSypFmCfrAl54z7H4pgN9Civeid2g0GPYADa2uNleoMihd29L
HsFYehiLvGyllxXAtdBIDsQzh6xMsIF/GuBEXMCyD7XSQcbs5jYdDNdWQja/9f9EP0CSGnTjVN8l
uw3s8TzELXvz1SL49NneVXJIX3f7EiF2TmnojedHPr9qcqYAYfwtDrq36KtzqZSRocv1qbAeQXTw
lz5chWoTP0Aul+b5FX7meZInrx+CrrbeM7LgbSY20UTl6CdkSJOvFsNU5TJ3t5cv+KR/HdbmYY1j
vEwIoHQB3+Gh5WPMbDmhvMQ4mXX49ofA8pwtCsXlWNvJwgdtpmlcmbfMms+Xw2I5JDFm4r8psmU5
5+WYhUJ1Xyqt/etlXxTyitFUQe6f8S33EV8y3xSuDJPDtuRZq2yu/nA7G7UelpNQAxCp0Ul5lpvd
Ds5w4A+roQGw+9ktSh4lKHtlCqbkNWEV9OLZmmsh7GU07ESg8Ic6/ISszwvTq1Eie/e1I/HXErxS
sUHHUZSFynmKUvX0mUa/hygV8hOzWY0J7vJ9B5DG0kNfz/3VGaw8aGbMQ5P/zgqvHiNBHTJ7fcxd
Xy//1Vo5v2mxXKYLNcjbydiw56ERZK2OWVTE/Y/gcCfS9tbajOmAYJBDbZQH/MS3weGk59GkwzdQ
QP6eEsDEa4VwZsCvGK/U/IGiIQhQsM1MDi8WVFb2vP8uxtSLpn97BoDshZLk3Uxnz/mMGbv5MOCv
C6R7TC1oHLMoCSjJaFOvOZR8TNaufuuiPSQbg+G5+hreGsljlaeHq34iCVTPUBB+gEpV9vUR4HA7
rbfGINTTPn4Z7RzAPeD+1Ry6SIYmlehvHXOtmiplt5BTPnHYSJ5+RYZX/J/pEsG32XCjFpv3ECA5
Pdlo3NUxpdbdjQg+M95mxT9A7EfIZy6umfm/zQexrJ1kUTMp5oo1bnkFEQDlLr/sd9D2LJrURTNB
wd3xTHQ6Wu6x1dBSUObBVxxri+tLVSsspoU4BTmoJB+6YsGSudqZ5re2qd9bEmtKdDfX7MQozU/5
M1ad59A9/6soisRPDFTL/252ZKS402Lj/uReFLu+UIE/S6cEFkRXkRWeYyN/QwXuqNY5BfqYoJ1A
BavGRp6J0wcixJobNPj2wqlCR7qLCP0dJYLuUI5Tg2J+6RSDOw8UVRLn/s19mR2hbp+To7QfUZQO
GKDYZwgRq5LeTBQkZWo+EAqvezKIvsj6m0EXYgWj0PaA7uiMZ4Ivl4Y6JTsuqYClm68/evnyIKmZ
oBZYquCpdFb6qZGwiua1cu39/RH0w6pTojh+QIpp/YSRCi7a0ZrlxJxadc4wLl4PKLm40Rhe28A7
f9ieQ1YMc7V23MXc5kNra3Lhcl3xH6O+1jxqUCA9VtyAJtdc1gn2rlflWklzgp2fkRsfNqI7fgpX
RHsjAQSdcjLR3VxnrjizMZPRSjF+AFppK+7RRuGXV5lNUp4bosi6TSKyFKiMRfd4HrAnqpONjARN
/Gn/dYDZQD6VImKKRXXBPZx5R7h2G7C/+dleDtbasyEadGg6s6gzoNDbX9mUzeUPO3HA3jum+af0
zUrheZPW4tdPioQnGN+22yTMEe+TG5QVcBlibGo98a3dWxl06rdnZWGqp+2vj6X/RKKolT2L94rn
7tgELjuXx9fb7gSDiEogp0ZejfuiRDRi887KBU0URNSG7nPWFc1AlzwdjXldRtqyoajADhpx0hiE
TRRNRR9fGE3lMKuT1K9n3LODQ9F4/hEKhAAoj8ml2x7ZzujZaiD3Z0MbxPj/fsBCAn2rkuOKmjjF
V5d3j/IpgBLpchRVNIpDpSHT8r3Kat8EnklZ4qOYJDHsx7ttUPHIdHAIJi7QoKfUQYHocVje1HFN
C12CiakAgevnmEPa+UM7QG5Brp32Cn7P6kXgzEG67Z9O0YFCD76peGGSeG1Z4WRlDcFcCw8mGbhm
9uS5KtiZArVVcwGIe1d7N1F9A35EefRc9KiOhgD3eEdY/lMAFLjz3xeCCMtipdchlDp5FFuzWwkS
JKGMYj+zEE3a169cUw2iNJwzRMo+g4IW9666xhUqAXAW868PdJM2PkpRsbcs4VU60ZcnvFS/5SiP
KeN5ZStKsIj9o0TTiSsbduYsIv2iVOq2xcjzZqf9bv/CupIZxB7lLCnHIzT9DQpPg/vz2hlyKVJ/
41ZxK1QNXbaKs54T0PK+5xs1EKP+ToJsKA5ETc4nHLI17iYNB/ksTd1GxHN/aDUfEa9Ll82pYgaM
qi7D8ohhttJq517WcRSAk3izIbEOKgZ7dQDlV0RWDqtfa4eh+VXt7j2FyhoFHQTbE/LwWUd4ka1+
NbqTV0PHn4yEdfCsssw+AHdhW3hQVMaIK2Q3iBIOiu8Q8C2ea/54qA4CldNO16izjSGtljg0DPrh
IG67vNruCdtEhRBpRjF5rNDhfWj0SMgHO1UOt2QBDTxatukw5lq9+yTQfen/oaut3CIt8+H6v4eu
aagKZSt4fljh0Bp1W8Qx4FVSB/7BndufRYUZQ7mtR+ajSu/2dt/x+xAsyQm26vTHXeO9YAsqemt+
y6jrwplx6tFPwobhvK7qFZmQN1FtVq5ZS/eej9fCbBOLsBOlV8ueK6GuZuLczftzMPFiXfsqk0CF
pFltj3Ml9US7x6VovKsRw/8LGIMZUV5ld/GEg3kBk1/ej0Q2TH+i3dja2yXFQaOQ0YqOpVdZ2sz1
vIDcNFvDfiOPm1PlrrrybZunximU++J/f4iGL+liO137qbRZpaNN3kweQGtdeaVzfnVf43xAaOcB
GrKZkHToJ6mOdYyQjD2P1jqWkcaA5hncZU3X/lZKvpJTSXCmsmLLoscXXTS+c43nTie1cVF8ER7H
3SAXS2WWSA3GhK1ZNc6vuMr36BrjDsvtGnAmaz/M859EKGizyjEYb4TE8TpusVsDeiiRwV8ddVE1
zPg1h686G8aHgaCPEbE5gVDOpRTZQsqZnTUBZUcXAv8XMD2WMt8FYZb+q8HLH0cT2mK9EBkM7x91
ajucOCtJvLck7dKkFLRs8EBcm6gsnF9ZoA4geeuLHzoPjoihivCe8qi2POWZC3hoFy/xqUZvSrhf
2tJVZavMK6nOOBUFEjJBpv3d1KiKOEnxWywtsr+WRIHkM3X4fEsmIQTwjQzK0KE7YyP9teFbNc8L
T+Q0qP/te+N9F9cwo9yyVk9+Yo4ErBqIgg0wvQtjkVW2HWweA2/aO3tQsSo1piCcG+TASKYlfAgv
JbzafOBJeXL/FVnnOe4ke9mU5h+kfn6KoEa3IojOyE3QFvLeIk1sEFn1bqoCcg/vNuExapICUrNV
ced9uzxJgm3dFi2EQsVYinmifEBaFs7KOSHpCzYTZEM9aH58QyycteX/qjQABhK5LUCOoL4f3Yle
pEy9qcoNeR9SP03d0zVePSVbMVuCuFzMyV3/tYNdQGvK0km1kQgceRT2f/EbyJbRkNI3D1MlPs7f
cemCGqxr1gCpjUFdI72DfjuxAeLwcTHTQkszBgx87l2gkjLUrXxb8sW2GFEp1oHQ3eufooeCTRCs
W4mDfV2NcPDK+reMIE9Q43KsWVv+WK4oNt2oLaT36Z5BCZ9TlPCvoeJSIgIbnIsCTqnlG0J8yVjd
BlTaWmBA6ABR9ql2TnUOoc3YKMkZ80rG0+p6ZkGJWRgWjoUZXurTUXWO4/eTLTL3x6eAy2/dVqjo
nyTsso0r/2DQCnUK9WqZQIbrul09S7UzyVZdm/mErJAtG/2i9/PHymZbXqeJqxIlMfoSLFmhP2MC
pK3O69B4fTiA03+4GJeSU1N+/v73DcGTOn/fJPy21PQWKL/drQeNBN0QPZ2U+QdUjAaOm8jaG+XC
vGkvKt7mAfsxzq2t3AC2pXp7u+btXTEN7f4g3mAqGURdyRXcZqNCKoh2GWlkzlrcAMSm2bOmtQ5a
HKbWIzS5NDqO5VETprobui8sG3yDpoPdkBSW4vVkKWbsI4krXoLS6uPEQlwyrxzOmuL7Q71+J9xu
0TAUUcVVCQMbC2Ym6em+8Xyd2HdKpSx7Pv0l6mKC1xK8LxF+XMG9/2jmwObKOX08g+USJcaQVkaa
3Rl+ngqa7doM1r6XG5hsREYa0CVmEcvSK3soO1XCE+no7cm0UXzvkHvv0mrAm5fJDhz85Dh8z0IH
fqDIyFytLqHkVgowM+UjSN9oWouAn9rERZvYxob5f4LpF/35nG1p8aTgDy02GDKOCmB0YNH4LKEy
7W239tA4Nde99/GeB5/OvEsTZaI0Jh6jD4fUCtfU+YfIazmmLh5pYYVq/A/FpKkPBN1NWmFnjtl5
IT1Wcqhz2dZQe6fhDl2NItAfMNN/hYH3q4+6aEkiQPtwbARIirsf6Nj20L2PvdtWY0qHX85+9bc8
g5JYKsHjp56ZPcSxV+cKMm3fsZ0TUV47xS+En/sGgnBQOcszn2EY9sSHoT4VCXp4MK2BhuSIFL0U
+Va/tWHr1FIKoAg6US7y6KCXfgptCRyEyMw01gXfZkWeNrXAH9DetORtorPtXjci/A3/I6zoi1H1
fzLMvF1SZI7gLSONKNauuA2vv0+ZoP3vpgvMF23gT31HuFsY3BnLOj7LUoIgjvCBDzY7C07MRQvs
jRJE1rBJRXpOTVWZNt9rfZFgGS1W8abteU7cO4n9/7yQBzw+8OfMU+px+JWJ6BpxNqbDO94b23Hw
dtTNb7eR+3pTUINidpgdzjMw0Q0Jk3Bn/Ajb2h1d1Gk7ArG8ODHh22ck1S7OrczbaYEumkiLmknH
MjRnWPmW/QB5RA1D8QiuK/72CzpIOq5ORZ1cUyMd8z34KbBsBezVIUBBtbOFIGI5h5DkAIkXzB1P
dKgizzCHvM9LAq67GcJR87a5sO29yh0lH5vchnEn+oZa1UPNvnykrxZNuZbypcECXqh4drXe8DYS
awqrBAko69LOg1/D0cA1FRc71KTnWc101hbnXg87qxMe7XFt1Rp0UtTgGJw8HLhTWsgYh0AR7yQm
C2GDY3rjCtY/GVxmxf9zKwT+h9atkgIUXI0SmuOZ1zh8DOU9Zt5rdXPXxsfYCvcz+t63nqOr8vwr
ar6oCMVmIHvyKq0gba/rWKdNLl4kgvejSHHm69h2Hj4qR8Dz1s2hAZ2qznTo9bo3IfEUhvPcuSbN
bAtctkrlNWSseuD5PV2GAwpg8wEzJa5iQkuLY3KTnkYbeRLKxEsRVjLHgo/Zb763VpWss2p//u9X
6WJ0Vg36tM+TdWV3Pq7xu8+cdTUxLo77dI5WaefvPwcegZwv48AgwYADlRwYX0Y6aYofVpyPYD+m
ZKg+KcZ2CqUZ5ZiAl4s0HC4LvbN+eSffDh23QpRHIGy6nXHFrtZcNh129G3TE5WthnaV39zL4IJF
IiqH9eyna+Sp23vLJOnmpgxKxSxf5RmhzhTHRaO0d/Xwe6HRjRjIihWv9XXBja+qlitZ6YwOxBD0
NPUeBRwVh4QW/mPSycdldyR6o2mpj4X2pOVm4oMuEsBkxZTfH88AsLPso8I5ZhZbaKqzWRY54Bk6
WKjmRJNQThSO8grMLJkvURnu2bveA9HOa/7ANReCFqrRMlrirvU5ZJwDNwm1C7JIxZfEMLmBMeFJ
mp8LwosRGKsZuh48t2d7kSNoYTzQ7y6ctHmxdV9wX6ZYY9YtCWEDmMgJam4ky6jVyTk/ArOs/s1e
ioSre1z41hw/sHmyHA+y3sqD/3l+tsn/R4m6HbJ60xJmxm8/7yEr7+NIFLDK6INXeqn+B0AbkUdv
qDOlZ4vMki7+Oock5vIXFDu+0r2QeCiqHeU4LXuUO4cBDYbYu+716liIaTPqLOd5IDHnzSvWzKG7
lbvzslqUlHE66e5PsvNNDfgLfu68J72ENI5VqMydOrfQM2r9vQ+EqC/LKDNiMbybWEpULhOS5CrN
Bzxzbn29PhAUcp12AeCFqziPsaNTcZdzhX6cjS3VpmChRo54TE4kg3mF+cP42wrgnXDCKZ9cUXAG
xR47qKuT2j52oP4hu1E5tSii1ugztDZ0xFBrlQk7jOOlBMjmqccBzPUSGYbLM+TZuW2PZjpKE5j6
4A9aWrcbz6PmxIyebNXA+cAfdF3NF81xFGNh6u+9RFDDnMXssUPs/Ivwf2ibSczfdRck8tT2cam2
Eba3eI1NH9v0D+OPyCd4N22BE90Qpk3sDNMK1yiLPRV6NTq27mjpavHXpneIDFLw58VZ7LY0qCqD
+nSshBNWzNBjdQSS9Tt3LgdDRHyDQYuS8W8li0rkdz1bXZ1T0ycrqatXnYfehsSdBVePlinFrw/X
2siQ4935oY7tbnfW2NO0Lua0eKAWG8RSvgCin2yCZk1EjCkUstpek/lJjv89oCRIm84gCdnAaH0z
eP4fQ2Bxmhtu3j4BSFwmk/Lprs4JDKcTqRc+Obi5IsbW5GSjbIOsnx27k0a0S40i0Qq+4G7ARhUd
W+qwCsH8+opsvRmsWruj7zh/Z57v2x3GHpHUsbbec81RzGH6NPQ8DGv4vGBAdoFg8EOQGZnmKK+j
CSd+CAMaNV12ODBoeOIvzu8pbsWPiZCYdPngUV/GK0t3D2M9uXFuWsnS3I8kwR3lHUBFGRxkQphX
4TCFzbvshPXd3gy/bLQkot1gdsA8sI2IERDPAttWjKIii3jq1w2qSVVTJmGYMg46UAbhgwKmPffv
7kKvdtpJ39f+XnhbxdUKnP0BIwuVNh0q7TPMKFlGXq1dH4uDrB2W9zzS8EhnMX/KMUelogEEYulz
weZKzMPw0gAToIbwGBeI9cBXljOuejVRjURzT46/L8dJlauf1U6t7VpLwENbtZiWu57tCz61DM90
L3iZOBimbZfmRpGuIhepg8yiBqPmegLz1+2wfzFj56pKQPnUPHi59Scmr+h5Bo8Zspx2UIiYRijL
y8hzrJJ196fsTuPkRFPhHEh7qaX5Qt/aFqyMrR6/K4lzoISWLwUDx1SaT+dOHVKe3GWP4DaUiAR0
72CiU7mnODeGOm3ECC4GMcGONshaAwFwoSgql9C1z/wclcRm+wVRCzIXwZytI9Ng9dWnGrfyzm22
gTdMQKyMd8ryhAOtkXbY2WPo0/yrMbCFDaVKNsWe2k8xMlsDEGnBEjrzTIPq7Xv2yfESqsZrCK3m
WUtgBmdjic38tbZ3hAwHdzMCDPOEwwNQp9iGAD6Zer7JHd7k4fpRLDBLfkARdSmFxjdzl0WS+aC2
Q9Xc5naTnbEuHesjnGVhP/cSEuPggF/aZ+YiRK6a62Jk0slWKRY5TlQ7taYWy//8yU/1EVNQ0U4f
m+b+yvfujMxWaQLvJGfhRZduei6MSGvM2aqtFUawyIejFXzmh/W0L3Vt8s3IST3shW6bEnAdOsvp
xHyOuK07vBo1j3rCBP1IziWoJryUJ+MQYP+3u/wbdh1sMjPOvJJej9mpE2RxZ8RsSqfId2/tC7hj
qOtB46Z4ENxCObZI+w6tgDKM+SDNLPpI+LK/kGi6DVf/E4eg9djLQcYNa5j0i2N06AZLtyr+nw3Q
dG9Y6BJ1Wc+vIEjdelkEn3V5nNIg/5zZIlteUA+QBGTGhd78Qc/SUNGqni61P8cWu9oDiw9zwoIB
Tn24zi75rw9VQaEcqnOvBtzVONGhr3+1tdjUJeDWVGflwURRPdm0sjqOXKq1v2rl67czsa7pGCNC
YseP8zjVN0djy5ca2BbnSuVsCCpAmmQlnybMUYNf4oflG1IbuojNYyVTW4gkcSNpcCgbBiMtjBo3
z+SlA8ESNo2TxiYs+yisVtBdGX3ocexrN6CIts//xM8wDXN9HPKS/9LdF9eE5H6BheTfaqTleyjb
VbObjKuJ3rmgeamg9G9N1Firp+WORFBHXKvD+BE2ExId4ijaW9qpXJIbjJwzanvzdFm25vdm63yq
PSzWPJqrPvTaEhFaOGs8zPCgXSiQe5OtcrqPdd09RLnrknnwgzgl3hGAFzT69yJQFu/qYg/lP0st
kfa05AH10sMK4ynXBY4XnWfcY81GB/7IKMinnjhRrQaIYRh9pHjUJmt8RDdglmGHvQGMoYQ3z+MH
SGbGu4jokucdv7ODIQYtFhyPNmt7X4wQW3H542EYhgxOOdz2u+Z4CVa6S5e0FtPA576v/7r3/LAl
gvt74UIscsNInZRuVHvQ6aTnRepGbKWKGzrZiU8vBxBKzEH0qNM+lBwJVOwIoLJeQsgxBmW5tQ54
6E5s6BsUCJwe2rIH6E8Fr+8QHp8Ta3gcrkqbPLFSWXdEQhKDhUzSUQ+rS1Ak642uYmWpfyOTNsEZ
aTYno/ChBIf0lP4ksWDSg4gLZI3vA6w0o0ua9i6YkORQjAqo18jjwR615RoN6jnMHH6uTHu/5+7Y
M350SLsY6XZ0hfX8pgHRKjNiQuf1y6c41Cnqp9Vz2A+ChEcFMsWa8CYa7rbUAZvpDAROW+58MvOj
WT4FwbVkq2CILAxrY1GRdgj/Cq7UwKM+4+oqNe0h+yP6JN3/P2uU00I6+h/ZqzHETQluClek8rSz
v9MWNSWbC2U7UflYEXdKK6PJLPmu3Fvk5pr0BcDUn4AmiMdL+ND3TMTsTXlfc0mCehy3GTcly3eP
w4lgk1JhYqCj3q9PS4uaWIZI1mJ9vfjEgi1z/LX8tkwkAbcXSjezu2iaDlP9peFT8q/bt6sNYSvJ
q56FKdPgZpq7W+VFlmoiLstRGbczn+CnFJ2Hhlx2O7OjTg+MODyjLmIFv18IgCW+qddXcRt3TUe3
/0iErrn6WM6V6gJ7SiQxAh/7GM2mHWeUCRQdfbQ0Q8TQ0OhPCBBb8+//p8mf6FN2c2DsxfuSZszs
Lb4cfCmNwTrc5Xgrmd91CPl6qiFMNkkM6mFIGC03koqtnqOv8e9f9CWiThHSpSFc2w7UhL9U6rsQ
DYql1e2OGw4G+tbXZJp+JTj5Hb30llK1YRUL+Wvy47+xbMWUMbigHooTArMkcCBVbNKL6KqFteLP
1xPY/hCMoAZ1x/nC4LWd7ZjIru5aRKKopzIsa3SFz7tC2gYUpIjBhUqxCYiP41ZSvMmo8tS28EVN
/GNTYfFkX4IV51u4qh7P5ObW3MOhFx0JZ3X3hCKZKVrV+jM0pMTic4ein5V8MSP6eDlWmbMRSwA9
i7tsV+xRvSKW4P5tN4pj3YKTuxBgAydPUU368SrLRCb1C+fi2CPQDP4m4Mk0/jOfVZ9CwNe3V9nl
To49nc9GWuN6arWa+QjERJbuPmmVMXXtQO+XMRy4IX9ouZQbTjCCgQhhvx8DLWSmgST0GTWGS+h/
xbk6XGxzKmBeY23cb9ZKR9iqyElPFk+VlRF1VZLHfvwMSFLgn8IPpaTmt4dpr1QOvlJz05uD0POo
3TmR1rbhBHxCOiXuFmDaOpeCt9JEUa5RnuDANjq3E2VG3u77uY3vMqCOUlErGkPYECOTg/MCaoCJ
79OCW5VIKCVB2OHv/Lh/7g1B+jaaOtpCfVLRB7oPapFUR2fkJiweTkDsYnTI3ydNgA4+5yYobsxh
Dgwa76GJ3jIbA/XsKf0UyzaK2bxc6uyHB9GI8dr2pl7oy/fDnZdYZeZjEkyjELngg13UtO3Zdkt4
wC5er0K7gsVguvu5+i9DhV6qHyxz3p6TKJulVzzu0mr4fo48ThzgU1/fuut3PyHv/hbRGakIj0Yl
MTq3dG7oopxp+4eNpyajYfn1aLawJ9ssk3CNggpHMtT+7OG2j9KDXLux3wVlD/KF9VcAYJzYoI6t
N5n6kD0nhKoaEMEE11vPtFcMTL/Lnbq54deC0Xt4xNcxeA9AKVSHtQYP2IWWW2ctJ1hvem/CekUC
poFm43Y3C/wEdX+J6wHbpqUc5yJxuSwnk7LKmCCcgDUcSKWj5eQjIfJWD7gUKTdkiGrEQIGSV+Pn
EYKANUjyMv/em6rOeZZ1K1z9+B1sLd3/G2qVnZWaoFFtC1Q3pdpNO+5pcFmlkXI1kfxr5HS2iHft
m5yVoNgGZacagOcI2YT3rOsrE3Su77QEdbJUl7wHKIktFEbHhBapohMZChya8plRJhyu9SiI3UTu
yBrpPpOS2apFrhyTcjMFmNIcaNDUOm3o2rkpaBNuH6syld53eLX3Lo0cx7WEoHLJglx8LfAlc42x
hlcL5VTvuHL3xPqlMm2pi1KyXpyIv/3PZbuqpiKh8lP7THav5hU9osbQfGj8H9XkgXbQP1h+N3wT
CiezdY36tBFJpISiMxT+MNLRILEbqX6pa7SKs65SrOpJ0V795moOhbJ3G650LHGae5XiI7fe6UEt
R/5whs8GxgxFnqEPnV0Mb4VR4nswXijUd52aRCtE0lGMN19xa9xPAvdQg+SXLKqo7XDxQ3FEHXQd
YUtLjN71CKPA2ZcVRAImD9AUetc29RoFDwMuMX1pH419jY/4vkSf3RSaLfXZ1hedhA1JNlNxGSEF
y0PaL5MtoJm54cIrANTNFKyhe8+FvYbx7y82jFB603IbVgyyC3/ZZsWaCtK4PdP96dDFyC1IfnhU
c4DewDa0/G3Le/n3qnwlMG04MqySjNyvyihBc3kWzpJj8lsAEopt47KqtufAB1oeX8bfFQnMLEAb
asb0eEkY+GQLG3WxSbvT5CCdIhXEWakw56eC4FipDuXaUt3Mke8rrmrJYGRcCALmp7pTNxdmyCIh
MGyJTlDnBxGvZO2OTk1UNz0WY6sT/jQwpIO3kRUi1so57duTfm/y9SlAw4WH9LiPROyPnVdTfoxl
AIbH1rdwVdBtF5NkI6baJsY1HdXP7IXVontXVcc6vGbfSb1l+7ecIM6KcZ96v3sT1An/YDQKh8nK
8AenwjDaGJEho1kNBRpjrKs0rSxwx7EtUs6XLrKXtG/92LeqoXswXPdQePtzzlDAytS2frAHJrkX
nMm6eQr54EFt4cyGsAy9/xZ87SM61a+28xfy77xXJWgcphR74H/V98qT6/ZBSVuBZrjtaBTKzuU3
LIbtUzvsztI3uLIz/tbyS8npeMlx4hd67Ijtj/fYKeYrXbgI96v8vvQkJPdxIdCi3u+RGkbA1mAh
gZbIraKqNfttfKWB8hzK9m5NgpAp6Zzrk/WmpsK+8Uz5OyUr13Zx/guPCKxe+xMludi/V5wMsx0S
w0FRkhDk67hzvOxbM3m89VdyrAY+pQhKtH1tHviyvfhbtYZe2svxFisegS/a5a+6DfbO3ly1Srpn
ihKGRpZa21jVF+UlAkXPJZEQSb3ugCdPHIcg8YPuiEEJHJeiUrL3KKjEr4gtEfC6+kEhOKZu6Dz3
Leo8yn0K2y77aC8maKg4BkNUREU1NBmPmIJvTMMy+0hZJf3D3tW5K83IHL7GNMf7a4KKsXVbQpDc
re6fETRJ+bswQavrIr4axgpkMPU+yUJgSabi7Gz/KPDvDydZue1U10rPJbvgY1jsuX9R3hzuUJAs
PbnfWLkDcTjSU5fGA7OzGLbYPSKPznnmoLc901OkdPV9Um6mzSConVzpcxQSzp0xoZA2suc7yY05
/bBDfh6ggTVIbfPqGmaTNuyL6dl5UM+eiXIZ3I3/rMob9ssuOwln0lPHk6xLrnfxsdeyi2y4pOXL
wI2IA0brGtA6JBCRZIx7MIYaZU53Mv7IttNe4weyP0bLcd5WApVDYXVhqK+/r7zl+8NWSZpzempu
C0bYhdDxYWMdegWd0SzFJYDXt1yLKdG2dy/W1O0oEnTeTTRZ2PnOS/bQJ30qwbGYQvzSrWxe+mDJ
ftuQvutLOQQoPMBThxKDafznh9quE8XHfi3hcKUGELr2IWuRSwQFiHfU/RgS+NC0Z0UlZJW1G36E
Gyc8TvvsGCFkKcWauOwuENlXrHQNxkW9cxhawztKMj9/a5aQivf7aP9aamZrcbq+NjqfnvDqG3mu
jw2RlbkHWHmSvHRht3Rkl58EBIpRoGe74+avTZ318gAa92XTYIwP+qd10gHNAwFky6nVJZ5+MBl4
P4jHI4KEtsaHwe6Vyf8BRU8sSOWXEGDa4GRUGT6SkyinTQttEilVugzjF3EJxCp0voD18S3Buviv
x5qHGG4qXOhad+sPzxVL0GylFjWuf+SNgWOH6cFPn+9AsKrNcDyOqugz6k53lJ2K9a3GjtIN5/BD
WztvkqgmmHWE2j0OWk/MCZvRTbgW8k3vgwYNWUnxec2bEdXiTJXpv3jOBeg30V44h+thX6iI8/Ed
XWGmFgigiZWyrrNIOHj3SenggeudLT6beDrPZSPc/3skvJilPTDIUR9GrlBK4dH2iU47fjRKL7rH
un2g+bc77PQ5xhkVvlyK3BI/qP5raPLv/xWqYGl3U8oXPa4ArEltGaIXjBIf4MO8EkmORHsYEEbL
M9RssqTBxSzlhoXcoDb+DLBo1tdyooq2d4bvWDP5zEz+6zilOeKmSaXW2KlQVl+i2KzRAbX47dIq
DtRes1crGi3yN8EYtmJMRSPe2Ykfe9nOpVGvLFoL9NmsXX7B2LxWol6ty9wOchnRmXPNYiFOBVXM
xf/avnrzsh70mZrJjwrRDFTQvZqUxk004IvNzD9SEF7UDKOWqjTNZm23RpJndItSFeC2cOXz6j67
aMTEamL5Yc0jwXLkQvxLsaCwVzZVQL8Sv2dRKyRfxG1VZarDPs547h48QTBXt/RZQQA7UNtr1iMs
Tl5gPLllPxbxX1zJsTqr/m6xD9G7MUXHNm6VVMySj+L1aKnuGfb7CGffNmuMzMbZPTXn4K5mghQx
cbUKrOU2mK9mfs0sYPLCDmrGYWlyHFas8iHhzl67QIas+ZsYsqI4PDjd/oEd+IND9jv9atv84wva
AiWPazxiaiN0JLbqTFqbiANDIuWVJyDr73q3ok6mmHjylKnxIuIS/7CZm6iATqByohIKpln32Nl0
66AWyyqYPfGeBNZLTWvwYtecgG46ztU2VthjNsN5GPdQIHs7Gn2OHDVzcbgzhRR6ZkTrviwdG2m+
OhJXITwpW7Q9XuWKFmU0Ggn59aP27D2+RaYmUCA15gaNQSxBsGQTg5rlpoGznkpBbd9mMYbzsNto
5CqkLVMyvgq4Xxj77loklllYjiDz3k8C2DOrCsXmgNw+D+idnDFjamb7ep/yWU2OqhVQY7MqjgZI
S7y7VZDQ9hBr04IrDGhjUPQ19hJNC0Id9w6ORlTgMoOILu+XgxQx8Wop9g1X4bT9Esm+GYR/wd+7
AQoWgKPGrU/2otxwZb5xWa/+gpgYJ0LD8abclXBPpWxlBhBGmLzWzy3mG3i0uACkGlxVHud324gW
mAAG3OKt5By9xn+BIyFDYey/leFfM4fafNJLJNG9IODH9PzBdvH1hc/W1j8Nl+pAa+aXSKXIuHsZ
CGpzbgqxztnXMui13VbBM4loLNnevXmy7/eIYpqnIyxe6YPLz0pQYMM/78fqu3XUh/rH9D1TwCpi
i5Z4syCYQzMM0+eZiVVa2zq20W08aJdNB2KyRh7K8PzGYTsZSI7oPYiFpAdPvx/xtK30ri11XWlc
XtMz0jL/snx8c2ZUVkLeOUA5knZP0jKVnWJTdW+zm6Xg93bfm+Pxo9Ym1+72TKKNNr778ibN58dr
EIZbfsytHWHaHCzWLnOn3E+SahRAzayKQdyJ9Qg6aF76qtEFlwI0By75C0CGVnYDtx4kGP9Xrder
ku665Zs1kPZy75jhtW7T7tWZO8HFFsPjM1og3ZfqSrw7aTybYqgdUHt7qPKQjjjDXia7PLp23zct
67CFJKAXiBLGc+N5oOaQ7Asr7TcD0SPhtkEMIJ888rrFHXXTDMXnkNjoodI9dxSMvR6TJRyzatWI
ZIkicxePaQJdwL94U2psazqBzdMKR217j68dpycxCGxfHBjnMnp8GqTIjgggfQZGZy92Mv95CHwE
Y2RKQFHPM5N/x/w0oTvQEGtchjQq6inEHp5DhfWVk1sqvIWWH1jn+JAPtyCqzSpc/11kmQOXHR//
K7b0aE/v79Yq/WKEIkrAqtWzRUvUbc73K+nJY2Db68enS86C0i+jhpsLcUjZwwe3gt55cTL63nkG
ZQNO5zayRB3w6Mt8MAjL7uVPZwmZyyuAMIN7RT9/AbyAE7voBFVC4h/li3HMF0RluYvH0EdOHr4C
CPaMhfFZYOIpvoqaWdSlMD8x7UIBccf0+hIL2AbmMKNIlK1WCUd51fBIiVgq61rqSObfooRyNoO9
7mwCycIBxLzG/YGiW61hd8+FK4RUKG9+P3Zk+TthH31bFYJpPI5syFO3jCse46ftyrWnfmJKARPI
VckYCgxpGN8dMG+BsQaswlLq5O5DeINtp1h0PnAkASAOeyuvqWqofYBNZVfo8Gj1G/KSsvnx2jY8
Geb40ha3IlwHahRv/U++1LmcvPQrydTlDz1yY1DZldMVueUhUwNP9Uek7o9ihVfRttPGcyNOK5gy
7IDeIIyTkgRVqrOJnKXvYWmv0Zl2KGP+bhv/IqGqvLspq/MQ6mQGYkATOqe3i4X2s9+OLw9ZqGDC
zrCn5kcfTfjZ/M8u4+/X3rRfTKju7Pp+kC8HsuTdtAba03e3KxS0OHFCmMvel0Ef0nM5QhjvB2cw
0494Hl825OS2wvyNwllkdk/sIt8FzpYG5Na4/bfrVg+68FtvzL1hg5h1EqXIES6ezha++GUVeUUt
OX5/2Pu8oW4K2FLKoN2IQSy/UowaOIgMRY5F2+n0yKttKY+CfoN50eW/YgMmP5QHX8ic9Ac44VGp
rTjQ4UG2MnIcSKkWaICaDjTOJTG1JQNrIzr5eE6qJxW9ZFUSx9x7gAFuYarJSBd+Yylhwyx1cWP0
28EViu55htobKftW48LLEEsHV9sZ5DazASeYW7Fsx6MM5jf3wmPwICPI7AWh0rFxRT3Omo4b7RYi
wscS8TS9FvX/Crdp/KgAIxcRHC8BSeCyEyVInrjay9GFWML/BKmsbxcKSkFqvYpW70+FHfZGz1o4
cmq8qvTzIc3OU6PmFMx20+5y8bMlqCMTOPOzcH8bUSVtfAhb6eWZXRMvzddD3ftSvdeGxP8QcNI1
omvHRz4oD43Y/mxst1dH5Usmg/oUdPc5d6Dc8HEEZ6Lpv4muaIMp4o/LSmNh+/w8HVXC2tKg7DcM
Lr40xWD+796bekw2Cl6PS+K/47Jvjt8m6XpMCe4RK2jCvXpvHxyLTE02tJw6MVuaOI4zjqphpuzS
2/SMzkvZrP/e8aVcg06NdIjC4GqRVb0ZEeQ0f1kd9BDVHWF1CBQcod2Jkws1vMAwOsrjExRBrchi
+5qVRildDLk1NnGKvMF7F+J5dvoKprTgQovxZ/B7xKMygAnQdpjpUAms/xNwHPptV+hT7EdtCC1M
U+MS6nm0Rm6t9AKDItVEFPD3B8DGX7tQQp9aDt3CrZunKsooszWxQC5GlvsWXH8vT7NPjeujHu/U
x8qsMvvznBomPulahn+k++GeWNt+SOegBfdnySiuFsPJVQN6Rk0/7EQAgvmJkZQa4PUzU5to5/tm
KIwVaRnOuZd9glOvV9j7vTxtfkId+EvhygaiAzZ05R79t4i3bnWIdAnXElYGcvL2UDkFhnjliF8x
rFptT+KGEMf2Z+betL5xaualW6l/b2zsXZ5oqjkSuTndo2zAvN4au2zmkmxLBM9nxV2Axc9kiW9W
07gfhjY9iabsrN3YXONmtsAep56pAtF3na2gyxD9P6IKE4J50eg9+yk54NNEEYdfYqBUE8y12isd
9g1ozvrvT8IYB/Kuxy9CGJxvtgFx4NbB6ulgOcBI4JV6WVUZRj2IvtlPFcTXqBtydCEdO+b3PJQl
AbQKJnATqhlbvEdtTiXenLMtg/ayMGntPjlqeVWj858ZQ9XPnl6ee1uWUuMsAJeIIMfxNfYEzE2e
Jag0hRoj8I7AbpnQouggPsmrjCLVVCvdaaXawKX50rjmtXQ0DPnS1+Qrx6UNB401tSUNJ/GbjKQo
z5vhQikrPj3lq+WkzImsuSULhVCb9Enlb49JO/IbX6VeY4jzCOIn+40NCrt8uP79/w+8GIW95pcC
XIDNRFu31/eBKaNa2BsCwYTkQdU7cYH7p+seozZLchaYDSqVl1NMM/mwpWJlMR5LP98RLyiH/QrW
l1SYDPDPYtRD6gzloifaCzZc2Ne8tH5KmCAHzgkn3OvvOt054uaLHtSPy8brliim9yI9caOoQiZQ
3ieVooNHrB1V0agoGA3r+U70LV2GfOlsoTBJ9CQKZNx6tenyLE22eNfdyRD+f6x/uDPyuiJ2bvQx
8J4W/iFZbZJ2lnE9m6N3oOxTJw5LJK963ItbVrgGzQN4iLkksIyhtvta51fNthtnTc7MGt3eW9Ll
kj2q/8+gnTYIhQxvEqDf2reYEv0VGcIJiDWMR9q/BZCs6hZuKclWC7jTfPzlZ27TOep+WUDn76hC
HwTDRL6uFRyQxVsS3Arq8mSuFB/LIR/zmmiQtcW6lcCC6GDd8EQKn03nXZ4T470onC3S2YSS6HT2
HpVaIKPNSh7iFrSIxNDSW4zXcCZSsNESYm0AbPBgPQG0odVfAbHKrk9h8Aut90i1o9d+MP/kZCAt
AEzxfhH2Ss0stcYjQzTJygjL1229QnRrTFL0WeTpwHzajxrxD+M3e7FULNewolM9RCXX3p9lO4jJ
X5pCHWkDhnDoInhbS2xOFSGANmin0985IbATNi4YUFJFP14lkNNOpx6ET7GRpeVaYda57teny/e6
1GlWpHmfouLuzB23lpOT7zH7ZQW7PDaZ2CD7nKQXY8XIXQr5pcFNsRs7VSwZPD65/FylysogoP2G
Ru/QQZGa7bIrInTLcJ3O0NiWSVjnU9dBjjtpKhhfemAKKMJDr7TWZiBgiEN8xSvJRfr3M3qyGrUy
4kN/nty70U7kKrmsJ0R25q3JagpDRepRJGJ/RZd+XjKnBgJlFyaDIAtcLxEOZvEwsRQSlzYLol+w
bfvUiFBwKA9jBduFSk5nYOkmv+KpqUJa8krnBcTJbINhHpMDKk+x+SGhC2vee4DQXRGtMSUqG+Wu
RaaDHNbhRr7s0C8VqV6xEicKiYcdFnNXimVHjids0jNI2ZsUO3KDoS4pnZQ3qhDZ2QX3ckyacBIX
L2WpG+kiIqOtKRVWNNLW9Kd5cDxNtV1DoAaVKoBEv6+tcr+NeoSKDA+CDPNADSeVuvHYmkw+9TNu
TzrUKvHGA4iu6pu4ikZLxOmGrAVCo8yuHuJE5REebfCcCRL2U88JUSc45q9+1qXw+MUgYhT+4NAq
A6jIEWs69mgQ0wGDvRqFNEO+pWEuYeEzPj590Fij+RZNd+DpEncgifoiyPNJI6W59QDCILTrCczP
j7u2mEQfOoDpzLgiGsBQXzqa/NM1TZ7iVqmP2HBh1SH3E4apcD0qmffXkKleSaMqX+a9H33jHO9t
R8DW0lw7+ub1vwf8IaWbUuFZ86BDmloRm5PeUSLoz9YsuntwW/fWXu/cjnWIMnDPSxIKcFaNJgsV
GiJ8jr9N2tYnol3AZ5C8FSXF9HAcLXpIFgCa5EquQCTm0CVAx+CKf+9EV4NA6QWZxC1w6W4QpaHf
AZRVuGHhDYyad0yoTuUWQpONbXY4pFWKo9MCXp+Y0FEGIWaSDm+5TS/O6TSF8wxOSArMZNAKAlWm
hCypW3tIzg+2sscQu0CVpaWdo/QqRmGOKSxUEbl6hLJ3GeYbT+jZOQX0vl2khUiYG2uQgEkS9f+Z
+nPeBXaMMvMF1x1NIj4UcVTRtIHPOlPT3pHuO9/dFr0gglOhyTk7KOgjx16M11eXuPi1bfreqDX0
GjhQ2xYDjGsGAuu1CaNsnkUi+qvdNRONvz/dxQRMZGTWwV7eaGbvlh7p4YF91s/39zIZ5G8RBfuu
5I8u7Cwz1w2npGxO7H0IJm4va5Ks0lN7XtUwkkCFN7GxaJ2u+SgMnrx6kzF9AZKe1eDPH8LP/yh6
71hSSp2jmcCjRPoYYGhPJOGmxmIQWhKbQwUpMSI3XDoj4jkbvvcXyVJIK84abutTiRODxgoAehkK
53B2ofLs3JWMAxrE9vRpVirdNyjORdOtGPGO5zdVrz0Z4YaPlaSuBDDKAv3oXORHTVwcKp3tMy0n
EDxgxtlFT4AY3eU+HVXsNnAnR1zBJhYeqNyRV6QEs0GGKR1wP6z+wDoJxdJ3DD+HihCptCO2ezKF
sICJyzx753e5SQPeWO8hsHre2CNNqaREIa96e5MNnXoZoLG3mksxp8F6qaBXbkTvm7fZy6biZD8c
5gzgtYusndnCwZtvrYCpsxS5wLOHV1Hak66UMnn6ENuvav+2xwfXsznqcV5KeHWllrtyoFRMCokb
zRKHXVp4A2j8PP15L1Kdgw7yWkf/2qSO5YcuAYJgtHVxUNVqcxRF/jkx+gDiySGFJjhRP07JbR8O
fA8s76ENjZmFJLdzTdfjXsOf8TZyW2ySnmpDLPo6/+Rru+vuKbOdy8yOHSi4eYPBzg+tzRNEpCMJ
Hjzg9iZ013jkCFLKRdDMsm/tB9JVz0EjLY6hIvvd2v/TMX0OoSzwGnP0B2mkKJspm5E39wUZyPgq
2qhVruqgCAegDHwKcur8PWSxhSZGmXvYOyTNpSJUQ9ZBO+r0ElNKNjoprJGfCGFm5HfFyImasvKK
/dPO6odcm8yVCq5SFUIFKC1aW8idORo1DP31cQSpdTTIVHIw/fLxTzGu4bxkmIyVhVdnPGOjgKEc
jM2TKhHvJ2g0I0ufl+G9R7QBn99EQG7k8SDn7nLN3NHtwAFaG4fYLKnh3SFKX1TbZTZteH0OH4Ql
+RD4GCrVWyP62qnXk1zBmay2eI5vLl43oHyOoB6HBZu/VMINxs7r/vc5zCu+ZjC0GcJK3QZepq+L
1b5W52i610Yc0/MUdOW6C2S0fXknowxolghb6y+V6V1r7pAdlQ9hGgC2yrEtHIX/zd9N4eoKKw/m
lmoIC8eoYAdAyzdcko8vtALJ7dAwIRXbjm3+XIu4TJ4pJXkJGb8dL5oUtSLjxri9CsI/tvOu6FvP
2Lr0KriRHXTGe8WyvZLCvY96+REC/a6kbracxj5Lk+Ac90RnGIHfr6NN8KDhWIqqr2w3iVlCFM4s
HCAHaYCv3kTxN7AYa3Tow/b/XSaQ1P6ootCDsdS1Ma7ohMIeKI1QwUTfrZl49ggqfCP4v9DhhRJ9
a4FB0k7Ln49m5lRu1PhCBtQ2e/aZRfLsnJdMX60Q+X7s4CRu1gK0d7IwO6j2XTGd+X602DkY0Cdq
knoPjV8gq8IpuLOBeMSGwxx4sTjx6zna7tZPi9CQaP16j802cA5AsDMG9tdc84jkD60m6Y8iI0Pb
FqPheoVRie57EQsBXFueB2h1FrjTNVjFBTn/pTX3Z+vZmIJInXN9erM2NyUCvnFNfg+uGVRexUKR
shRP23QqcfT9ut4zaXIIM3Gl2Tgno99y7ismnvewNZ2z83UVKUkXWimhcf2MDWmw17ildFmDxCRa
YVsnv6GeZwyy/cSCFD+PMxgZ59ma7TSjQflvkP9dzNm0CngYHY7hrLFVhMVir8NWBpgk3D91ZOWP
EkcEh2sAY1Lu7QbawMCrMKaDc7IWdfwDBTT+bdozV1zW+vuGkWJCfV5Pb/ksfUHE6PafH55YHf/F
fGJMnakYeYq9A8xmDKYurV/j2AWruXlj4Ri00KBVumM+FOz6eHuonIsOewWdLdZi7/Q2rShbgsiB
lPxPFNa8QNPv1vXprNJHsWgYtFacNDS64CYIiCHhAsyhOp+TaMa8hrhOoadrN7bF66CkePrgb570
4I2P/WBRkBPpqTP9dnF6U+01V/lWoH3cOCw+MOEJ3eBm+zWbmheN2Xj1ekJ6YEBW/KmKcBe31o11
CIyML+5+t82VShKKJhP690gTphLkrlFhY010h5ce2AVCxtFEzugq+jAkaIcFGs08R8mGRjC5uqG7
EEPlAhLecTsSRcUsP7cZkoEGJrGUQOj1p5xQ3dGySEFwrI10J/DZQT6mFSV6XaKoXZZPK1ZwujKp
TceCmbyAOUXYEhn+EK9NalWQRgRX7fXWyxz9FAL1bSwQO2asXM8iMzv3FigtJCfF/wi/O5CgvIDD
eMbnXfS0WHJqDz4UacrgeAnF6Lnt+v7cM/vy3m8SXlxwQvzG53kf9/P1KnygFWcndpWba31I1DlM
YhjipBIB06ssIDOt6JdF2w8TEUODejPOFx5TVLB044ozb8qWt6XRrrmfc5W29BOzpUfVX6V/SPBP
XpwO75evFCETmtgDasGfqDr1n9RBHxlIZ31gG5TepgLmURDvm8r63U1KEQgYwqIVX/AaVRNhs1Ue
eZPmmGgdzfkEDBab0KivRilQvhRgiK0VUsm7vPEOUlbMVPlDEuw6ZQpWM6yVTE98K5ibs9HloskK
p5wfVrx2yM4UxB2iKxfwEPPmDq/bJEWDooI/VIM3gVa3EeaYpO28qav9m/c/rzPCuIkYvl2O3G3Y
ofMHP7QT5YME0oyHL0LZF0JwAvwPxqWwEnpCiIxlUaV3HwY91/ZNayNNEaZGD+q2ITf5g3rhRqWd
0+ht+vqRILj9baX2TgBBF7PiEGm7ZwfuY7ydroFmRuObvXU25N1zY3rSwUDsaVelVq6V0INHvVBY
OHdqWrIuot5sMhm7H4CWKdUfSwugMyYUyQFzJWhYywsCIyH/2n33Ilc31OhAZO3Jey74V1OtzUeD
rssjUjAoKipcpb4tzOW9GVze1cjk+vN218XAqvrYsiuw6griz+FbEcscgxkYi/rtNW6mjTyBaAUI
fD3mPfYaVZzQpGnpA/XC8aff+EEqoBecxSePWSoJpkFiaxz+fMtOYCiFjycfeLa95eDTYxFJjmoK
xIQd0XT2A94cGJjI3t5SF3bjpl/cBkUV9nrWQD4Cj4RhvpNvoxv51sgf62QlQblYaYKxe2zHvYDG
2kfvaEeNwal9nNB4bAr9pXmcuHiD4bv2ob+7vM8u+kpH8152M+t5VshOoJN5ockzQa80SA7RppsP
ufuw4U7ImLpdji/US2kdUSsaHJ3sc5o5Hw8kwuYlr1xZxa5YtN86kOObSKKSdBEvRrb7eaLS8BWF
iWv2rpwQDN3bh18LSuh2Wp5yuibauQrXPMdhvx+4SqJT3fsKRlCr4oJxTYlftNjC4BwZucZHbnSF
17HTlpgt1CpttzWajwYoyITOqugG3/5Lgt7otE3Fc7lN9fI/u7edzQG2aCNOfBsk/7kk5g4k3svZ
JmpO4eJsGNeeBTUTEzuhvDTDS4IXBpb0jAYLhjp7Whq3bPaWUklcENZ33hRkr84XCNc7T1O2FybX
bhY6AC1hItDkMBE9GjjarGNxZFrFSOQWwC9pir7Qrv0Kq//j9+IkMe5bUgh5u5Lp/8JqinTTRzPA
wF80CJ6jP8DtkhB/DqWFfDbPeJqs5KYYxkuHjYXS1AZHl0FHJFnuRXQrEnvzesKOuWYAgHNPG5Y9
Up1b1STGtn1Byr7hnSOm2iT6g7BJe0O4Z1rQj8JwEdcB8Kky7a5RPvycmzpSZNnLbn5o/smBYH0H
qcJ1EKheArW7M7t46q6vh9bROd07Pj2+XJ1o1q/2D57Sssg0rU9XsMz0pwqMIbKCYellc8cr8GAZ
WzcjA1NIZsjajX6x/PqhpymZWd8bli7ZK6riF51bVUeBEj4OZ3yfs6K10214wzkrZzlj1/ZhK/AH
PqXxxtn/t5C9Ce5+ArYW+s0c8Fc0Q4gkI3B7KLe0v1B3KG0vGIsQXzd7A96tYVinvCE/xmRAb/rS
R0//TZsSmHzuXUCbuZ1HWwOfRPdv6Q0HB4Eb5roR1RY6AnWL62NWtyVdn6B51ZCSLcLd1aRQC/aU
Auq1cor6/q9a110fWAbCgXDhc7Cybw6TySur3HplzSPg3sP9xXge1GGc+3lbj9XfSjInX4uls5wT
2HYSeHuEuz4Y4MLezmATYeNcY4AmCvm1j9dFgRWkX2iWHwX41UlsVGII4CcJh6Uv84XE7BKcDm+Y
KjeO5dFy9bJJuOF8fzg+KIF9khkBhtDOo+B5o9MLEixtkSr9KDdTLzJTBqi2GzVWBpbGc97Z7a3t
GmlF1xc89uSL85MxXIMMKx8joXpOMpESnfsEmb0lLHfoCPz4DeJrp20CyRqduubdVwx14DLDStIq
WoO1stfrvPSSaKpDFgpMclqqr1aUv9qi0DH+mtj2Wfd5oIDDVjDZVE4yKiH5JCJNxkf66JTAl0rH
lAVmLadMmyNr86HGe+NNFEnUL6j0Kx9QkA+RH2bSE7UwtwXzHUzvpvG8559L5aXxygcnKaWoNkjC
vpLvVZlinHFLuqdfzQuBNNkM3gFMpapHwzEXQMqqV5MS+kJMN7/CEY4CvvZCvVVz78QfifFF92k9
5a2L6qTMRpG/sanN/v551Lg+SM4ZeAyCb1oKhokXm39bwFY6nqem/Rlc5iB0tyZP2gLtDUrsQhMD
oY96/rEBY9N3zrHjTqoXBW5SLKt//S1BqH6Y8REnnj7NctE2iyCkJhvxZxGnZxzDM9jpHLGQ8GKM
GxtW+h5+a8Adh7F8SVvoYXIZuwPiwYtoS4I74oWc1YbQk+SJESsBY/9dVvr9LVeBfypEXk6zTznj
5xRzIQgM6A2MYXC+8q6yE3SNGUn+KtGv5AVbP1AA7dlleeJ0WdwPzrjs6Yc3sNYaMPtngps0UyfG
f79huTnRtBpW3C07iv7o2noBnihCx3H/dKtaDLCMKGIeRXNJXPBAXKKNZp6wIQkja7pSs700zXa9
jU+vio/RuLXCW6oeSeGdthAyCAHllAeIL7ORtuYcmcrooNpSrmeha66/sfGPUaLsITIbEyzdEs4n
NbcooYEgjKR0WRCLFodFW4wHqcxK9WGb4PDa4GfLVdRmtz/1tvl3R1fViYdGhaG3iaKgfXcXD4st
14f/JNiXeBa+g/w2PZr8nsj9aRqszhNpaUgf/PKwyUMp8O8DYVkJOMgWcU8685KinN48R1jdIMA2
LJ5fmAT5e3yKgi6rcN74tOFOcwXpDgoONxF5UhRhn72sqfNEibUULbOQn4IqiUKsR9MdaEXbU1kI
IxltJjwS3R9O9eVDNIPeufoswiH+E9nmveS2U1PL5AWYJ9HOt+32LzSdCBnxezkZg1GuQzKMkFqC
nVaLa0rQ9fPOQXoIj29atH0Hzcq7E6jST9uz4sNaevRrWNK6kYGkAWduL6yAt+AWPgZilGFxqGkc
1H3v1Tnhdqr52lZatfHuRhcC6Krr0tAykOZNZB7q0/6DGtaFEpPfKBaCBhiV+rKOzQR7E+1QSZbf
A8gumxG+aEMPlbfxwaKfEpa2DnH2+hgM+hi3IKCIzP8l4pVCGdBXUzOm49cEKWve0sc750GXEypN
hsPkofltEDPERIN1cbiZlXGo4zB7nCl4LwddiCNpVssaw3SaU+HsQa4E9k8kRT50wkgeJImWsOtj
06J2TQ0REER8uJFHjM4ZKcJ6SJxD9TSs2KHC9ZXypoRtuDFt2AkMz7RnEm/rdIcOQhrhzUFoanaI
XU2xWAe0oTolViMDFyrlxxKB71wPH1tYyyiMnVCop4tmaMfByyq8Qqh1ZwmiOK5bh9xF5lCTDA+8
mSFxr+28Gr/8FAEalzlCpPWg0aEWVy9JY6+nJMZb7z/xIJkrCXbRw0Uoh0j5y4I88/4h6VLFHT0Z
LNtC9GFnoQUAh6bC55KWfVfcnfu91vOnql/4Hs+ADPm8lhFS80d6HCAfwGSnWo10wNnQUphHaRkR
9NyzUZN6YX85h935mlmsWNGPu38ZpeGbgj8AabJgLjbj47zuz9gFmrsxqbUixqb2TZC8M09HHias
htUCP+qGEwn+JJlwpwQTegPEY6SX8LSQTHeV1dmYLX7eGyiWdaPMPf4q/ZNqC3HBS1w34HM9LY8L
md3PL6jQ8UVFNtm5Gku9kEnv7Cs9dRdOnZIanXRCMgGpWIoiXGJhUbuMkBmYv55xnKxbOZbZ/tse
+83E6ynzLdxJYkQ1xG+JshFn3p7HmnE58pIPW5ZWhBfvoudxPjiS0bs/qZecpGgeztqDtx0OcFFB
A13XZr8xojzMe547hzOn6u6FNeqqkINTcOV+oH4dfWSecH2RQdDWt9IGTOc8VTfW66q4qrfnHlgh
hRRNoSdfTmi2LBjDQ0nZ91EKLbW4tHIQgutuwP7Hytqv/djmquEaVs6+OGNKZeOJ6TTxTL/TUzhQ
pm+mKrlCtmWlJ1bL45t6r5eC87eXAa7/w6ksLsGNZrffY1lKEYi8b41+XQswSAliKaVcdx0J00So
tGu8xfCbgMxfchC7ka7G86ehpxpPBjXv5QezpKLSJW0UstUAcha4n0ofxqK76yhV8Udk3dx84pNl
vW397WIzONDVExXxDXb6lcFGPvMaXmg421VFeeQGjYwH32TqvIwT9AkCp4wi9PpwzuOhCRVUPtNG
k3ehKir2Aoq+6ed9CzISnK6/KS3+4jIcF8PH2FTfCGq3oqAr0BBo0GN6wjhSEgeiZ6THf7al2LHb
P6hxZ/Ivg/PCXa59RQRTtRAACd+kysyUl3vgQqkpv6tQpzQodPMF9s+s8WgBfg/HXjgpwC4ysG0E
BHO4lnXQgx8oZnzINVonOwfNGDsYIN1LOtnAK7zCXmrys7XcAvnrp/c2GFbOlD1ZOOyOtNWhQWnZ
RRpV2gDkJjpv97i5lbTQssrYQhNvL6rl13nWxyWORXnnqbekxAVBwFvMDyn+U2cpOUTrqgZRQWxh
rMCdVH0vojvgdg4s7Hpo/kQSj6BXFZukaQac2Yp0PIGKQUwV5DnyhX5Vn3//VerD0qaFYO40Eu6O
puo6lbd6SL0l5Y9YlwXv0C/8WNONi1KSaXTs4q2B2jkFbd4zGzdFFiUvNX12io1CaATTgXTnqOca
b7/vjGpG/kxz6AIRcnDW8/8P2vo0KyDuXA51k3zoEUzvsxShg78TrhqS/P4poL/6SUN3RPiQBdpi
19YSxfpT4DXrplfwP3yYE0RvKtuSpPWtiw9T6/q8QJS+bDH+jqMPTdF0H2TOb9yDbxllo4V2iD6Y
Vifw5h2rDWYZ7RgTnEykEMjSp6S8R+eQWMrM7rNg+wlnJSuxURXOovj/gpcXnTezLNq6k0kASa74
AaUd/MmTav7mYf0L/fR2kiolru+LHKziUOFndLjWc7yfq+ioZ3B6r9X7fKC5zxxqzEQNKK8rnLjH
6J+mndGHlfmvEAaHi0qW6chEg1++Sv8Y6GBdSzNnUhXFxnndxxDVWC5Xgf0B69pEUlsRSrso9K80
5JW3T7hM/vB5FqmVn+dwXb2ueGl+n3m4nRlJIoPe9UZ5U8HqbftZhCUgcqUUf26QVGS+aQQn9XU2
sDFXcpcM48EiSg/gwSySzUAbxncW7VX8c3+H52zZ9BtEXOHByuVx6x79/XUMlKCaI0fDjKVJ2pac
h4jDiG+rsoNw0EbqWMDGNE39f3VkK8K7sRH8uZw/1ix148KamSMyFEQ8QtOxvCDN5bTsNtoO1VRv
zQJfIwuvVJvbBHl48gi/FvpmFvSIeS2qtQ3ahSU3Vpa1/A4yTf4TIeWM9zcjN/GGf067A0liqcDb
A8e9r6S3TGl5Y5hStk6NX+weSj4+cgGKZ9qH3qhGfSGj72atoeGDVwksAHnvyphw7YqX2xQjXOWM
bdJnysPvucoODhf9t5YtOKrlgN3FYVnQ6tiWMwIAra1nuAUMLfAMi8qnoGedecx5ESDvHEDEUH2/
fdAzW7sq9vZnOHtimL9CynPPBsn4HDDRHwlOtJGnRR1R1otbGtG6dTtyuYdqtaW0dJ8yRpTv10wi
jlFGIsqeJlrFWyAmXG2MMn9VhxgDT3hNo9ThU0qGiiq5ouH3SDuKlqRL6ZcOwEL05Sh4TV24q3w2
8/KcRwgEwEcavdgQHk1pXH3Uyp3rAgloNtag8mybzyqaVRvoBGLndsPsr6XlGT74QPNx6IMqVx0w
U5EwwZYIeNQeOdY/5p0oD4hYfOBYu1a6DrSIDN8zdY9g2aoqxegLfbM7RMW+qe9z9AP51QYQOYRl
FId4LT4UYJKVv7HDAach21NivUcTPFf2o6EFS54NOW73cXqNBA5kd+6AB/k/VteSp+DcXkPKs6u5
+abO45E5usTEYcghGr7kp8Ey0mQLJWFTlARq9kwKa3cQ19ONFk01L64Cg5NEbP36UnMbIfw6M7xi
dyg3w/2nq6/LAkm70z622qGSIMSYeMPxC37cAY3/eBpAuK8ISf2jI//GgE5CQvRhkxt/CtGTD9z6
HWQ5974N4uj8oyKBvxqMYzjGOfHzKTRVioefvIEF8AiF+03YBJ/sxvtDGbOzUrZKlrreYAtUuQAO
n3cu1V8CQ7YEmt1WmLspXaA6RH92d/aLRWBtRX0R58bXnsKSDQ70M8sOWu2BmmgulTIT32w/GOfa
5zaGLs9ni7mAO+zjsgxVFZHXWVJ/meqk3c1bJAM7Z+zXTrZV/DbJDPzzpcuRW2Nz7CBIW3RDQUYt
fUTYmpJ4H05Nonub5wo/1IgmYAs11qayickmmNvswCeRPxNBW9dpmC6p99iRJRQTdM6ZMEmOg+ON
iRzRiaABcFmgHcnkcatdzF3b+8dag+KzKYhYl3zLGZqw2KScFfwzcarq9FhKWrE/A5nhd3uAejBk
UiZfjNLhsTIs2IwUlexaz1XfG/UQgznXGomF3gmJzJKN4hQaEZiPxtr6zEgDsk1UwFCdqrCiFDZ2
KYWJFFdU9N96DA7AnouzycL1NkmVUk37aMAbITah8V+qE4izW3JxqygDec2JzP72bZzVb838EBCj
3NzWzvYO7IBDuUlOXZ1A2DpKT9L93L4r1JoZhMeCTJ5vK/ureoIyb4V2Xl7rq7IKkEiZ7EqqQ28f
+EpPRGCi6ImsfBy5PNqebg0ylZjlCDDNi5zbjp4K2yfrgxkbqxqz5rNzEa8rQNlHPepbcZJ2jGIf
bzCMfF3mUhnTHSYol5cMKrolG+xAWOS4ltVo9unTUE9WwFjSeBvT9Z/x2EFcorHZqpAI0kaaRtWf
NsbnA++Hm1s4oS6z3ZreTOW1TaKEagxqo05yXcY1SB2n2Fwz7KfbiFXsDSnX7H4BGeEFqiLpljPv
xUbdEyhoL9b0ZyFmgXflPuNyE7ONf8M8ahU8Dd2Jbv4YdcK3TPLVG3i3C+J+ENtCOeTfZETHbjhK
vXDD/7cuqpbw3KIBRFupi//lBUJ1WPWKJNTkVHpDc2vujZYvHJE+BsxLFVkD5YxpqLbzKEC5KfYW
E6uuko/cD3D2Mi1MUdtAGT0mrZT3IhNF8n9EeG8yhHfwvDnAzcZrxhdHp4Kvh9GO4wNO0Y8GJQu8
p9lOork55UhEMRrCDD1MQP/oGMqgCKslZXGlXmgIZUuqNagPW8llchhTEuTniESPXVqp3aUbSmhl
4RpmV2YQ0qBwjBesMmKC09/XfqCuhW9tvv79Dyy1+1VRzsTvK3rGcCRctUj4IfJ8svJZ5zyGeJw5
UVtDauy3iBEmRXXTbRSKG8Qtt2TmatI2ra0coWZpgSTpsp8OwMZgnk7d3gRYhaDMQsMKtcZHdK6W
pbCHgrWYTN6TOAg6XjOA1rph8U9AvSb+XuB99O8WYPrkB6IihnVvzhRNbQXJgvNMe30/D8Gvp7vE
wUNq71MriwGpBHXzswF8Dw6oay5ys9blzHajxAZkr7lZo1GRaujYvoEmIxy59HouFnOpgH/dhVmh
i35JQK98Tp5XdxbqqSAH0IDj1exhmbQUdFUfM8dothfVGyKrVw5t2x13wIy5qzKqrxn0I2WT2hHn
gb5EYc276Iy8dQpmEb8BItbyP0zkPePlqbmqbNkz1hfw55vszxOV4thMCWyxDhPB3NUoAA4/3bgc
Z1R461r3Q4C4mt4quK9C6L3eP36Vra+B8+z+0R5XnI79ZSgBzarccEEkXuN9MsdhKk3MPMVcyHCZ
vU5vBigVStIClxnZqURtVmsAaqfB8jrUHoCUiwgxkhu3ctaJxhO9gHX26LGAGZkOIF0sB7U0LQ9R
i24yzwOogSaGm4QEPMg3wlDhGdMtTN/k3tAuVziddwSiJjDfTsEYV6vd2h8+dKhKqSmR5ARfD6/k
IXc2sPB0jsPy2lHCwcb5kYFNY3+IT2nmMt9oJ5nE4we3GmhbLOZ/f1OKkUSSyzy6dY9bSZt7UbWO
bSbagXw1EMIps2pH7++pLGwl6cxDNt81QtEDcND2qKTlxh7dVRY7KbqLFk2GmIYfrn66DJnLq7tY
Pd/Cyo7ctjIGc/YQeYXPIbwpfDrqU7Dd0P7ukmWeG23AsRWa+q0cmgac57kUqbE1neI3dHBzTdeY
cv1yhoKE7dwMxw0GxDAMxw1U7t15pDQrhrBfCLWCQjwmwqAnt5pct6hpRWw4vmrQe337+/KZINvv
8w05yi9yjFa7Pz9cl5gMnVSqZIOW/pNz/iYUS3Xo+ITt5gnuRPDIyYkpTDM8FLY4vDb4avwtQrbd
wSPVm+jBunoZ5tfqEybRa1etgq2hungX+gpcPJTcXttWCp1F3CjLsSn67X3m9SEXLcN2FWL/+x74
72DNgA4HmtE/TPP5hYX/4I3897RGb3AH3Nlrt0OL3v1NIWRXWCsmm2I8Pmdd+8x/JiENEqKLjxym
AJa7zrlXL7hc53edEx0rcv26lpMaxlCbPspaS7XORN/VuHWffmd6t0PH0+SA1jzEypzOr3w7EGUU
nn8M+MqwndYkj5Z4aY5YHVvZWy7BAwJpXiP+IR0HKy9gSdTcfSMMzZdv8y0GJ9Dh8bMTeC+Ap3ww
Wvo8/5dBA6YACPEVaY6Wx9sB24g+tRfdJgDlCVwxFSR8uIgv/1SVO6T+C615ErjB5Q0zXbi+RQuD
ztaggYmgw0YHoBfBwsO72rO+6dPyy/S4msVtyAOyaBryj/fcahC9g5ISq6pzglSTXB1iOEWIblln
HseuCU+blEwUEiVlkVcGGyvS6UpIKGjcnxr0CTnhSdY/YjMnvkqoBUgw+DcBUA9Q2WK7Wqo2h+Qc
ANr1HK30c+kjmkr3hioHMPhdkOugAUehOAt8o4voMeNNXmipKxETcZZdy1M4D2Ze5WDLtKU2Xpqd
nDBMKonxwX+FlENHLHSH4kynldnK7f1xoFQppE+setD2kPzuEuhfiF4u0bm0aGvMNrj3ubaw4Urw
mEHdQa7Wwy0JKGXDRI9KX7DmkqjGxQfvbH4qMzeHp1bhHiIsc0zFRh8q5EkJp+N9ZDGJyhl+ldYU
ggyR13KUWzk5YxNGdI8BQHH86kFRA+Cf6QOuKLYnP67t1M8T8MkVWZaQfj/n3y+50ThVahcS5Jhw
8Hi1wHPjUMFTnx8qoGtw5MdtxBXPUzoSpQCVV6P4npvOPWW1Si8Kxcka4wKOD7AAmCeSryRtGeIz
UxakFVYh/Ev84Cbmq/CFV/KDKUOcA3F969qYnl4u+HmfHDNYGg7fprGp0jBrGuKVsvNCSVRZC1Q9
WydAiIMU6RDmAbRMc1mIXXd4MCMwamaaSSrFzOnlfxBNZa8QyHFnjw85v8cMtUeDWxuj7JXT/QHJ
LOBnWVAF+mO/r2okPNGvE7C9gUAFqp3d9wOut71sOZCZn2JGfLVgRGXzRoTGwy4FQXrmx5esAjpK
b+aaV8DAAkUOTLlxx/+nIBBq0KdIM6Uuf7NrE8dy3E9V+UZQJ4luZjmS1Z/jCWNmXG2v76I+kXJW
BATNbyEvgmNwXQMkejvEMrY8oKagVQr68TfcxmoZ9SrUQgxbnHl6Ur7W0+kk1PuipBzrVP9XaU71
t2KtceAOPhIvcfj/URXKC9AjLQi1pbr2gaZNdjvHw6VtOmE5uvDINXNg93DMXJbvFIs+Fq2TLzDm
6t/CzzW6Ue2J/BbJe18MA0jlr25Z9Bfwa7TWBghV3N1/Tmzu88nK3syOM4U4n6T4sG3kLaMkhQHe
GSuybeVqBkgjEA+nTGtrF7r7MKhjimzoemPob2qCL8rDDWwQ0C3j1hM0g3p4rEgK0xU+CvNRyONa
ftPVUV7djqGw3tvu9TDK+cnD+YrMWUdACAbB+hgc4xlbYMUm6f+1+8h2cTWYM8rVC7pzlc2agSPj
CwtpYxgMfIUkLI9w79dzH24IbtOQgfQ4a6CfmCcMG75cAxSWeyQgU4G9rC8jKqb5jPzv6JuiF2SX
x4Qfg19F0VR+WimSR9kWWH653V1LhqOi62xgc0qEVVdwuHEjRFA82d0lvtGECxLBmj6nZ0c0IIqV
5BQffU6lH/G94Sbf8fEmYGLkK68QXegXTaAAGDwlHNd+VA2e5uXt6ZoAeF7UEc22Jd4hnOnFV7c/
sOtUgDBJtZ8OC/Mn4/mfA1CZrPkRCBLYJxVy8ZHhT3BjmjShitGlc5UYljxV3KyUigGvDTYtqifC
deYGq7hviUytrDulNk+11LEFe8DwUhOxnpB9DBKRVEbPQW0qQqzJ0q+K8d1gjmjVyZ2RWVnLUAMj
X3a8T8f5jFB5/PuNyhWRj0xdkvSrwv7AXJzprP8stXYr4E99ycK8CwHEWbWSN0E4T737r7tdq1gn
izghxVDm6IQ+Ss1f6uQt4OI41479eddZzLrLBdGtp3YIfao8zaJOQEd38NJ+mQzTiibi15SMuVdy
+zEzLCQyn5xeV/vXrja1RG5HNXwF2AYVdaCmbEBlbP2F+XYipM7T/+Qhsht7M8PNotzztMBz0RA4
Ftbbj/mZmg2cE5BGJI5VNEFGraO70VOXkzDTDtLVt0NTpE+ts8wTU9sOJ4BdOZT9AZpGDIEnMzph
+Z+tH8Xg6X/rQFvGiK3aA7hH9yLcleODLbj/s2mWivJYTDck6u2LFU3aiOhxCy0SKdPE4BwT5mmt
rKiRjy2Mrrwj8YPZGcdX964U7RAEIiVG7X9q1D50cofnbh40tM9XC9BMfchmFyrkh1j2DKe3PX/f
5hUq/4g7y5bnMwEfxy+/8gYjmiDxpgWZiuxDRu+11tieRHK8s3IQxYLSGBf6cKBpZBobmdg+w1RR
sfBXJ7Sz315ML1HgUuuYSVdVUcG5fLk7n/VeEfeReK1QbAGF0Hef1NS6OCz1vP6O0nQQnuWczlf2
t3r6Z/KnnN1R58ZQr7gROYsYfu+9rRS576gfBaiCzB45R9tUKd9KPeDhaPPNL1TAt54rg5qlRE/z
k07xCvfnCDtoY70sCkPozX6+l3CRVN+RBImqSuYdVfpiDOHZ2JL19E7AbcoMckXAC5AILcPrvrtp
b6N7UE6CsYfmARt0YMDI4520Hv+ZB/NwiEs2sKbd7X/GPoRlQDKy/+gpWWQ8Ik9piU55OsW3q9Gp
+FZEJ8AyUmSVYuJjFWexwRKYBX0WTfYxQGI+pLH9ZHVrU5uEncGYxMk8GiA0/UBBAvMFqXb7cmGO
qOc+pldsnh+vfbutKWp5/jkSrC4qKtxZweAQLjoxowmCCiXCsy7CCwHVkbPwAVaR/I08oV9vEzKq
W78zt2pA2HlvPRMhBkGnYc7uc0TSan0nxmr32Qj5yZvw/34IlS0F2TLzisjPie9LLvRNU7hskwst
CvgdOQ9lG+2OjLz2SYJjk0NU1oFmJEejQXj2M0NIk9Xh7eDjT89kCtoOFqNLtzxIPMEG8ebwy7m9
uBodemgLgUtWGKIXeO4IUG2vqEejpJfmYor3gCjlaXptCmmuy1JlCP2KK4My9I+yPJ2pQbU27+Qh
R6dLbO+4/1hzU5VqI9ntUVFC5ITSD0YifwdKeO5wUKes2f2o0Lcg/N+fWFgSirBDHYeZm2st0AgI
mGJCrAkvCLxJ7av017K6XNArV4m5DGMel7Auuat4+4e9J1fgFaXsoADX0e3SvvONMZF2j3pT4s4q
2h7Z2QRWwIi+1SoV6XbVUjuIuoBy8jDlDnPkLb2EXWuRWYqAPqPW5bkFxALxKNEzJpY5jo7+UIS4
i6nce8YmLM5iCZROFbQB1XqdNP+zfw5mz+Eti5nvZfrrXn+/sXF/3mpVWNIORf4loXQR49FmxmQn
lTb4rAphIsHV/tHCyeNNA9dtrct0iBZtAW2qm0alo2tZIYzI9BL3jlzFerz0xdS8o0WhYM/+KK+S
1/7DtH8dKQe5ZiE0YYQvJUwyf2nWBLb7qsKtWprq6WxYWfuEY0hD994CBSoseYf9xT9Q/XkOIY1i
U8TT4rQzFOu7gVbrEVIWfdcnescnuOc28AfUsmtDENcl1N74Pz2QjoRkdBmCq/5vArb+m7KvBkYQ
Flo8lXHCp69/RS/QQ6aAhGSWdIaIbGn0w5/maqA6IizKhNnHO+0nUWW/t2pTL+oYhkbTTtXDxsHY
RC0YVjIfJSPczHpD126BFVB5om7HIulqbfhsl8LWmBMqJuSuSMA7TYe01qQzLVtjuVeVEpHMccvg
hBJWqMnmbc4JN5di17kv21ogdusaoGpC92KAQfTFLNbj2fQstfGEdkC0X7I5DWHHAEGOnyBMDVhU
WMSLZsBWVhwA/h0zj/mDtbrfSKeD7QW46b41Tu9yf6cErP0jiuA2rJNCv55DU8sYidG3BNw2xSRw
sJjeC1jt68qYk4P8WDIqdqEiQvuprB5n2c/360DDQtIAcBDunxSk1eliaBK17faSZ4ljO3riZnwO
o1Ap31j4MaeaxB7d7Q/P5cNOfxjgY/x5qgi257Gqno+O2h9nE3upDRNCnfmyfBZVdVMdP5Q9ZlSt
E/JKBrCZV+NjOwq3tuSjHoiesxCCz4rqBF5+n4HY2oCU8DS/nRt3z+F2NF5pfDoGayKUVSE3NEWH
M3PQ4HcHkr3LD1Sg5YyuKeQW8VstsuEtyzl20AJIcweZQ+LRsaBtFxKCo3FBz4OqLsfUuH1k96DM
/L93xvL292ijbOaygN2kpazFCsOtF88pZs2Wf3EYHs0of9D8NTy+n/kl2YjaeH2wnxA4DcUNVUwQ
uO74NDrhjCjWTcosF9iSdKc6t7O4PXTTaO9Bestf+AWZVCzvLv5E2V6dNjaeqbOH0w5fKrbUlUPC
SbUUtxHRhYb4IQGO0azABxauyly2ZBTXBticRCLRLbFK54WLWjxImTSkIp1zOUNM4/zKNxhThFP/
TxmtpyhgJi2Mm3uZCoiHCbqf2cO5lkXsOL2rXSkFfJRrbmHI3NwAY4DDBXsVgXr+nd2NU0pBSxVB
rrwgLBTh22qW9S6XTQWNTbR30EOoYN5iUSFR5BqOXRXIQR2th8QXZTAJ1O8DmVOEUJeVx7fd5Pn2
3aPbR+Jaqsr4YkHnNPTA+i8Rdk/19hHe28mXb/yOeS8rJjUUy1br6vTM88uloFyMtbvP51+Ph7ti
5ftAQWGcMGgQdYXG4RAYmmJHYW1Qs0pZK7XsCt/sXWqINv95jEvm3jPBUUYwDveIHEGr+6rrEh15
9QYPYJPhGCesndWIneh5xtjQXkE8dTUCKS6dN4IqfMTGJ3+T+WVy0I+XA8l4hA67z5xLFzBRjJ4D
2PhBAhOz2+u+v60TeDMUHSr2wGLvAPURgE6/lXkTtSnY/kefZsDqZlkjkhPFVMnWLdL4d3Y7I/VM
1o7VaADeVQAWDtYRqsBsolfRBaQ7DzMbgqVwn9FUn54FbBeZ0lBrYleR4LFfro+8eKh7Ab4ZbKh7
qPqQe6m2tw01l+E5qXZ2tCDSISFUdSP05oXPt6hsV+72+CD6qkVg6+6q87viw91t56kRWrmo1W0t
9y3KQNcR4lPv+BVTpWDGL+sOBusdEFXKXBs5bd2izAZD++W35lM5ujIHI7zzfC+Df63g2hucyOrz
TpzeHZS74lNVRTyDxMDi+rq78aZaf1lH7Pn3be3nZWW+ibRVGAz2QZ1fe9oAAUEpMokInyPWKIfQ
WXq/zUf2yRjN7fV+WJ2rEdjPZTaOzlf7Hk6C8L2UMQzCW+JEe2FrVk/qe+uFXJXL0gF3xi0WfOsd
2fVItwJ8uUYXJh48PhW97BZ8yQtCiVIYPLmR/zIFo1aB/bB8qqXMVjouVFv9ES0SHUxA1nDjLal7
IeUQUbY8NAx3In+J1x5vK6Z+1fp6mxVOPNkpTP4ojj0IyAidM/o3mrN1FDlHSmuMwmIuYSSHYhxt
BTg3EGBJkalakGhz7V7yZIUkMmmVXL+sFe6869/tSuJHWqOzAE0PYM1Ka5S9zoBbVldJBPbIXbB5
PGiCuZbbyQWF+MVfEtpJ+Un8LEJQ8+vtuorXM46Josol2V2hpDnov7zUnGfh5gUi2Rbi99+GNOmf
A71NrL4v9rBZAz91dIEQqwH69DdHk8jLzk8PEeMjtyD0/Gifrvi20eWEBI3PPyOW6AnrGKesfuOp
XJfbT//7J5q9GInaFO2slYiRFev8NtXDC+jvxSgTX+re8UgKBb8bHM2lTPoFb88VPV9FbleeCCGI
Gfubx8BBYe4UwN5ZuUK4/ek2DuGvo+ysiPOojlHSn04+KCDy0xHJ2zr+f+qhqwQE8J/BJsFi0k7y
ur+UEbeJdvnBbDgI5hEMX7981alKLgAigN/rHLtPYzuciqQKTBDFrPb0ov824ERx87+jeWciKzvx
aHkL4TJ/i2Pj6IotbtYW6VpjpR5wtbqPPJfZvwZKlNFjsCyb79UkbRdY8eKmpbyOSsNOl/KiCXKz
vy4vr9qK6nNqqL3IN8UwrLJPd6DuoL39vh6Kw1R+ndcsFeYO3awUXtdmXSUNxBqcFViMNYnjh+kB
gmMzhMXqK4eCSw8itai854Gw4Pu5sE9bZeN2V+ancnmZ7b9KAox44zz7abYrwCngtpRD6obLe6/y
zl6dcNdMk/B55RMmok059iR7pNmBpAjz1Cs26stSUOo5j1EcUqSn3qKEVi53l5gj6JpefK6tpIQt
HK3yBzKeArenFpRrDG88BRpgdSFGxQdOps4/+RSW0ewnqNoQVE4VHbVsdVqHTLDOhT+DNVfPD06Y
9+h6kJ0CxLifFUgFb2Lyx/JxBsBFZEEozg0jweiS8GkE2D2ta+b66YdA5nmMLvJwWpxa9qQU5eLv
6JvdmtknNdYUgmeKurRPxm6bs7sPfz/ipA03BXs11XzwO9liZGz2Nw1nNf0+BLCS3yoFeh4j987S
jThEfu/YqImJv0fabBKdAT+tGbgtYRC+R0tX6rnW4JTCT0+NUEJqn64yGx/F8c0HJ6mK+R2AKVpI
2P546gebruDWOG2Qi8zS706wb9Xr6eXKQf7AzU4kYeO7Mr3T5ew2Z8mahAWHhto/fug1PNKPH4gW
MdhghZ9Fj6IXoV8N1hlAD+0wuO+eUrtDapuogC8I9cPfdmU0+fF1yFWzplQ04mCD+jHNlN4Z6m1J
uJAHkI2tpFcwlu+y/xHfqxG/Q/vCot2nUCF2PnKHDsl3JemBxc1yAGKUdhV1Mz6SQ0MQ1oE3d/jJ
baQORyGKUIrcrU44Wx54bQ/j420X7yA+oDvdSbvQWmLQanl6dkABMNVIGqKc3tB5iJcyJ0JXsZn9
E2qRBzhZeFDkSIFxD6g32qPHDokypyCEfMJ22uU8NVX/fOOqLjLqkKTGCTB9FVKdg5Llv4qqcrf7
CXDK381AY3h5dU6rRcH+QD7i48rOrCzQ0nAkplmDaelJB76HUHGH5Y8hZYQA7n5tfb4VkAHVM+2M
xDCeyt0IFqkmS2eV5xOTUEe0iC4xKx1QzY7IIBJHMLavxmBCauCn+X8pPxXx59wHoViFQ4AxB/ZW
r4uva4p8tHjdULjhkrCR8gVJweO80EPTbVNOH6qnle+TdD0B0B47Ue0HSLfwMoXtadTB2PmKXMrV
ulnp+4zFTTSNh6QdNzEiyVqratHYjd+d62g56Qb9gjYCFzPOeC/facIfazblu/dDbyAgIEGoIjif
VOQhSznzs+hTOW7zYscQbU00NXAjFT+X5mbcGStOhCyLVhomnYXa8TddKlOaee0YfXoDuMmg/Ezb
AsfqMw43Hm0I+hdddVdIHGT7+NjgVVmYIn636jEZ7Przxn/L2nWppoUkQCwlfumcbVA6QNIutqtn
l716IMgDeVN1quHUSP3jbbZP6lMpB2pSxgumkdCDaim00zPrWFRcxMHI3Z96sXd4X4H7RU7B6vEZ
EYj4n3z76Qpa/XgaORs3Oxt1pmknym1DbmZzsPTlHxeoEMmzGDI4wEUCW9ZgerNRfrpFXpHxJAib
ZCrnwkR1TjZ3/RvMASelhJmZywhYn5IrJXo9qJ/O/Oq5p21g9Syg6/VYlhg8w5FRa91uaOmykeoh
2j5gyEcu/HoqcfxggZCSGaw11cFJIOkSgCHK3BXwSlKteS0b2+2LrWSMdv/75obpKq4XMt3GxBvJ
7gVg617NhQC5L9vl6gNLmhbG1omtKX+hUv544UQnLbSYssHwGRi9ZNiaGm+fqP1RtVryCDq8p/Gs
hevDwMlhDaVzOmtSE0yPkA/6th+/M5IOLccAZPNIFNyFHi92i7cKHoA0hKwIS3993zuOQRCKWPuN
KNUfAUO9cbm0n4R/SP0tM5JcyFayD4bXq+iCWkqb1AlRg6YsB83q51OSN5Hd247/HPufn7szvKwV
jcU5/LaZOikRungMZm7T+bV0t4wk2H3YDfdwu8g9M0GHSnlNKoq6MiOH8efT/9uwlDylcukIHS9a
GWL5BQQmsZxrSzvp51ybXWLwr21mTuqe9ohiLWRGGhs4uwnLoQ8m4JELzsDJl9j+SedbCOQn4kHe
RRBiekHoZT0T/Dx/kGKvUhsiLkfs3XWnnK0qGNf9HMBJEBJ4p7p7Fpg9Ju3WpxCBioeJWKREO2/W
s1LxVjWgw5VPAskBErcMvPVtc0Q371P5ABTjCv2H4XLB0JDWpeRb6s2p6YxNsgrINeR8F37/wNzz
Zpkfn7cOKmhxbUJ9vYbVz3/XqLgdTq7n4yr9UkoiU6g9Lc0xMu5z1rR4q5yIx3dcL5V1iZtus7UY
MyxBh+cpiyNZLUNU/QRs73502MBTjfSIA3K/TPYeS0PdElB4axPyO4CCaQSJfKE32XU9QOlWsfnM
+YyUUG9B22taquEy7OB/oS4t0zDa7Sj6AicTchy/6lNrIS1+rkWYUDh3cUArTM7tdmvYvWUaJ1ja
e1cbmsnLd5c/ar54Y8Wj/a4mXKUZMPvFK2PE1ldFm0GdihaA0TfyaJdZc1vQCZ0gFIqlSLc4wwpR
T02sgm6onJKOzCcRXHYCD3NpdXjv5hz43j67pPztJn/3c4x4ke45KH7WXPdD7351iPgykL5Y/ezM
XjkqLi3XxEVZwgzZhCisXmmwsyq555KNxK4mwqVn7IdIbYQ4UNPjHr65XeBsFh5IMnaSCk0v/ndt
fNUXpudrV1cG2t39CdWM/34cCmEjISUrXNMlWbhsRGi/o1qOHk/0GQP+48buCsQ/VRQ8Mz1/F7Ex
G4OUiKhXqbf6toMgi9r05bCteLV6RSxTPwJxpSrfjo59NrMdC3fCXZz0ZiTNnF94rTdCQ55nWkc0
jflSlG7jssCFTrSv8f0AnbIJSLyrsVAcHtGzESP033RmSoTBbTNTHoc7ibJTtCPDME+fWBUkwW70
sRI1ET3CLiJ7B33a643kH8DjXM6hYNJah3rq3t/vt1kObG4Pui0cXrNN5nXooqg3DO8ktkfZyx1/
JRV/joVvIMbs2/yHldjbwJ8fnuPpNLcXvNGnbmrxJWjNFVk6Hj6bxyxE6clRLtrUOiDUZmry4qdw
I+9kJXcmhE2JcgB2kLGCShcQ8UNBWdcUIE/VWbPw0PPr/Bbx1LswJuehTaommzPD/4z2NbG55K2d
76apqVDdE+NvaX9a/8m/rXV16AQI1EJmQ4odrl8l+wbSgJ57XdML2bH6Ik6zaUX96uPtmHnj6BAv
I9ZORF9HJMv/hkHosDjKb3fYtIX9a+tLRdoeeJqKQY67pk7c+MJAikrd7aPx0rnQAnBSnKlzOWYS
2mcfPEBZh4lPIJVOnV2391d0zznDO/AlMvMcO6C9kLFVJPV8uwuus6d4iHXVQHOKkEBVZtB+iy8k
wIB0YLa0Ly3mk0QDqOGFm45935aq9dCoKhYSbjYQiuV49aJDleYOBvZxT6pWtyPGjfqy/XZl88+T
pYUCDOJXhEozUFaapyKO5HnKr3DL6X/3p2FT8jQA7M7avty5rApSvIRybtxkWVTjR86jsnvwdMH/
pC+40xEKC5KhiIk81oe50yV7nm0DvbhISO3Hhrfv6Rjd6PLBe8nsmTaTdD1OwxRp/3Kyvjgxa20m
ZvtBL4WberdXG6a8M+Cm85GeMeFcZB0NzU3v3KHviEw8h1748d61ySiZaZzaHzU9VgUY35Zzk8Np
/O6WgIYy338SyCLnBncndArkf6IOAlwahatRs87E1n8o7bzR8K9lgMtR9cK+9VsqVXW9wYcJDq/n
jJBkbG7j9aCupLxkYPm0yhHJ4wdYN+WngjRuOUikf7f0Jcv/1B9a1zXlzOklqUXgw37AbrlSDvaS
Ccwes+J/oQcjFixoQGjRWzmPU6qmCqKfNuXXY/31U5+r9HYpQFa5vARGA0217S3AiG8P0YANyRwX
lB4/BDgVt2+TdX/VWXWL0pZZv4XnOWvgGwZx2xOm5e3ZCgfixgE7dBPW80UnskHHalf7bpttEExS
ytFtee3HsRppruYE/jdlpb4Ut5IBihil3gaFDUcc4lVAL/yseYZ2gERivVlzYIPAVQJ0AJUHOKfc
XkABH6xgKtoS2SxZ/GrC0b+0X/gGLy3RIo/6I02IyKYRWa8jHeTBBhrZLqqSketHOfbWQ/wHjYLX
AZEnP4+3ilPE/Th5Wd31PQu+2f7yL5sgKs+b8VlNGeCZ1xymijrX6P6pyCw5Jgzecw2ifjxTZ5ip
NQtPfsTrL5jSQIidf6thXhP531CFCjjfJ4OQ6od95bKO2DY4VrlhnFk4VpGfY6loO00DZX86bT7p
vd1ap8LbtO/+5REsLl4bviPnc22tKaZQCh9EL8ioyezJw2zPjyR+PdglFwnAiOCcrl7WzwrHK9ak
lJkftLMGdkPwFw726+Sw1LwbZC+3//juS/mdbG/NgEyGwleW3Ufyw7QStqRSwMnoBoInziysy8CN
GJkML1pYDo2PNSVoO+8luvyqZ0fXKs2WBPBPIDTpoVsg50MThi4QYHF1+IIXysBSFo2N2Jo9AuRN
dXWb71gglK+sneix+Z5feQCewrrC5JOqE9hSdRAkpg0Fossopo2NczZ7o2GQUYCn9iS3cR+iSPJ2
HmnaCob+UIuAxPn1Rz58DaPbkUczknFXYwUsa7YMuAXaougBLoKQKT36QxAK6h61RuXY/5CslZyf
2taMUUgpmrsAg5iunT91eENQ3+WAsvn3/ScCO/0NKqo8Nh9pmmlpnYFCQbPtaTif9XDVPxUWWZKM
tpfqZPsd30c9suq37q41HwU44MVHVL4uL0sFiaGO19RYumZZMGn45smLtWPEQYsQXwhl6m0yaCvE
dniIP5wDA/IUzrGiZ5mBKmk1ERsWGwIACgLZm892T1anFACve96Q5721XKIE1nfUOWGs05OB+SOz
BM8FEMEaJOJ6bEXjqmqK1R5m7ogDal+dlLg1UyhtI26ksoOMPZJ/BReJEiIImqZoSqBa/VdLYp5Q
ZmHfCQXFPuqTLpOenpLFLa2ITrXdFQkJcyadA14Z6gWALQrCAa0RLoSj3Vlvdk0xwwjKhxknBX10
ZtM37KtncN/7F0T27dHf5s+NT642+/sTDXdgqRp9tqc0kPJlNYeeF240cMjlv9oJtQII1qgHrBTD
WJluSkoIgAuQ8yybjXyUFsVI13jGaXFWUuMtThh2up9CB8Y7205c6PQAdyLxJOBe3sB7BR8CJJf7
zQS5yY792o7WoXq069YpW807iMsUwMZX3vdjJg6k0r0cuBR3cCRFEZMYIRajE6dPrqVDvGpJMk+B
oWEsy5wmOYxJGIAQWQ1GUI7UkVyl+HR/eX7H2+yK3Mx/Et6KLBYw9YmSq4i+tKONjVX8A2Q10E7q
xleFTCDGHfsjiVr5m87r5aiR1cjvXoNPmQtwdghuN4qq1zRgJPEM7+3QK5yyFOPbr71wyFgHcjnx
a1Qvf1p8ZlYmpc4VXJSzqPe9fErUTNLmeRQ4LNifX22XuN3iBHCxi6fw9RrMqCKJeGP0bKahvJN9
P6t8RKXdx9nA5PGtmOYGHsgFRxL9NXSbChsdYpalemoGtgXdQvSdYMpYY+PbGcdW3kr8n1bha//F
n9xkqgfq1rqkcYzgEwU5K5ua80H7ZRd9iPWpGRLMOfngUtgoBZ1vIHVhpBEXz9vkiUb1bWRR/wrv
cnMfTn2hz9fGQpkMKrTmavckzPe1ziu9FBAy2Z5GYTUknXTRAa0Qnc2I+x2RUcNb2EZ2xSBmXe/u
sJhjn7+HQh20KCeR5u3gB2roAr3dK399vMqGDrMMdmBhBxXkpeHeFo506Fc5304wbIn9w1lrz45n
pawCcJPpyXFHy5IS3yQuMJD4iJNVncQ2ZpDnTitIPjuStASiIFl5ldSTcwaTTZDMLFwNtAex9/3/
LNKOcZ/kU66hOdo8F3rfHvx3B8eogc95PApx7QkLXzqUb/31jcU2aH9HINIyUld0tjj0w0jQDCCo
2yfzDaf75aPbbVjlVNM6+wnsh4eOwX27z3RuIne98peFNnlr1Dtr3xDfKe2oSfqB6TTjsYlV7m/s
0/j/MyFPyEpd2Yxt09qbl2yMpP31KG71nKITclVLYVgZw46dd6yKxjLR2n3RliFm/kGXIA73FVyj
dwTe1IqqtyNy0Klpk7OizApx62LYU/gmkQw9COLsfLW63EOC/mLSROth+cM+H7KXw4YIZV6mYG5f
f8txEAZ+xjME9N6qTihKiD33xblPEc3n/HhQBb9kpWY30MNatpwgxK21VqapFd4/2qqETYk+UH5h
WW27OJhKZo2P/lww6UIDpyNbKh3ttcg7PUf0b6sY6TKzruyi6QmNH78M8/RUbYxLi+meN8x5iJ+g
GYH+ynWLd3WycnfE2r9BGd1xcu1YxJgT+wkC8jIG7DAJUnPl6MFidHrlEwg897fyEtVxIZOA/O3y
vqsKOZXL7NyH00Wu+KXOysloRpoVVK8VhiwdInIY3ksJ7LV3PtJON9P+7UnBKcN/OKPyoXe6SaJ5
ZGhB3Kob4KmHQt2YqpUOn+C/01i3fKe859Or+8gDijf/cJtRGEpeswoXB0Vms6bGABKVszceHQ8b
jF25+tnHlYnjtkem5OcQBIMueMGhNtx2DVVB67Y040GaEdXNL8gJQsN90FmrQYjV3xWW/jM5ha5T
SX+NoQZZjkFQWXDai9Udpzm/fQoIN/CxlaNI5mbUCjhRptHOht3MM+iTxt7sCKw8y8TXcqIUqpH9
mr5koezPDUGLR7vlG48MY4Mp3g3bBmxV+fR/Uk5UPFNlu7Pwt+2UgFGaA/rd1p5vhkFWCmHmvdvw
oMmNBIc0r0LiJhRc/FG9VhOO/kS669E/ooC7TDVV0kOP+fWTirFRJ4TUs35oM5X7tctNBQBhSNES
r+7c+7ewdWvH/w38zQxQzTHXw8SyjSQyJyVL+zI1H0uNknCEq153hxjsDTslUrUJyRSbZK4taO8Q
8G4eM5FZ4gMhxzPzhc9cf7ra9ZCFUhKUf9yN96pdqpVK4tiTdd+jf8Sjv0rLT+ipsG994JN/YYby
fogb8QY1gyeEIiT4jyV91K4bEtwYtB6MxE99r/YcMZgIIZ8H0SiZLXeVcXcRgGMjiSSlXXXwqjuG
T118iLfuVCIreZ65HDv0SK/7XAkKdOOn5qz6yH7oY+Xp3cgkDFzfnMLuGCEVJ8h0rImAMFf2QXSU
CrjvYC+S+vnLA8vtT/nv4D+AbGq0gV4C2Qd9lZN/hkZUZgLbz2/EmM00or20liAAWGojNzw8Z9vm
z0jbQ/89CvtEgU02GzN+aXT9ROFxNHGId/ivhmDEwAyXiTS/GXxsF4nSe02kizsfrolcxm9QcTkF
0a/arzqKqfHepgzB01dNHYuNQu20rLKpEufORnba3tImFBssYccZ8X5DXzyyikZtEClC17z5sIeY
fn9pdSMZQj7ltWeSxR6I77eIjiF+6ZMa0omOMMMRkJ3zne3k1XxFCenjtAU9LrIN6K4TemuxrVnN
UX8GNSd5QW4MtB2pylaStDUAEkOueaYTcis/k8D+kTg5777af6m9pSDcOGXD9PlAIlZ9COsOdlCb
RIw1qpRcp93Ft/zT3cA98Uex9wtu+OeQ8x8XLNYxs44RWHiZyWwIodgTlLWF1hNUsTyhfVFXwf6D
RHUo9nU/yoEFEKSanH/BwzKxgOapwF2duw0hmPV/H/UpFhkwh4oDX/TTQBy4PMQ8JW9f6M8rYjGS
QkTJOM7wHZzA2wsOJ+a7VEx9HgVqIZl/9PfMkXk+7TGkmm4iKVHCtof2jnYvzX+HxoTOa6FfdBIL
O+46SbrqVqCdPyhP6ETwXlc/UQn9/Nf1BDgJb0U/GUA4IzwsMpdqJJhfTD07xhk7kDL84qs4C07f
tPu1epniRS/xEI9h0/M+VAy853NUJyUCPYAFyR9gqB824P3n8jCLaAPuq2QV51PO0aUk/MLee08r
fIzf8IpGEsMI0iwoP72FbzrNordFhTfQjHXH50QqtIZs2fCGhin3G/SJbDWU1YgG2mubONbQufwh
I/1lFj4o0Ej2JwxJVsJ4iEFu4+5IFCt1MDW+T3N0DkN7mt29H3KUUbyQdlnENd0s1h9xZDmtDBDF
UEsyT2PriITVsASklTsCenhlFjwdC0lDoSpP4NRS2tjuZ4GSwDESxJYtiibmCbOCSTpT3dsBw6p8
Dk5JAi6j1rJRNkQF7hKawAXR5blm0HGjgLZsH3LkFegR5xzk3zujdQAZSVgS6w4uzPk76MsJ5nmy
DUqrpxx8Kmtk5l9pQ8JEa6+kLzdyBEFBHKSL6vGKFo970nuBvKZcb6HFMXPHf7RwWCrdh0h30bZ6
yHhPlxBYH1E+DGpGPBfxPhXBYA6bdr5KAWFFDB5Sh9EwT1qRpchHD3G01qbiHH40uJQ6baq7fMl+
SG3/fpoRzth/8dM/Odfyqhk2zlsho3yRoSXhoOWH2M36Og/wKwdkD9NyV9gp2DF9k0AhGvfuEtwP
d5e03SJQMUzxRx1vXpxVzGGI6ulGAAyd+4t5ExI/WJVgOplxBO+J5n7vtNA4lc7YV/7bvsxMWORi
x8APOenz1hnFaPs0XckeMJmRyzrjP4rrlukZX0x94pDvmfU52ql/Xgw0rYzt520WP52vk+2jTe2P
ka4vszj2AmLuyjv99BI48DKn5C3bMHvnl4NmBo5PrEXd+mJq8EDHXWOvXt7xDZotkPizYh7inBP2
oafxoP3h8rqUofsfeVuHJGqz2lAXTTyCHmHZUjV910Osm2K94jEOmJF+Jm0D3n4W2B2tf/uufrkY
cC7Ikg3BOhUE+Qu8o286hyTY9Gvz/xg2Kr5j7cJlBZm+I363sZpU3LT3LafGN0IUVXL84g5ho6ny
pyEyIREeRS5Gg0TefgLFkXvQN5tN/pr9Sq3VgYksmwjEzqu5hk1qpQ40VnMYLUyav1Z+Uz4k1fL1
m101LMtCNn7TaDvVE7Z1oRlo0BIohf8/fIXAhRZFtCB2Cqr+Jo2N2KT9ux6CSduZJlJ80SDoKEdP
/AC8UxOEVjKkQB2ycBKwiDVztUav12itCLvkoAOqALQ4yK+r+MCAUqPvxwbR/qp0Nlpocn7Usf1h
9FkyDK5qZtNXatBAn+gGUh+PDw4b+dv+6X5cFfFV4icYyxcGXgwmvhyMDIsJie6Lp+O97YriGOhy
f+vWym/22bIpGlkWgYTbR1txdKnJQSjVevOZ8bKF7nHn8x98E1UEJs891L7dr3S7vFp1iDZhqqzE
nNEP/JGmUJXnpkeBuNpsHJcJPKmfX3oWMr/RsH1tyCLEqdrUrlZXdJYExGNZxGapp+ytmPxBlFg/
f6XvDWlygwASDVfPfjZCoKb+zVn0Xv+5EWLuxBvXyfaUvQDxlsFsuiAjm1470/a99MLiEOJcZM9g
jRPbQLGBcWdG6kPnVJcdVDOj139U2ACIh77Gtdwz1zQwmwYc0quvzg5AeP1gpo8y2YJbMXJ6O4HU
+oWXS1PrI+NOzuBOinBx/Vrqu1pz2/p7ypBt8gYTQLM92QWWqi3U8f+fdf4FBd3Ebvsh/plTOGRp
L3tbUZ91COXPgSVyIWcooOPdpT5oJKRpNWWQV3cVmH9wfm3BQ7cdLRd6k+0KtpmpRNiSY+QTaWs+
yD6anyKSnsed1OBbYQAqNt+Njq7s3vuYYRtI3vCcCBI3/VpZttZ6MoJxP/H/FeeOpt611gHvj8Xi
hg0Me7rAi+xsBBmKI82xjwf4RlmCab1aZxoVkHN3iPY2C8BMBgOtFm4F4O3/8pL6ePWs65AHv9cG
R90GUgNahgqqGjaItb9jw/wcsUDO+7ErNvpjEPpcWuoSEhdKLIkunnftYp84DWBB8DYOxYi8uzRj
Z38RzHcxOHOpTJk3bZNgnf/fCZtwQlWhVf+Y2JFLRchH+cBdebmhE9NL1GRoEyG2qUC8Q7dgjAoc
C3JSCnTU0cNmWGS8Cu5OS9lYqKF8vOJZRt69QOwCR3d7hXYmHA7bvplV0wmiEgZI3S+ekH205ZzV
KCUEZHiscAPT8a56llvtiACShZzoeVmczAm6Ku1x5qBjiSN45c83DdLj/JKJf6SyLZTnsV6AAlnd
i7GoV9g2ifrnJlk7dGZSQCTtC6qJyiXfaRp9YDSXG5N0FqAnW3d8cVnIvAF/M/+4sRSqebhBe0To
tBs9mIl4/r+diGJCsvGUGAtOlP66FxSUF18oT0rm7X63JTxYkhMTcqbH+Lc+cc4daQJo1HYdIHeu
vDMc64qzw1+HH7apsfA6KEL4jpkXo9/2m5hPdQY78KO3MGMVItcip7SVST9m8oUfBZzFoTgZVP0V
MtAdIA9Gs3WQLoUBXESdygFEFxZP99JupuCDGIIYYlKc0TUO0FguESDivW/BBNIAT2h2sfhOllN+
Wc8tC4HSOBZrhzXnJpzmEs/R4sFPjrjXF4/l1W7q4lzSqHzW7/NoCqh0ZCdX8eCnwM6IlQjmt0iz
ocdbpurpLKva9FLCZCBNamk66FcBL1e6ZMuXomapQQgG0XCGLqdrh2jZlznB0jSvW4L1uhTY/klK
6Zz07HIVp4aEDU3JV/Y/HCVrsedvfEv/MfTWM+XWMzLW8c8mRQ4t4F9sV9pfmMvzKp/h6P1UCR9y
HiMRyxg0FJdKMgqHVkhP5TTd2yOufyDjohJp4+OatfWSqmjL7FyMqxaLmHKyijq2QKjEzSdltJg1
/Gker+CutOexV/lr4tDdVfJWtmNjJxbrNCyEynnL8itM0CbwD0yzXea902VQVdyEEB+cm+CD9eUK
kqtHaHshk6M5q1KvmEaj+nei7xvbBxmsix6Nl7+3aiMGMEIlNiA8LQkhqahncETaogo+5oaR5swe
Zmb5CI/3/uzEnaYawu/GlVyFe4TbGZyDXqG7KI+s9+9fUmve2o2GOkIk3tHf60G3W8GV1KSBdq7/
HM3p4U+ITMNd58C3xGypT62CRb/3+XSQMMhDZHXXZnzut5DX+n66CUWbvf7fSYmSf8k2qxhnSLkQ
Uzdy9OoBzGZXzgOgq/+SRKuap7CTxzGUZM8c3TXTDXRE2kcaDp/LtcECXKpOuvIoUl1dtm80q2Z2
TjQ2M8684zC6+ZaRVZN+eDqd8RdUgUlXqirVs/j2XfD7Jf0IeERCkVCxYUv+srzKIe5lDEH8Kvsl
FOkZxiTPMv8/yjLgh6MBmrG0mJFILlQWAkvzh0et91xEvDlIKLXcbVHOtyQCUV3R1ooy6fxFRCUX
zXZtI90X99WVAaLgqDGlGNi2oQBPCpXxQLdePpJ2viaapI6nr0tO/07fcmJaofiVApFGKE2qGIPl
XS9wWRqnLFPfbAR//eU0oAV3/zeNskmsEOn2TaGER/AHknsNpXLVjpA/UeQh6qXQZSmBLnRbMGmY
kHNZrQWvSLmUhMDyZR7U2JOZq/w3g0238KBSFUcVliZT9FyBalpQtz+FGq3nw3o7A7d70cbGppGj
UgrwIO88PvevtcZeXRzWXdvI2F/55zgzffaxWzp5EVU/7Dm4yy0y2czjUpXF4mE7VIXPhJzNGUWK
Lt1873wMEg5U6BYIEssMIH/VrNwcVzA57/unFLQPrm6UD3D4x24q29zOeRm1qj9UtVY95xrymQaZ
8JH9d8tL7cL5jx2RpfMXc/SFRIv+nCXZaZePL1Gd0RWWOeVVBXNIIddpAslcfQJVlm3n3VkpybMd
maaU6Mniz56n1yRZALWgDZgt0/k2mMsaUhdv8jp8BTxJIN44nuajQLCZooUV72dpZ1BvmebrTb2c
FiRxTl9pj1fiLzPLemd9ZKtsVF3beJ1wZgS3KQsMUBs8rijn44/3k+tUMJkH6zAKJZO6jV8/nA7M
gjxjOeutMEyfg50K9EXGmURBlUy7/g2yoQeRyEjIvjKsaw8RvFDoJSjUg9aeW7MWLYwhyBKRiNWI
EsYexsyDSJaDP0/axw911h/7pDGwFGmYg4xC1SxJnqYHg3cec5EULUOb9oiZfDewUx03qwz6kbe7
QjFE5D19sslsM9lhhRuZcNI4FYK+Gbe1jAuFt/PO94vcuVXO17M1eFpkO95MEm6pf5zgkPl7Dbea
SlYi39qixOl/+bFL3dEK3z2l7/OxOrWXPIwEVfAWK8AF6Jd8/yK1WIp7VYWtPCKhbDFMrRWvdtOg
pTMtUQaFIdZEkrY/a4K9YQwpFEgrcaJmkIapkcmqJ2NIHiaWRXBnL/OCq3l22Ft9E2rAqw+RK2ko
SYyJZ6jPSJMamr2zSYhhAf+6S4KaACMBGKIcs7/sTd1r4Xk4gXOQTmHVs6n0LN4zerRkFJWLFen7
Nc+I/Ysj0CzDk5pH151gQuG12f7uGL3NHloQ3fdKfJd0UCzVkYm3y0ILrCHfkTVdEZMLhlPbHgw/
mzv3DtmQrWi3xcSJNieh4is0h7ZfKhLJA1fFQAuPov0H0Qwg7gyEb/MKTMu42vrDS1X0QlbgrZDs
FSAsCrOu173msZO7URZpEGZRqCzSgS6+X+lLELUHfjf/UNw1xks92mTxmwCuRP0RB49amC7nAS+A
jIJXkWvuWtGugydq5kGjdJZGCRKnS5YNqurdCe/OROzOfreZXPhVQv6T1cXWdm6U5MZ34XZ9G3XH
3qoK/SaoNEkQ9Fm4dqNb1j2nuIjojElHjfiL+GJQ8E8hsSwdi1rHPbb5tcuek9N2BCEzZ3nAPrWt
fAqk2iXPaUoa7N9Mm3Bvfk+vnyPyhZk5aWmqLLPhKHFSAAzvUUdBoqSJAhGMK9KFomlo0gnG/81o
S4rM52FpXKB6gcMNiPFCQEguTQpZNaTJzOVq2mDZUIjPSY23gSTkX4CsFDPOfSeXZGsDu9k1pu4H
/xlvPwI3FPb5WIkBH620VlU6w+AxEY/drmPYLtbD1KCgVmenguf0JX4mWZ/Vgnn5gr/xGFBgRd/r
37fO9v5bkqYkxCAQca8/xP9BPJTGrMwl31GElMcPLbs/IQhgS0u4olyRigDwShvlRdT356m+be4q
deQgPTOzS5+Kk1ISWCtNwy2tcWQg9Pq0VBBZ1a6jmMO0/FAr84UCDEGumt+BD2ioztt1ZzG+mBAh
6vE2WL5uWDTp/eJ879pv++/VtDSXmAiVBxUnbOhQrYBvl2SXp2jXwZ6hZdrIBvzS/3FQKbKFHPmJ
zAvYzRi19G8W786oBtEixLxxGeUEPX0OZUZm4W/obksU2Av5nHm8gT2Q5AE6NtYsgVYpGM2DPzJM
jqOrdUcoMFefjuJcUuV5MBdk4U6sdNDituUlnZ1yMI4Whvt0eiEiDNKZMxvKEz1CqHiJkbXojDWO
ql4D4FrpUKu+/ZTQLROdADcjggzItNdvyhi0qjwuMchqJ9LqHtZA/1NpKIPYYZE7bVO0gs7Gp6fV
cr8NCZW3U5487Kj2tYMT8tcHynh7irQ6bEqhFekcEXQCeCFr1NXNoC0Gl9to9zNk3iRp0bejMs+g
Fh852Q4uA2YmrB9s2BaszMSWYOshMK0StKYpu/NABciRMgy24olS7pIV9ETYr5se16WNSwWuWEUS
KqNMB6IvPYGLJvDDNGZSzdQ4yWr1Mrlrr2/91bJBjUhoFWFNRIt7HzI/gc3UqlVIw9S582KF1oxK
1+SItx7KqJMjjDzb0rpgZFRayLQ4GaINR/hM22XXPoXxKu3sqDzbAWt8k66Dqm7l/236NYKEgygp
br5yEwpnMftHs47EDaC9ozUaUPDu/rT9DV6tjNC9PJy9wR6DgZeVcLmvGKXCKfTifWIpreggSmXe
8Ce+jW33qhTWA78JsUG0WBsCQOQFrvIq4CUQ/2qT8xwhmig9d0Nd4Fl7OqWqKmM/XPDGoLlDR/JW
UBcqqZWrwoRpKVnLigadjA0NfT5A9PThUx+YNoSGEsPZHhAwt8Qw8vq6ANCM1OvEBu080CoJe8D9
+Bs7j2yGEnAfM0CMkvs9kqT+YOc9TJAMvuGB6vO6nwb5pT38wbVO2M8ozRwQPAxPfJoxYFtkjsBh
xOfeuqKIZInwWEjTtHHTpSjNBTcrDlhhK/l/EC4Yg8JzKxw2TgH7sx/9fUJ1JPVj0wIrubgoMA/J
4iwo0VgtgIAuDpK7r967uPa4F6cNzD83SpetoBEmO2OlTNgtXBugxTdlSnFzvQcfRT6oivnP5FFp
ampc1CLlfjtSnXu1d2Q8CzVGo0Y36mVPH99Xm47CRx/YgL92WcnU4aTKKLzC/MmTg0Jwo04u+toQ
oD82g3aFfjdMi8TBIK+nXDWs9DC0Gjch05IeABvu2QJKmbgQBWB858pBcO4MlCcqQJqV9Ay5PDmr
XyFwcB85TjO6HwnWe3fRzrUPP9P0UjLYLRI9VELQyh+r5vpIDdPH7fm2DjvidP/UDFSVq8FSQw+j
1GphzN4cehLMtzkXHdD+ab73nErr8I3Q8aUfgwoSfoRE++982GCSiZoB052dASh6Wdoo8/6hxGVi
GsTsOQ/P/OKR6kASbhzQaEob3im7xGflgocX4ZqViFijpTd8kZ8yJz9ePt+bYz396JEiQXCDBROI
g0kbKNcvexqigI1kZaLbzz8VCuh0x7B37yjudq6JCz9qcivUx6USxi+E3RnMvG77X9hG5038mLjT
2StQgxcMIblUk/jYpSbDCd28s5qrub0vFYqxblEkoZ8OTRce0XVKYSA3mj/Ueu2+lXr2/VVaVJtr
BDC0YbjzSFuFIapB4fAhgcenl4UVDKc6PDTRBP5UPr59dF+UHyWBQOvUqp6x1IVrEjsC6WmfLpIH
psUGqQ1SlQ2i+F/ZfBfb6Sna9FO8akB1vuhtaaZJJ+HXLicP0WaXnS1/mdjhZP1uFCQMXrj2ee3a
JHYNZoAVi8J3SWpV5ing6j+7/2NFz70vnER7TZMHg4vs+PprywSrNhOkYFuzy/vPzuYk9gMwNcPZ
QgAL4Qc3t3/9aMZ4+02j4cqG/nviXvLmJ8bP6aVBVnmr1CpJ7DvA5oAwEfLG08uAJor5lewQ41ax
McE15HVCqThsvJAhKntCJlnMQiCnbp/vsS7kN7B49GtNHM4X5kXtalt0xxdrGuAY/qHoR+7Tk1aJ
9jl3k8Dag43h/DmZnLf+sq1hnflE/J/gbV0oI0abKe9gPfPU3nc5vvwXnZENRd08cEl7Zuvk/Mtz
rBMw0xB94y0Wl4rdokrc/w3nPmsjR9dcAGvsW4Yi+IinIn2OICDteU75SKohQkkSdVPB7KxK8QoK
P8kjKHJJ2F8tIbEq0g2QXIRoZuyBBzKnRkAW8wKqW+w2qdlsB4hO/PCOXlwcEGUv2ypFPrzscLhI
y5ignMhuw5IriTAYVYz85vz1ZcYb5TpMMaoJHX0r2Ja3Xhw/ir6YfwRqvutWxHzwnamwrJdory6l
l+Ta6IVdpO/1i7fJus1JhsKxMi5oJa8/vB618dGyXxaoj7wqfi+lPS6n2Gzv3Y82ix2i4yTHmONh
F9kY9RAkwuj9/ZTkiTflra/Kk6FPL6/Isu+diZzzB32Yk2r5edxuNbpKfx07tHgIp/hmYQ80BvOP
GAtU1404K9pqg+o1xkph9b9ZT1Tfe+3b7cvtZ6zJ03lnO02dK0G9hOsWveC3gwJlsBqio0ZfVx9E
dArMHAbCmd+6+OA42y0A07JFGSYxSy7hjA7mAqocyl9nblerP2aEKf/2ROuPrgSlF2ONnTwmY4Sn
qPmysGukA6KbDUx62KH11z3ugPWSCFnVdcNwn9ZUaRQakJ3R++UFiU7R2iPvjyEKLAPzFYbSB5oT
dSc2z+8Rbj1RJNK1xUXUb97TRiHHdaOPbfgAdWysk70SOmeEpOBCD+c1x6N4x6e5xZf72gSxF/Br
EYpKo11wKEiUodQJg007Jj4vELcInTpxAIY/iO/lfWailJ6C2N2MQG1VYwLhtj0+Ntx7tDxfAaTc
eMoFEEfWmtigB9mBkavxkB5Wj2ulS7+12l/czQO2Z8mQz9+xmYPvqltODf1smRVk0SwDDcQjfsx/
MnHebpS9kcTopyGFFl65sQaTvJTD2wxhW4Awxfh8bZDP9k3ljgeHrAPxkLUmZjjAdtVNixxpHiYC
DiNANn1Cg96spU3Uxl0K0DlBTxIg7E9WaON10MXdKxabN1sLMcMkVlLTCxLKLfxYr/C6s0ePfg7O
PUuTLZRQwlw7eYLxNW7goXbSyYmVxx9gpf0+j2PdiX/5s78QpbjX8N/SvNw6CpcYD1+oMD4tKgzS
z6dCNKUqmxozbD77K8Ce999n0hpxEt8nealtHj2z8F63U6YswFNxrSRyecWjGGBAkRGpfuhTo/Zs
MwJrTfjeTeFFPg7OEa7lhAq2Tuyr/mc43nkIoGC9tKmD8RZkVRZbcyASicDVr+bwcmOc255+w1fj
LnIBub2zn9862EkDbLiwUOEbGAr8+jszWLnCMs/X18DOtzCPTsFjTEh1MjjcXDhM/ymnTnKNehw6
FrXiP6BLScZfImNPjCQhwDxLolalbHh7qCmLT/+KOeJdcbThwpBOLoZgGWcaNKFk+Qu1Am/Lb149
IVEevWWJUWJs3CYgLtxGdC4+mFS9QIRDUOfaSoY18MIPLzmpKyyZubDuAfM350GVKI3Rob7kplG2
HjldRr//bJIgflAs1uX4GkgNDXrg32R81bIcyd7lvB0RugG+YZsqRvrKMCYWr3fAapK0OsL2MzN3
WFDx7gNkMQYtOfxnHVCIn6K2E0XypuLhOJL/cffYH3ZEl7xdow4U/fZrUFKLpJP3VhywrGxHv839
NZkm6V1OY012Q/fW6gIJfIZxPZSYMUhUkrT1yTAPmWXckdoOk67gwnQfSt3Tsxl9/ZeCklbWDJA4
eYa4s3J1dsmpl+MeNVRvGtuBK8EPMd9/dvnBMiOSQ6QENUDPEUidFHvz2vBMQki3uY/qtooJZGpI
vjQbFEEnGAgGULu0GErgsRP2xnzZJOOYPRzDxKJgp3lo1YxArjRtKUAGvkUGjj+MCeMQR10bs33G
+opUi2Be1bqkFtipGdPT2I85IOOVsejFw9Fc3c6j+OsMtSZ+FzkOpjGhS1NPeuHmy2ms8RsisaH+
+2QzKR3MkAmHjLYPbHi1UEyz1opO0wNkP/NHOYnLBvFNQVbKWEiJTtjRBl4ntXrawS5DbjioSVmN
fYFg7iE28O3/NE1RIbkdl99I1BPj9p7uR6jhJdMIvNHuaPGKukFDgOpp2RVTEcHMqi+8Iw1AK/81
bJw1jhaA3DgI+nCaHjdS4cdjwhdohLhzw/14HZQG0O4kM0tV6DymXxZ7y3jPjAvZ2+jxl9EFwPFY
K38j+rNy83fUZhGWfjNGnh6qFfPbzJ3fEEfI5jdzlYImD8mCABrgVIoS+9Hbtvib4VQQBdcpBptN
THNrc6z356X6wtQi4KzHGGiGa0olWpehT8aTCI3FrESQKHW2tU9Een4E0MEx2/ZVlSzJDbgCgE/z
d/AjQRcgf1db98WelHf8KH3Nb2StQDz3WsXWuP3GIQ//OwoXQkyKiaPJC1teZfTo+I63de+dPc7g
NhNkkb/H9kOTk+aJKPQXMVN6ujUA7LSPPIpPEu7LZ7VOdw2vTI08JcNzDd/1E8BFFWPwhL2uJsvN
hjcZoHHLnjE2fYCgh9nP5sdBbZyziP9j+SkXaO2OvP7T2mHa63dPuF8PTazPSNhXJR3BGGP+Dz10
X5yTIAUHHC8OAEAWkTTrDCoMj+J+fEjuzKunbpzsNqepuae36fcQh9N+hzdhs19sFHSXYxPPCTQL
/aB3oD9s6cONzPAJPIf+OR8pZI/sN0+521DPmd1dv26MJQMfAEp8Uwulg4S1Pm7EfQWpdeAEezMO
GnVtp8tc72OgTPd50th9n+MHHdMW+YqUz3mfrmwsrHg7Gw2DvUO9Y2jWf7jGTqE1aReyBw/WL/zg
dNkn0VzKevpdSVo7VHQg5T5Aaiw+Rwl1/Ez8snYtjKExYeSarcP6qGHK0/nBvyUMTTOpXAAsXCvr
d4d3b5O1F5Qb6Z5US1crl/8crevHI7nKgYKVhsADVQdiGW6Gw33e+SsUDsUUPq0WCWRZJruY3IE+
4F7u+EtlEA6hEY/rp5hAyf8IHDN32gBxrpcYEFJjzl9eQho4p+3kVygvEhdEIIs07CWisFkoWxbv
v12pETp3eURfveSYs7+K9A+FL/3vRjj3VRT+xal+hZL+hBIFt/5X1q2uJRUzjVIX8sHHewscdZPE
9go7fcxPNm1tXyanLKlbVWNNSWY/LPR+LLWGX2LfmOYtEih8GK6mg/2QQESZyCCv1KYRxACwcuyk
KrbG7PfyAy116AS2CUaX/rLhIpXDkpeNgsc2w29tFXacfA/2TpQZJwAdpMDtPb4oqmpHsWJMxnQk
aWw4iHIcI1NEUkmT1OhgnwiiTmkVfs6b7rTviFoJs9Ar5uMK4pTP7da1I9rQRBj6HH9kdM9zE5Qn
ehYetb3AaqObFs076pL8etA0dfWRm3ZNdIKEXxjL4Qc+KQkWMx0rJOeHr8tdDiFAmocMEI+fA6rp
FGwrarCRqCrYi1PqpvjqLn9r41SLh8fIrG6v8htjINB8mR3E8zQ0pV423acMQayQh4JDakQQ+WV8
5G/bm/P6kUKnR5vRj1W4AwQthH7DL0zlcs8FesoD9GIb7U8TpGU/EPN/kMuu0n5r6zCIGjox7VtA
wGLoGD0DHKsAxO0gyUjc3ApRTpDhcjXjt5HtzLbQs7F8XC3thlCzx5Su9IintM/Na4I/QeOnpL6C
a9ipkjvxuTkkBuMV30jJcmghIsx1lyMu2UYiF1gy1jgzR8P1PkGROdTrp2fNBqgFr8GVuZcZdu3H
dxPWU8fGlnakXU9oZz/4HrqaKJhGa2A+TWUZvcCO0Xw67a6GPuXxUZkok820oqo6eC0gKHISdPw4
KDmfWWi0K0YuZVFbRslcRH7I++MWAAvCvWBPwPN86J8AA4IvSfX3GSpRmZhY9uH3BZWemBk+DzjH
iDZgSmXAtsx1SwblSkD3aYuVqsqwAZpoisxAJmQDoCW5fUU5BKUWZf0/EUYj1fj5vuihdWoLzqAX
l1ZVNBfIJ+o2Uem+3hR+5XOUkEOXxH+QPdsNyjRXP98bQmCD5B7IhVpy4UD1w4nh7vWgx1KpmMQS
CIAAAnlIzIh2VQJqzeMn/WF41Xt7G28H3CvcOCCy8GvD15Co3lrJksHjhwBl/U1AMBvTRvQQRKal
qH20EC3blY14yEbcdjlqOgDKcAi/bG+BmCuxokF60yPZvXSVb0gfpiZtC0Z8ctnn2eKHIttcg1BQ
u4Ev9NI0Wy71HYKyXa61FTp2KWDWFdnIugIXReR7Sv+1prcuZ4/T26Fx70JO2N0pYpEeaLNzeIyL
xfIQohm1/gW+1Co04DbzQ07ka8LMX/YYoeK1WOzo7jvJYSO4zjnFNfxNnPZGACanCt844uiBNbRz
oRPWS93WWFXj+pw2YeYXIj6B3qmIJVzhwsE6oqeHsmnTQDDR4yMuqIyxYA716byT1zIc90Kk+EIe
Jy2mgDFXY3uBbkxFZGo4/JB2ckxjoa8XfRNyzgT1hS3JbAm2Ps2hkeWV4NUaBc6FMbgIZEsi2rvW
kzOQw6tI4fHGbS6ICnxq3iGryVDVcQRS19ujWiurBXvqeZmNW0FCyVlEHcI1S6amg2VFlQXicfrw
PB6okLW4MUa9uvbE5g1e3pP8RA5zmox9DysVX4J9+XZ/tDKo2YNyz5KmMcAqRZoN1tE2y0gkyhgq
wsIp9CYfzrElNMliOORbZHX8gAUvrbBNv6W/xAB5WRNdqUDydFn3B3nhaJ8I4q6YGMpyueWYcI8Y
LgMtuNA2CjC48E5PnlN1TgEpgt9V+xfx7ppeBZiYWASdKzmfyTPrXdQcysI3EWX/s3n1ii0aNnSO
Y/Zv2CAQMS8/PTqpQfPdR6j7AQeBImib0e5mz5QTlw/XbijhYROep0UKSDQjSFfsvK3ClhIdpjJa
V++2SmJOkna1iFtnolOf5RGmC2OHdeTT3CaUHdQLqT4DI19LVgdtoP0Pq43cXsdGvnrItMlV63Op
SOMc+rtVKpMZ3OtYruqvyELMyrmsE6cjmKzGb+rwR5iubI6hHioP7FZedsDy8DoD+IZnxdq3hIKI
tDsmdsGJjWDRHngEU38JUHW05wjNK+PffwXIX7KDb4c7wwk1p2w8fxP1xsz54Av++wVcheBt0Fi+
eZwLJhSp3u3WJwYQGK7p0cHz29xMwlASCQXB749+eqeR4lIml4odtbIucLjMO+1deyzjqXM+NDBW
MxnYlLAqFuW30WC0Lp1brdXJs3ubLojhknqDhV4QdFCoZhXS4zSOPA4lOnCNXXpONhydEoZSScjv
1aD04BlrtNgz2L4UClanqeQxwL+beCOqF1E734W2p9D03/EUk6YrKqJcAVutpMCyQzuln5uEUP0B
KrFloVWdG75+yDDobXTWylt5EXnXR33WOg7OOa/tvXawuGsJtCztpHvCXYh+ZwnGUhhh9oOF3rHs
8kdx7g68taDZ3dYosOrmI04twWL/OUTFf+sqpzPXj2vzyEtEbA2cgKMFx7G9SOJHV23nsXcErY9G
A3cPeW4ncxPR95EyL7pw3j5YvFCa/vzr7W9AmaImyymjsgWEWBFbxOxVhuKpTOUE8Uk6kbWcE5Ar
Ri88T+OB0vzR1zT5c9hr9YwA+UACt5LzRUTv6ooP/9gZKgQDai4r0C2+FrguX7XYyS3EejCBT3wn
CHZpVaRtz1y9hO2emU8uhp0cnu51quKENN0TS4QNP8nngU0e1q77thtn/phfMAeQasuLjn19qZ3h
qfE1pySi+OeyugtHvvBq4jM/fLmePmYFSfckmhiHmelocev4n3FYfoF27tKcGd5G/TUEdvle9L1x
i/WyDUO/ZHrhN3m/Me+/xgdztuVlp8kGT3738QvQDs/h+9DBFDWrWQfxXffcSVs4IzfQ2bCOgPLt
0U1RssJGJDOU9TjTl04NF9prTHQ43VUMQkbaMiOgQlBCl63+fa1wvty4g3BnIzQTLdXkJc+6Wr62
gUsngYyY3plYW3tvA8vmhuM6VsNIN22HKycAj6ve0pGBnrFlwznZlTrqKkGDYEhWMrDX3lTyt4/S
wa1qG7h11JXroOktHDFgzGJVORpKDykIgEYH+vxuHQuXCSulTukx0KeEM2DVKh86HcBJMl1wgqpR
u9EjvWZJMdNsix70uNXBmYm+zFRHelY6EBPqJqAvTJwkTjMnHqMeLbCkxwRgVDhp2GXJCkeKh0Ya
dCShJL3AaZGe1H1sRE2gSwtxqbf6xLXorDP1oF/NFeDbsuw/7tRMheTKN25YmUAP5e4/K+2exYuK
nMTHHJDFtNh5/U87aUY669w6nneU4AIkMdvUrGmQlIhHs/V9s/nIn1Ha2V1veHpwbywIYC150spv
GAj/LS4kcQLSelp+oSTRxFN88yDPtYW+O4R+ENhX+fX7335AlK+4m+/JD3+HfhlbVIBgjodqSF4P
eyFdBj2SAAXh64gf78OkTKxWC1/VitWZZuGK3kXy/ISTvvteX7HJan6/3WzrSkPJU6rDvILqPIsU
tElOSe7zj1KcVqtVXArYSvSBGCIVsvt6PfKu8T5v658jv+PEcrOppS96Y/K5OC8rSOxa/6Bd6BQk
GaAIeYDWsRUzI6tQ9nFIMqfAK523nElbapEqGsZJPx0NPSDSAbVRAm7nztc1EcX+CzY2Mg0UA6oR
/ltrqnY4LCYbtxkdLOTHheNosRMQodx/gvTlqcjiO2/LwoUF0A0FUd1T0m0BSX66x29M+aCFuxVD
3m1VJjthVmZpZpXEiKyQHaeXFcgvH+cw/h5VkgGGPWjIFi6SR83MzwzVD4mMPbp0yIOpjYd0aJGu
YkJkNATaBiXKsqJR9CVfY/2Eo/jms0ndSdJDXHa26DMDyOCdvzwwx5bO6u/NKlUI67ehx2Ic0IBc
OYY3i9g3yjdHIgqAGaXCYB16fm2BzIO8zrHrRPWxWz1Lb4ZjWYMXGTJ2UA/Ly0K83/sOf155wLMf
tXwWpjLS+Ms2FNUdhAOv5uH10ZasFDLEL/ZK2WZ8+u+371Oeg31ODN1A15wFJTSCys2Rnpulo0sl
V61qLyIkfasQOi8Lw1QD57HgYD1YqFs3L+ifsJgAQDo7ddSSZqdA9ymtRf7InGZncIS3HAm7AYul
RlQY0Dejqwt/VpDSfF0m35V5RNKDxpJy9jq5l05aI74kUtqw2OtPhyMLwqnz5ofWGkEswZDgOsTd
2CUBp4NFjEzhnGwwaKZ2FOrig6glQpy5PWgzoXeSb8KD8G8b77JGuvxYasUaRrAmzvDaiqTe1lTA
hCRw5/GD/psj7TgUMpQ5MUT7x4F9FzaJAIDsX0pRiskjgVHzK+LPSaUbaDr/S/wDF+iZrc5FD1O0
oQ7v7t4uIqChl2dhoqwY4SVuWSeFU1Rhm4G5vG+QpmVKGORvGAj3WnIDAbSxx/xcQD3smpsruciv
XLdEP6/MIeW+R5KAVkowVeGJ9tJObJPb9P+Wj0DKPKQ5WD1zMrOQTvcQalWQMyP4um19A74MqbXU
tnplXctSYefdsYMUOdsHA8cNO4pH98lPO62Sky93+NiIxFL4U0c5K0vLvI1bJQovuldV3nEB7mi4
9kbnFmhoDEoeGnUg3XoCMyv4cwr9ixFwkgMCDSeQ2U546jJtpE8tauw1agnTlSBQysA8nJA+njJR
1aJ+zWmdCiGjkCKU8yhX6gGPWu8OQ5ALVkE5QaWGUHc+khReGt9ceV399Wg0FOGlmMjWnRBQKUOm
Ag619JdAu+J53LsMdXE8ljDASlpR6AxHWLu5ptK/+mbfVgeeH9RPvjcvhPQDSTakwWeOhZmjHzCH
QDJNBioRwI77Ttj+UbFaFqMtspojN6KY+urjqf7V7JJ8Kg/+zgaHX6nNe2v8I6PU3ulDyBLGXsB+
VSdwPL4diONZMmAX5sTT5nXm7t2Yz5T/7GF52y+zm7PE2bVSUDlBvJHq8J6l3o99tFgqF/A26z5m
/e68BqPclKrK1SA16at7vKDBxMYslNVBdPyAW9xB5O4brupoDztLhPTDDf3XyDVgjv9ONBZlg9Ma
oUYAnCQExai5v+4SF1TVMDJYhMJR5A/bvGFoppEAGswQcOakrG6MzewWiDS/RGUOPgNX89uubvjO
WNhdaYY36Ri/QAd+kp/uhv5UBDNX2yXmw7I1wnoN2z9BmkaEHyWfRlT5hThiyr5MyspoSXz3Y+m4
fd9O6u/RsOIaooXs2CyYGnN0i7kUb3y8Wes7riD5g/7R8qNccMfcD7fYpN8DLxn+ZLitxH2yhgLa
idMb1Z2ZvGbnJxR66ybwVTTKYRzxqWDqaYCgIdwsD6QQSJizE4TbAMDyYw4ioCu3pdJSUXU06C4a
QSbZzis3PsJnszfb+NVTkEUQU/GT3kC2IAV6+gY024UjWB8w2w5B9cD5lt3a6wrSZn/cKIgspizW
t0L9c2ZnIu/KUXC+xOB9FtZoVopQ9Yw5MsdE5uuuQIJaUm6KB/bHBYe8sC/yZNCgv1hy+b9B+l7D
PYlFV8BRWd/gd+x90wygbU0d94wby7AaJA82lAkfFNQHU9cc++YmrjbATtHi6k/CK0pchqjoj7Nf
lmi1/KX511OSnpSJ1kxhVwwJ2131RtZnyhFRpJOrgAWSvewC52JSLD8qEW6eLgxcncIyphekZrCB
8sYvBkicIC65wArBoREvreCKFt6b+SnpM2GQA6R64AJcWNbjUKROZ+jlELvARIot+6oeOH5Jkw2t
0NHyjSbaXyjqJRw5FJtGbh9nDMv/uZXozTnnHGaTgo7jyF4xm+reQE47TS+x1Tt7NmeXcehBDF4v
vEYSLGF3vBQFaqtqqZgCvnrleVRnL/SGuerhLcDN7G9JzDRLmEv+yuhghVtuDQytqUsoCaqfeYe5
mnZ0eOuDMLKUaDd/fZcd3frUO78fAztjGKd1aiCcNLpijFphmGyfDkODIqx75vIdrUbj/D/aNdAT
k/Dla4LTphARQYTVhHSmw9/T4SyYbYhz6nJGIMMTUUtZ4x97nDz9F/SJK7u7whDzmU3U7vud3Y4G
YT4c3qPpgYu3bgfq9l7WKVj4b+snmamc9HA0fNv2wT94OlbHyF7cZ2mlwc+YW0+PCkDe35jZBEyQ
XjJ7hdVC+3NSa30eq6AzorQ5hyNAqysEOxhpFdky9/TUj9peJaIWcBOnaaSQW5RMpWJ4B9057MEN
7fdvQCyDaqvb+3c/N+0nmJpc1hOTQhiq5p4FxjfpMp+tFodU7FNx4ue5E5cRT67wPlrFTi/vdXip
9iCMY5EIwNlMOXdXDzmYTmbYZGMyL+zTDZZH1LQL1oLIrIaKJBUwen/IQZgpfClfl4mE0TtE0xqc
EKG4+QTLelbG6F/zHK7BH549hfqtAG3Av3e/Eht3KL6WKIR6cNhhzUQrqt8AKv1Y6/JxutQT394+
HiEfdR/tlUYDhctFba1a2QCxMgR4jRf0cKmEXkezkyKUBAmL5pcdlkznmb6nthmt6yYwvNze0DpW
6pReAcRXPvWPjrpZWmsYr99ipAq1LfNsB9G9aOF64bqeTc20C6LQGcywIhdmJ/Dj2XtV1fZYzan6
DdGsNFGljOB2p0qvLpvwCYrjvdYwohj9n0ICHpWQjtlwhF7442KjHvg7IOI5N9TABCWEyMK5WIHx
MV7zQaDe6Vu4x7xfQNmFL1Na/p2Ap995eAVlSsRzZRBqWXafm6+zBPFPtRv8fEnqyWyKbs3C8pUJ
aNvZKCBnWggMsogbHLM45eVgy+TiXplMqpRytbv24AU0X1N6Jr4mIvcj4+/pa8vEnZWjtJ/ZkFud
tLXB06/cO84/inJlkdG4fjSMBZVGOkHo+DxrpibbvxsYilVrenQiV/Qg1g590WkkWrWBE3+WU9OX
AMbU7J4ackSsjDIdgwxOIIynAZp+r0uDkn/IKLiovrv9S6UisXVcAABSLTevfDwQDYXsxh8hUdSH
2I2SNLpld1iRfU/AlrE7hncHMtJ2IjKLeb5Q5IynYmhHXGCar6HeJQjb9qwghnP81qvUVjxxKFAJ
pMOxTlH6ZYVnoSXXu5b0tCYwUMaIaLtLVO0ri2fbtK2fKCNkG2AgqLWnFEGX0l/0ZfUhCWCVkNpb
LIDd/E9O4fB1t0soVgWZaNVeaeLU61IGBNJdB5x9YckbyIc1maXFd8Y9STBq9iHH/xFYjeJ91Y60
OrzFAfWqjTq2F2qI0e/egOQY22BzaCysPzV9VsFPJqeEYnfeHAEvXXl/rUf1xuOI9FPR9aphPouq
79lG/e/rwDptrjoGYbV5A+/Q82760Lw+tjHTtgjkS9TLcnAGQVO1WM+AXw+jj/q/giERsRcoTQfD
7Ttmd3220eGzKMd8XEZ4dqiOCUeS9ewFqEe8Za0qXjBkOr4keFU41jVVgitD4fsE9egomFJREfYE
6o/pkBYMrMaA4DoLlZfC/K6gWbkm2YTMKxT53VQznzGEJyymurWGJXLZF2GOyeGUZx1You1JtP5q
wMQ2OBWFixJpwLf9tMRtgTqr3EgfVTzRPZoEYh9tbco1gIO+mpmw+ez03mKS0R6z7uu2eYpK3N60
Z1uttZQAyQQN1FyiDXeJLvn9GO8e7uwrSYlvMPoFQO63bt5vwP2VGgIvlh5CY4Gw6iJJzK/sud04
D9vJRNJ43CVCgGa/VdODggTyayPE+vCIV4Wu2SGDIu8yT3H20AHhr4Mi+Oy3AlIDc4BhrWRZ+Lh4
5YqKk4lv7satE9LF0bLSpXyojp297l+4Ifwl4k2c8k/0sCHxyU8nxJUhYGSPEfGnD7R0nkKlpKeW
5Pw1F2351QcgFUW3BELjn4I1F20W/L5j7lz/tqkPZ7GM0+lwDfMpIF9yz5/cDRAw/GSp3umdqkQ1
09RE+XCzBeFWLjGtJFgY+LYPD1E1feBPey6Rpw/8gxdv73gRD9tqOOHdzVZPd1sNFguUi67MCid6
eJYdRNxx5GDnqBSu/S7GG23eZaXi4HJm9Etve5yMMbcUHPEaLQmvKfU9j0UmmFi2QVdLTj6ldgMw
Cfca0UqcUBSM/Ni2Yt8540sKIlN/9jwE1eYmYHBqzK7Ie0K0bWRzp2aLVKZx9I5DWF/t0a92hMIW
JHzWTlA8d+I95CTO30RT3zw3wyZ9dpVVN2D746T5mkyWskCegEXMV3i/hTZq51Nqhw9fTza5aCIs
16lha6380DZgsOJe4VrZr7C9VqwcytXeS+KkOSKFE5YUJgrrTdu/XZm+YqNLhyhCgLz+1F8IcXAR
cCQPSa3jjt8yq4FQXRx2P0wdho8wMxxY+O4yL38vnUD16crCIVBRCOAYA+owm2U1SQ3KRvtiBmdE
kIkBWvSAI9ZrZUb9w+7z16nYwUJL5OmUkQtoEf1FpagfRJAFAgw9SgdBfqEkuaK8LCaREbj499oH
gnzY8Z54KV5nNgkQCWHZVgNDkMrPUmVI3jCB8L+bxWLUfn/YZaJzfs9+msrDJ9fjmzvRfFp7QYZb
Ohi5GRzydmkbxdk/PEybxUklomiUolAq75wFix9mlMU0xzraIAbv4o/UK1pwofcDsukXV+Jyl8Pi
DBTiBwyU48Z8x/80DbKWl+zS74eteQlccfMefL14AHVIcKFOLYR4HP94H1HAH13tQxHMG78SYcB4
38MM/DdzjghbOE91jrPiivYH5Lyvl2GY0OQxKoWAHKjJ8caiRMmJsQEfAPqQC5pY7a5wvosq+q3s
VWadUYxx0+I674QdS4ealEmCLRlPUfP1RGrGEBQkV582BGQH+aieGqZ370rQzSZTDtsU7MugD7PY
CvpenUkZ0UNYb8sVBKB5HljlD8MNCpJeMrfmobAd8AU2IjfAuPTnDjqjt4NoYHrD0r4bI/KAjOIo
5aI2tkL7mEwKqoK0Oo/zVjHLH5gmA8ZQNXkI2c8RcrCh7cTwDUm2hrt+3OsFe3gBOduO6idW0lJm
CEDQjMTy4osI9sSikYHhYbY/lj1MNzuN5dKazd6L1VMR9n9mSgS2iwW2g4dil6onD0Mv7W8r1Gk1
I2Ub9vzZOzpkzCf0JArEixUfhSlQGoJm89U9p8CyJVcWYD0CQVswGCpdH2jY2lsQv+4b09jP14aF
SvQMgDXJrPt1k8xXsfrVASPdjKKYhUUcD5nTEUpfeVP2DGuo/dahLk2znwZURs9d1E8c0bseDtG+
wFlHjUavHJgREMZGaEHkMqBZ4RmSU3mSR/rLwwQJIUDGrpryEj+bp1VG9BGjlfPuK9tSSu6AVUDV
H/KlZAhtt6u51HIHy2Kc7DNgzFRUiIYOh9kUul//U4+CN/AWPuobh8qCHJucXjFHqSOXfJNgcMKn
ZbOQKGvFvrykQ/9o6HoY6ChEmAa93mCfIPyiMzDE+nADjnhthDpGL82bdAo8Meyx1GbmWH09dm8t
ZfcIhq5n9hkSkArpz1d/NYxRtSmh69qteMR78nuARQm6mSzaq4tO8uzt3dcHhPK0mDQ1HM6KPwZw
JMrbYN4hnQhZAQ7Rrc7RU+w+D7ZVlne+SNJx/xR0qzJwIF60RDPirjTuIAwsEqe6Y5VZztoxaR6G
MtfAEhykcgZHxZ7YQ9/xsozy/xrcdXL7HY+N64r/P775n3E/G3iEg9Pz2XXIiF5gxWWvA088daUl
VtHxLfWQOhupBa79PYNFsMv0P8ScKIizOxdz78AGbraY/d0238hnYQa0tXj3wegMa+y7tgmYeRVU
glkfFUtlcJ0gPcGHtxUO6Nc1PaHcN8NQBCqbpN+xw1AEn/j2PII8QGG0FWYQDuRFqe+k03vqgdBF
xQO7zEJi/FNFXW8gqxUmYIEQ+WgW0IFX6gpq/Vfr5wnHqjp5yJZ66G+HjoOsow21i5wOxdfAST0n
Sq2mNacJbQ9QJYltqCsaSALGpkx17zIZhXBKhr6OCnf5XOyHNNbP3qRz3nSxOB2894DBZeV0HCyV
lF/BbIkdDqM5j4Xd7+YPynFWf28gg/PnHyaLhzFq5X7bPviuiilt2mwL9WP91/Vjzyyvquc+Tc54
WcqbZ9vsRTchYF9JoY0HH/0dg3Hl7b1e83lJhk/vUhnKO/8uEhj8bfaJx42/5cbWbKgoshZBCQJk
RgZ5S+4niluWijymDvH0LQrR/MTYokFOuw+ImM3pcHjBW7SYTc2sybB3mgnMmY/Ij61cdFYtFd1h
WdGA3MpCvX+PetOr6YYREv2C7ECgmlR68ixKrS6LIFyRBpXJGMxrLaDduPDl7JyHLP0zzUfY90LP
mBWAyZi08Zl5HnuUpdAmRQvy3O4QYhk2D+8BdY0JKplkoF97CQFo8wy6PCGGde5sWMvkeTvL01sw
vQpmv//mfIznZhyFbDLADneo++9RyJP25zP1HF+AuK4YtaS6EzCUY9RqC9y1BQ8WBq7G9wlL9Die
ep1CoSCUpGamWVz6ZHmSoxmIP8O/soZCOmlzOSyK0/ZM2l9lYdzuahCPpbx7ZQjGqM/SboI8z7Cj
znhL+q6k6pgIWUMNX4riHOCuAtAL1cofMB2n18e9Ap9D4yNPmXwQReX1MkoA8C2Iz0XedGe8RvZM
5+YKD97JHUnEmRB/cc5n88/SEzPnVwHygWQKtbz3to1zOM6sicH/JtuxHun0BpKDr/LGtSn/8q3+
PbsBVhNqkTvOO6Sgj2Zm4B+/VylHIY1FNkswkKkdbaK+ITAkW9ZFGsVjj1FQBZSB9shD1csMxPaw
d97BshbRraWWV8VRqzpl0w1NbiZZBy3y8PL7qGPwnorETf5sBdLLTtVr7JcVrwmB1m9ctIikI27u
TpPc4X22PUnliyIw9bB3LNQPUJqhgO0IFPY34JpUerBUSJK8DsXXR9Wk083pcyLhE3qVRciJ9HL1
BjgO5Ii18P9ICZe03YWaTCP0LIz6EBRG8SHfGTY7v7EXYJRfpm+1Jkv9ybUp1ZG0z65nXTNyBP2O
xB2qVJfFUISswjZXWf9VXi/+CC4oXRzSnxE8d+HNuQRbECD4zBA6OgH56j924T6KDjrT9J2dLBrx
B3mtwwNzMh31b00+B0MB20+MOGPXv6SvhLOfpEgcMJDcnMkJ30LkGu43r11hZylu5WzygGyCRV2O
Sgc4alYU+YU0ZmdLwQ7nmyRKFoOfSTN/gzqnjY8FTLEjV7+4xeh97H9x2gYDddu3eJqwfHaemP8D
FRYckm0ZU/HWRGq6n2pwBrTVdKxrXm8d+uRf35iGYZXXrhCxwyH/d6d0Rs/mAHk3L0WOFyzlSadB
/rvGu1GNZdE2EP+X18DZ5RWBFIU/XDD3n+fSRgBHBNxSHBlIW8a5yyfPrm/s4nbIEc6yTgys6432
pOO/rMeq+o91NlP4WDpbEZBNxPJ8otYwFzLhfOqLYBUhEmR1UTwV6cgLNiqbyOr1y2IkccdorNTq
EihaEkta7VD87sQ4KNxj6Bs0LSg284v72rOCYHZWpfsKb+LSONPE89d5dA+9whSot0ILz9bFiRQf
vAu5gLaaS4mdn0LhwH8c2P4vpQ/E6+8scvKjwi6hXebMGW2OEs3DhEWK8bE2FwZJVqM6RsF6lcdz
DGS7+pg2VkSLWZ5br/rSfU7jk4rL/3hNH3fK/z40j7rS3JVM62q2PO1sqj4Og+Lx/Zuq+dON/bLw
bvq24K+8lkoJHYHmkYEVvLquyTVX1rlO7TDxr4XrU9w/g8ZHBe5FhMavBCFDszDLxYTWIsi3dZgd
pcMwuOZYWtWpP2wruFZ1sqjzqOeZTTcPyy/W60kGJ1Q6QnxKzUjDnOAY4p+SOs4/Uht47irmJbTv
tkX73PfhoyBRWVdoJjN2+cJ/FkHvaYMtopxlfadHgLxemuBMggh/4c5IkURFhXdgsP7nrjmdi9Xd
9RvmMdE9hndnGJOKKRYObseesRer35diJ52TDx8YFy9aAKVCuuYXRtZXSv3S8gEWZSn/TYI9ZV//
yhY4WJAH3yTeVydbNvHuRXnALsgqzhj4XjCuDpyJerXReHQ/tc09U5Z1CnaSKAp2q81UKuBqIfJW
CQIUxAzr17o6Pu7Yyx8cQdVSL747Du/3NaoqqAUZEO8ouqDfPBPt+XB8KfOHSLKNCV5DaSfKWSX3
YPw4NvCfodhEw7VZnmk29fRikxDH76i8lKsFJI1oMYd7IZcm1rWVI4OjLmC1VwyqxusDKSOJ8aoH
9wvzb5gXjtUxkvy6kabNAlo5zak+cxY0ye/LOgUdOJaTQsHHlacVl4vukKujDJo8YS1j4duReNHk
Ldu2drStxxCy9TXeYAupxPaxJW8GNOvOhlOynomkVvLJ3vO3XrHpwRPs8DdZNqYHhWESb3fhGRpp
IgZu1glGTqrTJQsGN3s3I3lv4R4XY3q49MdlDXffaYXHdhhAs/d3AkDjLnPXvj1JXfOKOT4+w/vg
dZBKwefM6gUVA1GurOrA3CH3VwGA8LYiwjaADnzzLLd5IMSXi0hcj7tqyyfASs5tSUZaIYcHm+f+
y/pifWmCEK8fFui1IiVgoGnjB/B7pcyTJ4A5KMkAWsJaxegL6hk4g4Y5LtZAPQgVlCyBih7tY6W/
L7Bg+p+w4wMZQqs116mSeOCm3fSTXmx17PhSfReeD2KTmz7ijfA3+1uSnby6X4Nz3vnFWxvDQ5tv
RcCbkwq2+1EihjFTNH6AC55gqlOBi/esajSreimhStOq1dPbVOepBdmWzx+mmbWcRhrnoaB+R3zu
ooZmCXqqJXh7Mg+TzPdqAWOaPRetbGqlWwLwpmaLeh/mWTEqWNIocA55ZVPgtIsxiyo8baVVRatb
KhChzr9jMsD4Lkf8PWyMA/T11z4bqr2kZY3SvDSSvZ3QkcVF//Olyu2SJ+ExGMDsDMOeHMeqQzho
QmwJdYfZMu9VaQRW0zlUxJ6J5CY/llTno3Q1ymNmb9obtRHLafekBJd4PsmxHrlGYXMQ8hzHASNm
rQMDdV8Cn73rfpitIwdzgbPhFsx5pI6JTyWKGqOecMiupVfBIGp2L8xVXhbXQgyXFBNKGpteNp40
ntLaxrdhW01uCuw2L0oUmFYPBo5evD6Tlod/SgUHPkBSoS+rsipp4zKh5f/np7gMcTuwFzotzhtH
gpZYfXZ08StCsyV5mou/ojiH4m/pmB4r2Vp43MYFEUX5t2SsWMzWoppxHRu60AsOhE8paoKIBJBT
6MJtTjZ0IG8jALwqfngJHYIMKMxcc8MA9iRlAxEyIAJVu1sjdlsbvTlfsfseUyhN8OyWxw7pvlUr
pJ9ddwVJ+s6CDSZbQX3x8yn0MfMe43/QrBnTiwXPZGNgK76C1FmhJOeHlN/QlJzX8BOMnGIIPteG
wpKv60PO46eiQSssXHWxdJwALovS8YXaSpZ8zyJuFTp3tiwARc8RJ+m6+Z4v3TaYTKMoxOKjre68
CwvBcWsPhakNreuUcOtHwWcQxm/7HVH8kqGK/50dVADqrDS8JdzaVnof3/315tUWsTjLJZUhYvP+
Upcm6CmgWr1z4Xa99CW1R7Sg33kCV0JEj3lJtogusVPwe14TGu+dDhHwr+pTLTkvRK0kSAx+fEa9
h95wXOiWnp6Rr3QMR9lGZ9yNLYyZnajyduMNBVzGselkrpMqxNd5Z/elKwEXxzGEQdMsPciBbBqf
JinArkXtfcZqeo6sz6plbQqamF45GVPTaYdPFA9oStm2MK13eQ2SimE3L6lDZzZyUmBle8HObs+n
MJ9jO4BoEsuSNPYVrXAHJ6BbIL534FzKCOvXbE6dV8G/qVCXAobXa9QG1JkGSLO7pbffSuQBWMr3
8H8FdCTNlMgBVUgjhyK56r3s9MD0/3zetGS6csdnrycfp1dK5Qa0+rysVayjWt/wuv/CC0wMHpPw
ZT7ip2aEU1sOP0HzARmqqnh8RZZYHnfeWAx7gguaNXoGjzARrFs60WfaY7G7e2X5qc7+7C06n842
YMVpED0ayTQpafb95I6HTZ6YEqnL1XO9WLgps+oH4dPSAIiRhSsaT9Nt2QDe8EwneaYqQCbP4n9U
4l+4eNIDZpIEqm+5yiOm23LDZaJ5WuerkncOh3PQ/rkDiE2//cccpXAjgr861v7QaAwHD88DJX5i
zXvHq27P1Qy0cyT4hEzPN2pAsaZca+bFWT62p1LQIbJhC62yYvje6e6LGqQ++uMwHlWFP5knAx+m
Q6ovoSseuhs40hmxS2D6E0nUqqGv+Xv/ZtWfp0zeYx0qOKwCkqy3YMRF9rvsoiaxPHHVJtO5Ra7L
JLWnNj67k//mHuL+SLkFEAFkGMxitMSZVrDd4azc9UzRO8Q9mUb1qCj4J3nzLOKUWaEIA3LIY1ce
mpHnnYIXd+mZZXoMDyajyA3PIJWydZLV6VGecRruzte+KHtB3o3qcODBqudf12BwDDGM6/nBbn5P
+piA+3oV95Osa+6q3litODVBRwIbyF+z1O5Q7xxMUm+GHcY18qnjf60vu00ijuS2tfqmGUDwahbV
RcndU0ha1G18HA1FVEuAntBD5f5S9jnrlIur25OUM1MYiDFNWBggxhrpJf5wctdjSgs1TzTNj/VS
s5qXEKKz/qi1vGXzBXhJCqlRgp/Z6bmK0q1p46G6uDXHnO96mRFnMrz/UkkGzEyVZkoNIJuI32AK
g8WWPxv6PfgOi04bVvR4X8vjqUxk3LwdX1+O2CAuvUwsxyJnkVEzbYpL5Rb7cpa2jAJtwenNBOKe
13Yev02jjIL284a3f1E+N9kP0DkoTbLNEFBTTN8l+61gTIvrBIoVRoNzqpZjZuhrgK1sBSmwe8Io
ruO6Jq/O9zydVSrCGyyhd+oujaXk0qHC8Gm/SQ7U92cs1W2vlaam5xZxJb5c6/9dnXurTt9cxViv
ImZwW6fAgts3ehs9SFYdkx0zCSLbTfv83kBcOe7pdoxpGpcyZnDKcD07bbXaMDOp/EJtAqnwP6Rn
+18Vf9jIY/TIGFklKL8978VDClQ0ss5IDzdeVgsdlO6AoB7uAnVe6HRoEh5SGtjguuE2DyIkLLLw
5Ap9fLm/Ty6E2MoJi2bK0N7MIVxDet+mjC4BsobvfA4/doFiREiRTG0cA351nq6kwH5zgOaw3t9B
jOQXgu9vylIqXyp95jxyoi3FIzJ7gDvNM6X8ULMk84UETmf9F7LQsDNTMRmkgD3QA+DXu1IxR6CI
LAIJDMOPWuvjhPA/xl/gtlPXls1j3HSLPxs4iMdHEqJY6VSPc71CwPHfHEzTYkXRFYKhjpvXLZmw
iMsRV+aZWH2nuMnxLelxTPdA3rq4wfIpwCag3uJKPyYujzWvl+rtHywNIx9rdrtLvXnX1FuJROqz
tH8fnNmY/7P9o0bbAk9/BKuLJudFsR73F3X6LqpXkgnXeL8hpvWG5rUh1n7YQ8n06NaklcZ+g8Ad
KRKQv69Bk8phk3iIOLvidU+ka9crak1TcLdAPSFX+4ZbZ6W+De8j0wH1obnfblI8AAFSqUMnyBGu
tWvAmBXszu0iqZzmk2+mzHBa9LreEJCAqTy6EBmSocBC9T6B01yA0WH8WxVOtJ2udP9DEzCfYrNw
4JFIK8P5Yz47Gt4H7A/n/P+8nrGBurmMXei8e2b0n9qUCCTDaOp8anN7j8gYm4bMAVcx7/THvmLp
oxBCvUO+3apR8ZyFycgMv1AuuoS2IsYANVQbpyyImfSAyKuK9a9zS9cIfQU5in0o2EtToqqvt/MH
jbSSzVjRDX0pefaMKZ6DgIgcIqox7XnTQznUCEkuenmKGajc/XBqrKsAai+uMHNRxpPSmx633RUO
ZleQV92xA1SV1R8l+gWU88nVqpAXKrNOC5QjLjNMIQ+lBgrPxjmFopZdtEgplXX5XTrWXtQ8RUr2
JDMT2moY0ggIaYdkMrkPh5hcdrjr5pVOGqGTFriSD3jg/Su7llVErDgWS74A9sIvbokI3V7lFZOi
vw8WmUKRAel0axGMVLSSO+XuakOwq+mYXJ28zcR62ybgRRYqo1SaWZPJx224ih0W6/O51vJI3+At
TZLBxOoNEW6iAEfkAiwF6M1aO44wWWDIukxM5MpIEHSrc3xBwuwUGBRCvg7JrHIk6a0g10pwcK1S
UYy3W4ByMgsPzB5Y8LS5SkeIl2qrkBlC2loU0Di0+neKnVI0eCnMcnVoNFpruU1Z1DrBNqiHPnH0
mxYlQPvnU0197xZnz0vSUkGW2pGLkmsY8o6hWb7nVCJ1iqYopdyIkkVcoy0FXsE0oVHFSJ9T9Q17
cLJnlXws1brHb+J/GIxn1AcdxbencEi46Y+GRAJpr5gAW+x1q5qrknAUIVh5TGeCl2v2MlKc1vIp
B38d2q8HPfVV5ZD9UuyG1TGolErWIk/TDHfTjO8qZmGD2Vc2ouYDTDidb2nzdy+9GVde43cDfMBK
X0dfvDoVuz18TpVfo8lLhUYwno09uZ5aTDEnJSildf4TYHmRXS9CVtixlCRXEvC0bwMnAN4Z5Tbd
zzOUce9GEm3e8CAlzNWHYv4L7dCj8Vqz+SjdYXR4vCL2Rg2jvNGiauYgAcW/X3l+5b6VbdSBwZIz
res4S0FnzKsqnAAZUMvl9aVWP2k8LDkSzeBakjXQKnRoAHfofsJdPdjm48dnYPq4cXXE3uI+ZRad
UMupDWNX0t4ux7BY1ydgdUCPXfRnXjom3sNkNiJJlKJqWGP112p0wo2BfSa5T5JOul8q4abYKXZW
eD26A4FoSA7eiCciN03uzSQE4Fm/bpb3+DsFMlKVjQx9rDsXKfZXB1UcrDkfNTDgaNdnAOPu1BAm
GPjgEACukpPgtJFgUk4kAziQsJOfNgPZvQ4ONnsKgpnpzZF0yE8oLEQNeCn8z+Hox8EaVBddFzu+
LVzFs3SHfCk06KpsLZMrcvnBNwkKku7uwTc+Kw2oA0tGels+QS9u5/uMdFMwSEX7JshWbLQH8tyz
846e2+Xj/Gq0rbWVZOE4p9cI2/oUFzytWQxGDkauG5X1mE6+8ZQ8JffSzPWTHiVPawpTi0h5KAGO
ZecsRMFiAb1xAdeoubPJyUVYAHPuau8VyNzxvdFU0C4nWokjh9zwhhABCX/Flt+Z5aHve+e84bhZ
+WdPdHYYftdwP1ucU7TjWGHlIgujJas+LgF7/jBfufQnbmcBww0rwIVuUMboUby/33WZZZDMn/DM
Z2dFRAdToxXIBoDuZ69Xvab8BCcAYxy2yO1TxTSXZD4kEDA+8Yj8mOGGEMfmRFI4wEZ9bLBogPBK
jBKDRceQ/Po6KnpUVrUVxtt3CiPdKgkNqP/OPF7YKoMD6/7TUI76BrdDJhnWNRYqyQ2YGzcaiBZS
ydMR/+wNvZVLfz6plY20FFZcT59mkKZClpBsNRdO3FZjlLHQy/Ywh9yiua1cbSeO7rPsXwQh/vFg
aac9IrE+S30pcDEjmI3Ge+S7ijoiIfVtrtBOs9ZL54HZ5yvi7AVjfV50bKYLPaymDIGJCyJp9cnH
g2d6rG3Hoo0gU49N/YOXDEhLHp7Kdi++MN3BL4NL0w2eiAt8IprL805wLSYTy0TNwydZrjSdrEND
Ia0oLl1yxmEQx7v3mzuonV7LdVXr8BSmnzWEI5b1I0wm9x+VMqRxvWkuhpWsLOiEBl1g0RuixX5M
U10dSinZR1iQ36v9gvf0+inHUU9Ka/b5s+6iSSHJOgyyIm1w3CuZBDFWdY6DvXgSRQTNn8LrIPcw
RX55i7yBXDGpxz7aFysXbwNTy6o6QWHd1oq2Lt6pLZ+O+Bj2fs8arNiABWhUHLsrKRdgJuPgYtU0
I1bGg2wYDVkdCcUzmKT7lJtaYwhNaXJLEfgD2w+6CZ8impD1YUXerNNo8czVWwfivBBXL98iSlTQ
Nko2firP/7xM2ikzGFDvIinru6V49DZUUMSDG18OWboCEdmajrW4X0F2E2AucRu5rQeiDoI1ZEGM
/1pvnUNHmbXOVDcilpaSxSZXBLpr+1kAHeH7BCVNDDvYq6Ei0ksYu60c5YT/IAeRCHtruIjR1h7K
r3QXBRG+xB54pQ3QfAn+m4Lmj5AnfVqd0nUtTDN2RRjlGTGv0QxNYmK973TUA9ky9/YSK/zRoeDz
qg9hWtX5nTRDhV/1LbgdcLFb2GhQy1h4qrzCKaaA0YTcAAAOPfa4JjATmQ7ZD1R+MvpVVUEBwKHB
SwfJ8WNeYG0jVeT6MZzaiXZqWzH1EovFN2E6MwGWKfUbbExiBvEkzHUs9iPcstSdct1GDqbut3+Y
p9gZgkIytE279rrClulkisOe3EiLYJ/7QCCuYqB/6SJf5joso4swn3hoI6ThJwCczLPUa4MtKWdN
k536l0Qxgn36mqXk+wLuSpZkCAMd3+/4C0KfgYaXdoHxayUck3Lr3ca64Yj0t0DW9mcTVe1jI1SV
cW0OxIPSG1z441F9u5BbmUYsOAyXFRBCjJPtjTjIbY0G3DkLWoZGqRgsmy6jOsTY34NrBd93mwDP
8exL1iMeZYui7XBqZ0hzhWEUFXOsLJZeJcVgNCoDNbCeb5yNQzRVuFW4aGpWMo6wqzcpr8xRq9zP
EvnbUTYSSjH/POgebRuJTLHunztrgqpnMtehcu2sy24SOoTOPmXFJn3S0tVUnCaR0emuPR3Qus51
qsqAyH0C6iSFJ/q+/67sEDaQ6scBqnqPZQMcqOZkAkOLiUPxf+DfN0zMB3d8NTrGw0ICl2o+8Ap+
mBybVXnkrx8UPttisx1d2bvq0cjtL7uiS0TkNQToFuIEgPDesQEYvvFr2PNOoA0dQ6l+ZYDkk4/U
TU8k9sojyy5pHGiBSxGrUI5GPuRcoPPTXw7s9C+Bz1+Zh49gPeqZGlTTz+eW0BhB28q/qZ0txVBN
0INR9sTvY6xnWO8gf+W3tDlLr2OHqrGBLhE8YpUsc2wRNhPPOR0iCPfRejrer25XmwrLsbJcFu3k
/M1AHiyOdrqnWP2W8fgVGKa/4BS7ZxYKQ5dmpB1N0KEgz19vTzCmhxY4S8aKlyv1hZ4T1gHcyGBw
3SUTjw2ZfrpY5LSNPKyROq4U2iPXgl0sPqdN2fpua8s3j2cuUDrpddtSLQQ89w4n7Kkl7w0rgY9J
o/I8Ww19BAWZTunHTe8ZcionfWWU6EQ6Ym+I+HBVaqCPklc6mtx80foO/bO2hxTtNQjEXSQL6XoA
qmF+DFj+GlHqnWEoxjskQogFGJq1c0sGcsachOQDHhrS0056K4hwFTOIalfrfrK70vYnJ7jNYlz3
tgyLt0t4caUnsBdRTkIshiWiTHDpYpJtZqcGSUjdrwkDQ6sv8ymq00bxmEPyDCXQULoBP0LiAmfp
laJZoE40WL4huPh1SlRMa1WVZs02fUiA1Hub/g0xKNl1cDYib2jPzm5auyd23jYJFYk6LBQHpmqp
8lvYhG8JZdbN0cFZKHHkOXATfJgoLAY1JORtTm1UbEsyhOHI1naLv7LP5CBO8Ju37vLj1COZxtSF
Ew7HCBee5l/idNe92g7HLe/XbtgF5pVVEHmR0O/Ab2YX2RgCRl2ik9gPC4r7KqzP+L/L81zaB8Cg
qVMYrsbF10cy8JIRwYmsOs9iJIYthd4Yzv87FlAV2wtnrGt5E7dJZOAxbPR7jIzKaKCtU7OnuWJX
aSYLHspP9SElY2+ivsDLaYjkL0Vkl/sljX9OkLCCGTvY2nOta6D4qZfIk3oWmeFxlx1VMT/UYYPw
8RNf9JqkIk+2422TF8vwdBlhFikoUwfIB6A8lv9lhxMNaS7V3pQP3q6PTe/XCwOZ9zCRhq0oYUP4
lmjwnXfYBQ1fH00GBxLQuvYytMctmDsJlTOG0ZqgCwW+RT/shwZkjBG+msQOjycicUo+vFRo0zSG
W73LzMoqM8Yufrr8pPzGPfE90gOVJniqpMPgY65QQkulYxT36td8VV9jU9ekqKiEFzXWJvw3ul/B
dP7pozn6WyZoWKuL/hrXDpwg6VHQd/R6Cp+XQBEc6lWyM3p+gdPqo8Bsam5AFgTA0cI9RTpGUOZ2
+l/VNG5dyLzQ7OHOpkQeu93SUfqCUML1qtChKK7c6TAblsGPoadd3vOidRtCdsWoKagMIEAFMGZ4
fb+bR8RKJSI7JU+GvuJWFFPVi5KygW6ZeAYYR2X0V/I9j+6rFnbd8mlz5YINt+gsDUqF0YGutS55
gq/WErxYVTI2e2A8KR1a6qzXmH7oL4tAINfclmahyjxAXsB1DfWlgFsvdQnaL3LsNLx2Vd7zihoo
L/lATM/hiYVKCplR/ulHFFf9Yt7aSNbGI1ztO2X3uylCYHScQgZC9rzXNlko2bzGC9PUOBigwU5D
PDuQUEpLomNSacsP88CLrg9Hl350KZmmUmkTD472f+C4Ej3R349aDAdXgIrn8dW3q3V79K4/3L5O
GYKno5Cu6NTvRZyngXG2lTAAbsFgvXnWQnMc4PErjDzZXmWk9NoPZNU2Rs2OXneHjP3YLpGdp6Gr
UER8YQbvikWRXpA+Jgdg9mDghEHjU2fgtIE7Mim0tpSsgS81vtUl1a071H7lerx0hhQAassg7LMT
lMxEPGyQsM8T5sYErW4nw6TkAzwwtMTlYhcPt4Ton29D+3oQmD6wGUaGaVvMeKXcgwi2W7MwQsU0
ktm8Lo9ATZdPWgG3vxf14cFVu/gXYh4ykCfBoNKvxPZRLxBeRmmt4lwC3t57m2jI5ubg838v67tv
EyinhsK+w65oJUenBFv3RYiArlztqoN/Dtgk1uDn1q5JUTpLumse3E91nbZW5PKpPVydtg7XKHOA
MNOO+fwMIJuu4phiGoZN+3kQb3flK2ary8JfeqWpcFwZ2zbEWhSWZSUqQBvlaHXHElKRcAQ35sgu
WiC+aNKy8zxZw3x2SfgArP80wMzHBhHuuitkOwz4BwfR1asu0KVbt/SC8biYO6auU4Inn0p/o0lf
K0UjeddOjuPA774SUlDx6TLdBoTTwWONnCTU+iU4pJkBBUmpFAr3HOC/wkSYBhC9BxzdRLvbpnZc
V4zVwQDgp9nkIaRRk6+CPwR1ox0cy07om/ilXyjHQHjG2jsqYi25pLn/le7FRRPdZIX/6Qdok3dZ
jV7SCqySAZsFTjTnxLz8J2WZJxP663Cbr6YS/0Ih/i/jJOMldwi87/Jgzv4CKNdQUODzsMuaIMFR
BgVZQyWNa4nc3RaxO7t2yBXhOmSVxdPk7IdIvij69PsqE9krt4OHAryI08SCvxi3ggX6Le5leCya
e/8yfCYQ8YjtKHkDzHFyPPBvKalnNK/ezlFGjng2Nk/ZnGYyFYR89at/d3txf81OZIZe9eh96s9m
iczcm8C0bYzIbrBXeMjO57XmHp+pUydUftDKF8TPibj+qkwgootabOHrIFwyCitpfq6E4KLDT0y/
jld6YxASBUS/gt0Hn/2Qrq5glgKu58CBmDxyCz4LD9nDCxziqua9p6pPbtLcHAISMqyMrUsTldz7
/ymk2Pk1LRRRnJTDZchfDC/N6n5F7eWJCZ9qD6qgak3XygzlNstMEu1dB2FPDXXrNwe0DzSTKjCM
/9OgORODBZO0uL8g1W/e1ezV9Rfs6cvdaGyh5MDDzxyX4IaQEmpjx14lVEkjZBBExTe9Hn20B/pj
awJw0FELhr2QkOSBa/ulY64jrTXemo8Y2TS5rxDVAvtb/GfDmRl9c5ssgjrJqEUXLPSZjzMyQiF7
NhUHLCcod5FwS4UfbIe1M6/fPWailYP8jdDN2b51P24Xj3jm/gq11VpBWa2rH45eM5CDx/8l3JxR
HrFdiVEeuQSZrKa0Oi3bqihiAeUhmk3O1t1m2rNSBIKp3fCxRyOG2y5Pr9FRG0Pr2caJeIMplUpM
2LtI0rkM/K4BsX6/8MnBpMarWwez9WRuMPRgoqT7EX3LH/C0K0uHbXNooaLoaMfJiQ1nSuJLFG7j
bxCm6OVX6N5N5rJs1ER2G0k6Nlno5ETUGljQF44Q2lNiJmw8l1kp2MtgDV668Z6qXH8nUDqcfl8G
ALFV/sJ8CusAgDyghr8ORwLUFtdzM17nVjjGmzdFmroXEbHNX0bnYrdZKeYynOdGJMB3WSSGiuBy
upLkbNQy+ZRxwzZRvgtE2v5ORumNENNJwuhgHTSjkn6ccr1GAtO6d+/U2dn7aMjAb/y1+ycZkkOO
hcSA+eJeQJOuYQTMatLieKC68snyyUqv0lfFA350t+NWrcY0N++n0lkbRGo3HAkJSEEUSF5DJWhS
xbwHWJhcwqlIZJ1LpeYizp9JE+l/3KlGZiT7ZOeq7Azi74MEJ//MzOuObR0OtmLer8rJHnWNWBct
o0monBzeLW2zEtvqiLuDJ27PkHDMUMtRIpECaE4RY8IjyS9EceJwXbC1Pc1WD0JGSEa37ngKEatN
9qVBGdezJqgQFx6wVYFmqzCnQhXmlZ+1Zlc47gU2rD0ycZg2UUAE7nAalQpFUzHfsYN9is0VUTQY
zY+7MS5R6qtk0yOdx144LBsYk/fS47MyQmr5G/0ULDdW2VH0Da0kiXs/0jy0DJoj/poA3kI2bZbW
qbkf12yAClZ+wp3N2hXKuATkhew5XInIxzkcZlCMsx1dpt0DLqf3hcEGEHkeaaLhn/OvgOWZ6ocv
YXaLUyNBkgrm0LRI2v+bT8LERu8xxtYoOIW2rQ3UsbLt1xBaLsCIO2UboV53qhT64tprUTzmf2ME
1O5V9oK9kCM8lALD64/KrrwBX2Z3pAlOTZHhFvOgrhDxmsg1eYniyN1reSKpbAiS86uc/cA9sdOx
evQxj/tlvYjcEWdFGMqIQH4rwcqz7XV6qpOW9YV+r7eCEOcxUHOwtLJCUExhpQRyKK5ESJhDMdn0
DNVj9+qZcY9fdstAc4RKjV6RL9FMKXlNyVlVgYdTaSu9+oucS8Dv8/ZXmsaUPCmBETGUm92bCAnk
TnhpHKD3/WXudklD9cp9iuzMOUrGExCfhY+n7un2ymaJbYwEL0WYl3zhpV+IotC3EGg7F8gXMTPG
J+xC+yepQR3AL4/f4CWITwie/eVCBUbdA+/wZZ2NelL/RzRHbg58zDFJt8Tm9JRAlqpfffBhnpoJ
FCsNK4Vs4yWubuX2LLxBfUpm3O2Q2jSvxeptBrjpQ9s41w7ZD6xapV2d301+QMEgczd7T3KNbtw7
0KxedFY+6iKmvUyQOXICv9v4Gxy9qaAq11gb/IrXrrEgLlEv3utnXr2JAqaflc/u/mDUd7K7aBcM
pWm01pKvMAaLAQnhX7qUcIojX+6wHajDDT/Z0b9ptnGU8uamoNwkWC0JHV/l9sLHq0yfScYqtg0t
dqVV5ak3Dp72c7DuyHulMgJRRup8ieltgZX6zg1xgIB1Hkj4gQgLA06lR7qv3jdYqU+xrSwq4t4n
7YwKCVOebhL/JdeyhM1MI66u8nVcbkyiwk7fcYjaXzcTf+bfWxJxAATvNG3LpveMcWa3uutyIqnG
+TQGHrXIOxZvV5RpsZzkXOx0fYGP44c75dVobW4J70YOHQhg9/EtRTCBGFcQpsJZNHMps96db3s/
tDNjYDd4N/WALNXb67GEGJDk9UuW9AsqAlOfyDK0IVWaL44tZPPD5+dg3QqWmtthtjWoORqWNLpl
arqdVqSZS8TRY/NIDap4oLZgKua2mtPWt4aQBjazi75BHAih0rlrzmKx4VGO0SLtE3g05SYEiqmG
CJkWCQ02eAJAGJ9T08xF5mEAY4EEFZyMIFK5iPDMmQ2ENx+XqDhvn/Lhh1Z7Ij1TPDJNw9Pk/siv
uy+ezTFvbiksVzDu7ICDkQnlXzdjxNlHIx1CeaZZ6lcmnY90fZuCQ/1UM79W+4rxRntDxhpicj9P
cSjv8hTXO5KHHqEkGIeCbddKjsLQrbeGJL7bvzUT5ynQhVChHNDBFacU9nRffratOSMcva2/Z7DX
5pSoBs4ANF2DhLO05IN1vlOHArQmwLr8cHn+gMuxJrpxYZHhJCHgWcsCguLUnWyT1pGrWH6Nr8Bc
pr3OLaJUL/KHmOeYT+WQWnq4/BlxvTsk72wkLVAZzYAm+ywR4jhSx7WLXEbAJl2h+izjGEoRMGO3
sK5j1n1pMFj1//H7icEIy8MDiuAvR0OD3GDwFpp/cpoJcodDwTq0y8w3eoVvu2YMQfBSWGsCmcrW
YfRurp1hS1H4ex6uS+AWbKOmoVppCuVtevGc/hedUjOGN0yX+XC9/4WUWmOUAhGmXqoEj4g4Y7wK
PUNvCVhKbe2QUUAcdKCl1JND19Vpdo7l0awCub9bsxsO5FYwCnZrmMPuqwJIIs/cjqnnffzofxEq
TaU09UgD0hyrpk8Nu4GUXKjd5GLrOEJ3gTQgWTttC12fUagd1yG9QtEBLdfx6lil9kzw7XovF3Ox
FNUJSN63gtNDy3FZUOc6xLkZ/m14CQZJiGLZzUnjL0GffuYD1ca86hAZZ7FkXHGq0zCCwtySXvKO
uy6rQde9+jnr/eRV4LhHnsguj7XUTbDI1tGUT5y/nesqE9itTEqGxgQqP3nhDtHMA3Q3TkTuMmoB
wm+/1+f8YDLMS5E+YdcnUWI2sIkl86glyZP8VT06F6Fqv+QSm8St/l3ufWLKaO0JmXQvgVms+0iG
swGRN8/qiho52+KWtU0vz6XUUi6jtTHsv9S1L2+/KeQMKxu6KYicEblB9RCbKPgxU2AJyVxXoQnI
Y0lXelMq52DCVPjKvb7+86PPSy0f2B+fyVO4MuPAJuPdYnyPt46LhnulSQnppwXd1M6xHzWUaLlu
uTp2sLwEmWKQ60fH4MRtmOOfVvfvKIfafzsx41CekOLrCDHcgAIvPuZ12BUgEhyZU6YqQ5a4ceG6
OGXAJI/pRYIg1xRn6kAa7LBr6MyDeXaEZhpZzsSYmwxH47s8/s3GLQUBCFkLJyu37+KjQX8PBMX5
KK9Tr8yiL+HppUuQyNw5J9VjqlLyovHfskiwEeHjzT5nWIFnlD5EDH0KhiEnpDN43Pr9S93NPDNQ
YGgwq0jmOpSwAfBOLtksSdORPbn3MYIvG7ZhZj2v2B1+PkEWjsO8PhI8iaRO2dFAheNI7yVBIhSo
yWK1yP5NQWgFzlUkdJqT60RmmN8Qw6wVXfn5Bd82Whf/MxIQ9t2/G5xeZalXTDBcjC1DI+hqhoQC
gg/p5eshrs3QWhl56BwwJpDE140HATNq58NxDOfgB0PZQ8szu11sydLawr+T5B2OoDuKPHebVlqx
HwOJqVntq47wyB+bgK1JvsMPP3DEcvEbN64C09NHone94DWF++aOSlwYxLxT9AY2WW/kUzEn2lvu
VL8sEmG1zZQ3RPrHF9FPyIGl/LfV8rc1bYRhK4IcoCfLSfjqnPVj3jEp8rwNcaPyh74NxVckNX9K
ngx1+tQqky9WwxRvibZ+nggnuu96rh3rT3MKpZR3NRIs6G7trcRwNJEdpqA9hbxOmqXl5pB2/mPP
Y8lfLqRYfG9bQGq7JcqElZJnn3wfSM4v8dGKFYwpJI46gt1bfiWkYJSdGN+56Wxd/eT6sDvahMx/
rdeYQdalfCkL/0Istesbvm5QcqZThk8Z/V/716oYMd0jtkpH7PZRItSFAhjK2fxYP38rIuGU/m8I
qhFReUMjF/lldagIC3h3mVivnloG1gEk06JhFp8ynLjrXj5gX8/tI3THaHpA4RXe2NRNZ36k87vQ
CHKPxprzuCOKhOmMhN02wDzSKwOnAUj7NFkat2spuyxGRY20z1ieSPIbhbqUlzRddCCYWEC3YBWG
y4OpyM6TrRVcO5vIWXpMEsEuFzngNsPjhwMsxlRFadudX9Mz31jcGhVM50cCkciH/TFdLG810Z77
x5g+gNZiYEpPMgJdWIBZwM9UJV/S6jl0khdPbjdPSm3Li3mWqEAeW6OHKwUD2mNDzAXI3t6pMUC+
N3j6c4Dge2PX9vz0i5e6sbhPGuT7SdHkZpmwr1DKYR2aPXj4jQs/zXmvG7QbBmNeuEcF26Wn7WDC
joculaqc5nVTaEmyJWQ8XdwAoIhkWMCKmAnVUVCdmdNva7n+DYgwXteGT5Hk8XuGQujxMS8kjgkA
VFnDEteCKSaR27ikZ0I7xmVw9eiFdZ27Wthhlg3VGBPn17nbreSXt2vXVZ5QJ1cVtB23XeOR0k7H
+imnJ0LIhc3OWjayVhzmxhtVWpbteBXxQshHg0fEkFR1unNLlCb8twr50ghIlztamUeA47smkkhE
GgPzEev5VRNsKEpkudLLA5Fug0d5c2B7PMSExKynrmqYJnkVD6HtH9P16D4HoXFUk9sd3zlNGlSg
a4cDLp5Zz7PpGmwPAUmjpkgQXa6JTuA/KX7iPXpDG4GCGSj9iFwvqBFarDW63gU0OjrkQMdNWire
IF7weeWTNxxKiBIyLWC3yK/S1Ee+Fn/eKhrc7y5tK9N38MBFdQRcmCIdFGuACbhu1cT1dcRdqq8N
0sFx4RkoOw5/AOlvZ8b1s4Pjk4xdcQ8xQ8gl5+hw7Ma+ux1/P4WTO4chofQ+0zu0rfmCR0+evt9/
uxw99j5FxGVq27YJ5xw3gb8zrOje6yx8SA/lopuxM4dODzFuQghPHiyogM56lscfS/QYiu0tRHBN
llvrnXNv1qdFuC9I4ZYqHtHq5qunURB/k+AcKv0yl2w9Kw/7iODOynB5eNFkoU/orGtnrX6MF3+9
IwRMMx2sE4cXZQtekT7o+VIxfO6SA7Rnk+F3WIbB7j8fqJToqjLFOjBrbBDBuwlnAtfkCzZl3pCt
zk+Zy2ZHSns8NhNvoQq6h0Z5DHzsiAtvioGj1oTe7aAij789bwZTDkyMmR0a5gPZxcc1QHHkYaN8
g67z4bsiWkcjbEKy51A4whR7Jbo0ewZd/sjyiJNiYooXhJcdTAOKvxYt+u6A0dBOnE5ewUmZAC4Y
esMliDocS9H0slgMUOO+rVTFfky/YRZ5opj4SgVXTm/W2K7SacmtHM5Igb3PrsK8A7ulDPw6oXjE
jb4VHQ2IpMMdADOSX/vvFKEjLTjMu0HYScdmOqtVLPcCmhWHpTjlvT3tNLh/18LpSwWpIPAIdH5j
TcdL404ozpSaz3qO3rQ0L9iGuJTlH7VH1DG1fid3g/TDTEVEiMkyUsUn4MR6MpBqkTQt0tKxCBCD
Z6PMaKQS63GHdnxlFN0K9t84hT2aBc0DmkSQt0gE5TIWJ3iPkz1PKANgNQoymp02xrMDs00DNdo8
OEYO7jAmqzAJoRncSi3GWx+OtdLijP2dtIN1C31LjlPF2lynyDeCUvFZh9PyUxy7cSXSWU1exk/2
Ks/ydGCAB8nkql7ifpzAwLLSD3WPYzAPNgNgk2wBv8x5O2pv/nDJJdmVBVy4XU1C1f31GRkSeduJ
+A6mIXnUoAsB9RMtd+dSaiih0dSJk+V8GdPC6aMtFD5beWU0+L0t+3lFm5zBDK0InMZRXaD2CF/I
1Cx0T6xjPDa9pDu1c4Vrk6O3lMoVW5+JNt66xk5qb53UyWne41Cr1141zGmVDxiFnh2j12HYXdB6
WQ2KwqZctfR7ZTJfz0TxHepz8erXhLP8Phc18EV1oKIr6Kb7X/GrJa0NrmdxyKgDTE6dXtmFm27H
AKkpSAk1lgETrLzaamA4nSaZYArYFJpmkRaadytmjpJZU0Zel85btD9bKh5lJckXlQGJGypPu1vU
BI5faMMYZzz+fY5Whu9ExQVrhD1/8F5qc4m6OhMpmEEcl0PV7nB0hU7pDI6dqhEVpK4vW0cfUx1y
ujoenlPdUiaOrNzuu2e3x46DUMKXqr5A0kK414njQpyY2fqBlAAVry0fNO8iFQnGAfqiSUTX2nZX
1jnKuqQ6Y5BiKqsjTz/o7AlLlFcWZG1lVcsbT7sCSKC8JB2IDBBY6vXjohHl9pbbH/bTTEREK+e2
oB6X5ZSkAmX+8NlPrzCLIPYf23nZDWDNom6d1eYH+Qcr4db1qJVYJMyo2KfvL5skYphKYo424Mte
FwiHflrVrPrMjGd5uqaUNi8I4jurBvJPhhD+ypcs167+HOjSaw5WI8Q31pbT5VWFqROzQAq3ejaP
ROk8+gzhgvL2LQt6pgObxzI1Z35DfCS/9G5lzabHSL9NbkYXOharBVZoUtbRDxb7m8xbQJoVSaMA
To+baYtKnS7l7zmfaGBHSJCHb4plnLB45CTy6Lo5IR2L/tMdpqYksVu3mxsXAEdZWiHu19TrC56Y
5tgdneQj75Y27Sj/5I0kOzZK73q3dtFJSl7iSVDWlDh5E1pDLf5KNFlJn5M7gWMT4N85vehjomkt
UVQ9sktuzkiCBUmO9SQ5Qpms9V5/jMfvmRGHMeGaM+D0JN6daaGziN4wVyuVL78+ZX/JQbFqRq05
s7G3gmgZxv6yAmIYDVt0jd7S+qihgfBZTAMVCuNUOSalVq3XOyCx0roRJ3t/5sh24F9bQRithqg9
sC7ITy0++nvYosQ3Dh35OUMPodLNo1aKE+msA32o0PD4q+ZatKU2mO1q7EpVV3WhNBa/8D8t2oGn
+1EPvsTjl3rMZfhZmST3Tj3YRkSqdMnhfxCwQoEOT1eyfDMBwj6ktRjG2dl+MMhaaoDhJPKFxMdv
oU5ty5y6OpEtf4mapVECqLUQuocpD2yvCxWYOC942KBnhi8GXEgsTvGrI3COWY/nHY7VsaK00XQM
EY4KkRH4UEIJZln1JMq2LKnVerun/GVsISP1T/30y+PcpuwJxqw1VdpEsR6gytNZyqhF20glVrVV
FJfDKL6UnQlq2I1hKNhUb58LBM/KgZvcdcGlEyhEH4zMgFd+LLDwcfheRVxcfcff4cg1QMG48wQy
J1hDmVtNmoetNKSkzCTLwe5I4Y2JBBSCFBsygIkEwKC7NDv6YqimWJpCYY5y3J2e5vc0IhHYLtz3
vKoV90gDakFpr56ed4efLxj7wIH4FcEy6wXmLVH8n6LvcyDAOS/Y3227V4lm65JPyTSZ3eycji2d
+khd9445/F+Y9atkRtFcTlglKkvpK0W/w2z4XKA/i0dkbpxgbuEWMsZYgvYYTPWIhMJKFCp/Ycm5
amcnUsvcyki9SEV/CoNmCum8gKbav6TT2GAYMbmmkEkccn08VIgHlQZm8Ya9CmNvXZVGpCox19JP
E9Tpw7yAVMdsPUuz007cJHpkg9bW37jDyWeBeluHvNBJMSeR3z6+JnWr4rRPJ/JAE7aYMXnJSDsg
fhGVxyCZKak8VB+Mc4PVkCyDFndQAqxKCZPbE9ZeSalHS7nb3uH+0JdDBYNJZAJoPPUcuLScXb8i
ZiPvGMCXZrKnspwEADv2gOaXZ3nn4p1q525YMbjoHzC7UPpBvpIi78VNOw8+2BvjX3K33INs9emA
DM1jIZJTiB5Kku3YQuHuQsTKA+J30eCvOCKG9yzK+JKQOPM0S7DE7YYNcvnWZikX6HoOcmXFGpEv
OQ9BWhkjaG03zgsnwjSFE0onApwYdXbqdkBrOwXSNPxvk8pZajB44H1NqHq2B6inFXWJz5ZSNu6R
flE8heawEVbwCAy0Wa8voljfQgidvkEV68PQzw205hMph49prHF40dJz4m4i8GMliHMsM6YUeiYZ
TssCyi6TE//p1eIpmKN6RHqTefA740tVk/+JwBlFpoBebBevVxnKDfyV2dVfIzO79zVYBgbuiFsd
kfXLiEyGyIRS9DFBzhiXoHB8hWfAVNi7MaX07Ke/h+tsn6sRuoeo9V2GvFtY7EwJtckwoHfQ4g3b
WqMhykvozpptX+eV4GjLYlQQQc9jCHp19KJJc8h0/OfHcWDZ+58xR84+iAUf7AibTQC3mXsk4sfH
KlP3udD/Lv0M2+KEzOdErHqaZNS1O5zNaU097xmgeCTloEIXxCiR4VyZW7Yh0qKiNZk8gMx5Lu7n
5q4Ui52TkyzCfnWwAY0ssD6dCK5pUOisvdWK8fVDerHNz9dIeenfx7CnHyUCVPsvB+Zi2r2jL2aQ
f5DRLX3sXTRvSw7Pjy37og7PTUt+7PeRUqf45RQHX4cUlqBVTqZYPP6ErjN4So6qSogamKZL2Grj
uIMx0sTAgwdMcs30qM+K0WYFauKmwMC6kYIfgpPfat8YhpZMKh7ZEspgcjtsKhHyp4TTCTtP99m+
r0QIm/WlN4DrOTNXcsGUzJFPhV7q7TG5L7U8fi9om315sbu/W3oI9eeN0Jb0n6NjDZnVCXLAch7M
8SXluBYh0UxTTGJncS03t8c0xK+Z5y/eDj4QGR+obikBejulRe8P7/1SV2H/HRPjHL1NVhOaEWm9
mhO3yHsGsG/+SzKQpID9zOv1MwbdAmHBojJkoJVRN/Ozc7FOq6dfnddK9aEhGu3MOy3AIylwZjqp
+KGhEGqSZv2ksoZhDLzlrsV1Of0T1NVSUjG2rlqnWgTJ0N7ssiWzL7T3w+W04etoDnnHZVsSokt3
s7qO7dqEgxQOcbFVp1AR1fNFRANZy7PCEWI7fmfMCWIZDd47v7fQBkEMm6muwCHnPcMvvy886OVZ
NrFpR6meDCJnCTp0lLDoBxKl4U0BtCjBZm4C5HHo4XCZa739Z5L3E++qqRkAEp48OBO0i2pfhbDi
AwTqm4w120jJv6eghuZnwYA/v7t7V/QPQWG9nxuXEaawq2zk2l2Ivlu+S+A+0ywbNhX3KGpbKyMd
5CvQ/b1DN5iKMCG+3Lh5swxXIhc1txi7h83S4ImGZLAIQZSp1ZO/UuP8rZiGNurFg/TP0bRPLpNS
eVW/XdJk64Ad3992+QpX6CmjN+8hyjdtMZ4dBD6pEc8Lzrdd9YtekIYqVzOB1xp1O0M8rcuGxWvO
T7zc4/TaU7KGhaFRMyNYXgM9ocxIKavk5QeU2oFNB+Y08USm20XBXhfc5kt0mjEwVOrUa3SLo7Hs
0S9w2a/SFPv10UEzcilycysPGLGIDSMQ4JH5Xfqh6YTIZlC9bspOK+jSK3dySxWhu8PKIh5Hvken
ZZsQDgfiZJxW9IdjSZcvPmtAQJ/5tGzPDD/3q0f57DX7SvzjcnNja1Do/dUY78mD9ZZB6XP6JZ4t
jZ9SdcjuDGVSFRrWXQNke1uz3xdRUjTqd8OppXNXWrdFKrmr+ncm2/2Pyf11bPhUQQR4o7zV1kj9
7a0gvZppOIYAUxd05lWMZj0IQ6AZ5FKSRv99E0eZwrIh/MmLHiNJWKA5pbdM1y1h3FGkywyW6GnW
RBiVGDTWKLUM1eqiLi6ZY2a9uLrsZEHGviAnMcQqIVs3FqYYQ4CuL4jy8ilJlvzb2ShngzJEaYkI
cqiVDK5ecffvDYQqWy4mLHRSJhKzXMOz018EnVvqwZeqeyiCa//9FbcAc0NGIsRMfyg66oHk/h8G
zJyKa5H6Tg9AjShDdqwnsG6mpiWv1070nIss8AgWEoNWWQsZu57TyEaojb/zBrW0suSri/VdEGXy
I18Skd7F58wn+92zLGp/p/HbcsuIhALL9/n8qzwpP5X0snEsRyX9MrIPMO07C2nmJxgc0COQriNc
+Cci4lX97DcghDVzZwDvAJ8dBw1uxqFCa753l5ifJ1SgmEFfvYUQE1nzH+3FcMAIOKWYD7au1kdz
zaV0HFJPtR0R6Z9PvrreQatzKjB8AErtLBRXv9REHeXDV9fqfjx7XRnhTz+5A+2PLPNcyzI+NvAt
6u9aCJbl+AgZpj4bqtuVZ4EQTD4jQxi4+cUhdJ9DwGcPzNu5uSB3G9Ijo1JysGRp5eUFPGj1cw9M
tvSzpB8lDqd+zEV+mNN0VSQEQKhGD7QGS1g0Q5YJVILPcgglCogXVemHX8H1WNtw9V+4OTmUHBLw
xD32FrnFL1+e4lOOmQxRBpvVTeUrWx8klD2R/t54aed5hB6r1YMxTuJdyHvqS4wTSDq4Yhw+qzKT
QEmf9LbxO3Qoa68io+YdhYUM+6jXPIwxmPXhhtEvOWRavqfIVCFtbJHNrOVDngKSGtu06aDYb3kS
6MpYEYqbmVAWkuTmS4qnFvcmUUwHj90nYPGaG/2OCR143zMttkZXInO7usb66FLapJSGklK2dun7
1zsb1A3xjB72pFtwTTZhBTEDW99PNXsfy4+3h2hdqLUFDre9rrPd2T6PRYw/wg+czDY7o5O1SGXY
tQ2oympT1DmwTw9/8/Hp0mtw6xLSx/z3pdiYw7thbQQcHMv8SQxwKOugO3IJhTzmKCgWpD1J3gqI
1JCePCj9Lsu7SyemVApPT+CPWDZWmIBEJO1gp44ftb7v95Rhkpil5uViZxWKjykleIgVvQ0t92Kg
tT615ZXMlsu6FoKeOGD11uQaDtKZNAEKTfPyaVDjEVxmjPqJk3Mr1isz/n+iz4Cisw5Z8u8GHcQE
0EANAtCIhlygP/kB6kfkqUtM5SgOg93/jHsDo58+E9wkpYhRa0B9S9Hm/m7VUUtM889JxpNALyyn
KzkDu3ImmJGxUe9s2ZzdGLQUlRWjJbrDeSpCPhwttVhiw+Nwyu7cqsLEfFeEQX+WVWnB5vrQdhxH
g4zBavf5uJIn2gz9UUcZdfhKIxyD6+J+xVMCfq/IAHxvgtABu6oHmaYyoqZefCgnDzrK7D5BtpEa
WQcV8O37I0yBXx3XSP8J3UUOr78szhhMTDDSaI/z9ozp0BT5XC5iwPoa3BY2uGsB4Tycldmh+OUo
33r8I1zGtKRcFZqZBbxWGGZiHVY/JsOseXKT2Ms27fWJq/2hvIQg5DoyklxAZ3Ujo93NdZ0tiTZ+
/SQtVdTJY7tNDySyeJKQKxqI8qkppS/+MvFtlaQCSXsY0thAhhLg0K118svO6FNM/kNEmUYJacRg
Pz7h2z4BMiFodaItVGbF80dkT9Z96R0EBvht4m+vrMokVNDGLFZW1Vdv3iKyPebFpSspt6fzyQfd
cQobbMi4hvPLOSAxV8YcyIRT+kmDWCzH+3SzCWSp+Yz9B6/mjDaCULX4Tu9bnGQi74R1CZJCQqfe
xmOx40idaUxPWlCd2tlj2lj2FeQNzDp25uX47Wt2PVOx5gLoP8oL//9OSbbl6GZt27jkZ6ODIkrV
OQm35yNJyE6JOHvgHwn41N2AZWyKgOdA1E9rL6KH6J4AXxyIE56FvCXJ26BOSZrmZjKrQ0/MGOMj
YH+7vnBgQbZ/iZSUoIXDanP9RYhhA5tpNeNJlftQ7KGOX2tr/Fp80CnwLx5Z74IF+Km3d9BU1DHr
Q8ZrVqPxxp42kHNeI4TEYL6wqwHYdxYc714vm4VxcDviD35u5eD6H/oRcW6YQ0eQf3iP7jLNzezC
7bOXUh/MSpHj71cE3wsHatWSXlXMSfH6q8dVdlSk52UQj2j/+Pp+8Pt1ImeCYSG1Rjuu8dQe5utI
jSwl95YuoJX4Zj1xBGVeyyUXefzi1jJkB20kjXbS6lysXShMXCAEPp37zQViDRHcOBBwlpCzGRga
evUr6hKyNbz6glv4fKkvrLuurHZQNfzOQqNgEqYJ69PzfyTGXVTigDntFOANGJToffyU+BdYFwg6
R4AVXtDVTQMHMhdnAPnEKSWcktQl1QBsZPD2U4Y8usNtPTmmlgDATXyPnQLl1vUnsyNzo/FmX4um
gJC66fA8R+S6QwPi+c9zCIeOhpwwpT9qrR6g+xYa6UnMJRvRo06gAwHb0yxhnICzlFFqA1hdbpQT
iLYz7LE19I3BNk5suK9fLY5OsRZy9MiYBiH++Y5/iTF9yM4EC5YXl4YE58S/HmcreHxXWF0oeEQr
vl6pyddLmQ6J5AUhx2Jc+h6vBHwwMzCJJLTj1iNgufmKXBP1f6rAX39beEn29LM3jTpn10ZDgO43
6Gf7PpgJO9Yzlf3Gwvzk/AuBNWrMSI+wvF8hxfSUDaKPCv3HmslIZUyv7+Wq5kcUmF4QfNBegHlY
9EU1PrqQjKvtPwDnLd7//VlKllWBh7zu4bsdTkzNrLTKCXlijKCWcUnT+QyDSAlLpRwx4IwTXMS5
1AeYtBYUy8og9GEIadFKpmrRiGpRhGUMN47flMtcFIvhrkznSN7nUlG3mzcU+mxK6AOZ3cHNlNBH
PhmWiWCnclI4ZBbbvYorbtEK6rf8ZBu9JGJnDe0MDWFJj0t1GxmFD2V6ZjaUGy2+doEksTPWIXLr
XEpJ5Aq3EyPfWfvU4qswdPY4/f4HWib02BIygxYP7rvSi1wDcXaNkypRtJ9aS4wyfp+ZJ1a2f7Bz
/p87LomhwQxbaxo8jG15ZIFkqFpKS8jmB/YH9nto8Z2hNr4XM7P4TS1wN3sM+MneDgHsy8l3xAD0
tC4CvWzOjfaKkEoSMiuiiDb0T2Zc9yskIhmiihyePEDaQQFPoUPA2HGzmbpl6pSaEf2WIKFXeH8P
RwyGWGXKG80hy0w5spAwlc10mwW9OYuWnG9drmMo8K8pfK+H3gfW3XI50A6Dz0Pyc50XlR2S8fcQ
TqyUyR2cxh1KQ+paZrTwUvgaficEPxa7lXBwrtZXyF3KIUk9k90TUr1WZ2Ywwpd2gGp0BojoEAX8
UNgY4LMT+7VDEZOkoYfBtwpBgl4wZpTaWAKa2xxybXAjyaM9eiwkN+5AB8GuHGWxT/0WW6AVkplr
alScVSKz2GCsbggnzfCOfROi2M3aq6bx6DtQ2AxrY278UbuB9PIg36TYhAUuohYZb12N9hZOxfDk
m5VCWj3dQyUjGxcrA0zfvJgH6/xC8pteICYQJIYeEMZoJYRwuWXOZe+6tgGNjk/oKdkqueSnl7Wc
KGqwXcm4eEhilIJxt8vJXBd9RrC1s8mU2hCZpaTcJSRouSuViph+VlYMXip9dJdqQL0zkCvyn3yQ
/uc2TSHhY00VZ8he61I7F9Yy5gNEmMBe65OygiJAlZZWkAsCji5rZkVOF4fp2+bSaqwAiZLetupD
AEF00Ya6TOVWyS2qqv2cYa9sVdHnO8RZWnKOG629FAkRiptnDq4kWS00oeS4aT4sRWzjrwABLYDj
Bi8zEKmzOp0uMkgjULSiyZnxbUd2khO6tu/IKRKHMCerX+iHwKwLyfJm7G9wsNaK6SrHD/KaRMac
JVa5DuA7wYy7dotZaaBPKBRXQZmoPoZbb//0z3aepogXjyNgjZZB60L9FmT6vTZpSZBK0scD33LZ
TE1gqAPgfl2g1ipP1RjaJMD6/eRG+hPU064dRKVi+KY+QiflBj3qeYEMi9c7Y4/22sVuIWQblveJ
T6i3IZOp48Mg+AM7QWCnCxnGWCWtV6jQkz2Jid6vBYg0D4MqXNbuc8aGurnYtYhjAMXwV3FuoGBp
yfpEzBdBLrH3AroDQgsSEDE/e1LfTjGagx356itD4ZV19kmlIzFHDqylW9RU8Hl++SHGScify9b0
E9ToQrPAoboIKYa1uKmxHuvijNy+QRiFno6XZJ2fZwRMYfMY4jl+DNjJNxyQrCq4r3rPnsW3mUVs
k86xnIPHdFeu24K6Gu0eJMKffIPpxmbavdNJtDDAn/IWPEXocVKkkunZmDq1R6TwWA5odngKJ3GW
WVek0BKr3EPfTWxXqghGgG3dvayxOnksp5kiif0jXJvwMdpZ7I2W77BXQTAtpDoXBpSgh84uU5vB
Vy2Z/EXWtN7BvkqDsFYBlkGW5zHnfTW3Qpv92AHlDW0/9HUXN2dkebsN7llAACESj6zBtc9aGX9P
M1lq0t41McTwSEJleE+2xfedivrJtcBCQof04HYZcvUH8mrTBWa6p22n56Xugl4GWh7c2r9tIetR
+Wbmcv8hdGzjwvNhAiNT3tc+2BY51vKmHBWc+HQGulR/tpKs7kHc/pCM4DWG4pf/m9ODDn9/zYvO
VdCpK8yXwHNmZqH/td1T8+qgW2aqghmhyOGurH3p8Ec7BW3+bSeYfRDj5IPM9a/iwX7hR3hptZ/j
InDmpKJDfBx3UcwT14m4k+CIsqNU98bEi0uffbkha37XrLPcQvoyVlWFXSVwectiv4P9mQZfwQTp
6JdViIFb2ntSfiniU7zZvS8s8JmnxP9ieoPpZ1GNF8PJVwL5GAnE4+gqU87dE2WjauD46eqXQpvE
/blBnKkSpRsTKA/pbSVkFTIDXp7APqBmbwatZ+X5BpygR2iVbmHuV8GdfrfNJT0fGSnGzx/CE+9L
l2b17CZnlCbO76mtLQ3oSjcuGy10YAa9Abt5CqcO1O2NMwHNjd5aKZQsqK01Efw/9jxdhsQNCRgm
cwBgFNg6Ntgq712CT4Nb5I1XUzjQyL86i+oZuqCH6XNkcJ8rQlWWnuMr89chy0wBU++Xv/mu2uSF
EN3c+iMBqS/rh6otqTnZ/b6pMHpF1//NGio3UJpY1SOsll3lT88mpi+ZNj7We5sVxltWQ9ky2GNA
acgboAbJpfdrDw9ykFB+GBC7G+UhtX6D9UCZA9aHRg/47xIyX7gAOsL7CThnjVbZw7RA3LC+mtsT
yE+sDy+Le4RJVH6HRZLGLGWPfskKIw2QvmGy55GC31vpTNydOf1CyHaTX0JWMkkp/clTDvCr93sv
Hj/t7kkhKOU6Ak0y1bl9bB7zTScwyMwVHkBv03EV3rd9F4f8aDiCL6JufbyhHBXkyrvqD9Ka1Emf
3b+MfBQ6qrrHRRKugweWKXIpOAPs7vBe5mlZJAQuLrOMyLSYScF8vIL8DpPJoyPXi3xcmqTklqM4
oSGZICyuc7c83XCkOkl5E5cUAoTBLvKFQA1otLhzsnZ29hl+ojIXUB0CW8jBf/UhPzSIqgXK4eKQ
eC1J/+w8Amuv4c8GDi+4Xjq5hLb7IAUnDQRo8oOtXN+QZ7iOB5stLRlLpcqdjKyITHPMDPGtcmmF
lYqZpTI8CsYOmNc54AMewzAOq2YRz1L2kuR8mJwyOSMp0glrGG7fWBt+L1YGD6eHhafuPxwXCh6R
ARzh4jGEzekt0NtuzLoJb5xOGA6Y05pbyMeuUOuBQMLG63vAPBz2hxV68QQD1+sll4yzjhi3xcOE
ph4ECH8wKkJ/SvtUQvbZxp0nHu++LdXCNhU2apmD1KbKlXpr7UjOcXIWquI7HoVLscKFqhqE7BaG
lGLwO15PEV6prAVnfIYdym8ISqIehJ5ufDZbIbylla/WMj1KcA1gai4NHDSDMo+W+5eUXvu0TnTN
0JnvIa2TbZBdprCrXy9xv7srmQda38U6asfN/lJrhkF9Jt/6gQwFldjzhDApx9oF5biBRgVaOCEm
MIVU5uZO2Ey1+RP47eunf/D4LI1Uj/tKne/dMgGJMuTbVRH/l6sVQ4Z+wkmp2WoaU48cvriLOSsW
/l71fTC3XUbgHOSwtTNt/2G681snWa5pUTNHYgonpav4aed6Gt7+cUNh3u0cXWL0ew6i4fEH5Qav
LzhMWkF7z9MsTHh4+NAfuGkOP/rm0+wkcb/FdRQlhFrYj2/epOD33FJAP9MpFzR69CdRam0OX/e+
bYwD+1b8Y0GWnd8TIzxeHAngZZC/jREYS0EVuFiPTypRVa9K+2UIm27BKsCD/AZq+oP+d1jGObyE
EkaqyuRyBsDwIAwHHtD3QNovvKCAjQotsOKTbfHTxCseOqoFkl0rcQZhPORNgZQMSJ7jk2mFu6FU
/Qh/Eth+zEySZmCIQyB9mfPgYlopc+hpLS/9LBisFI7l1H3Y6WEPMAwVzBkza8cHUtV0vIHnFVkN
LWNG8xu6tHMjRrnhk8H6zYzLJyIMfug16Hfc48lwggXzGJR9LMqBc8ZtjBZwQDvpnZXEHCm1YpdS
YvvEzt50lVlWelr8IlrhmWhwuqTIaaBUva2IgMcSXb2P/M3EpDVDo4tOCs5xwk5JkPEUYr1ys5/E
2BR2ENHx6A6U5/VwXDehFJ40yEF5+w197eBByU71u7vod7Yl1Yvf13YgW0e21gVNJOsg7xF4rPdG
6JAUOpb5GjAQQptTqPDNvqYMZCYcHs3kb2aw5Hmik+FOOkEdRjVY9iDWdwfgHHM/5Vw9SUk4HCYW
/Z5kL7dwZiHFi7I2q6NcaZ7eQNXbuOaF5zM/pwrR8hXwC8FSu51U9kV/aH8rKQmT9zqyBREMSZy5
CDesqgR9Ms3AuF+sbvifXVwlcMwNoaaMfUpL09iL1rG75YHiDVhhKB+iH34GFnHw+fm++n8HLEJR
5+lc6o2y8X4Q20YrIxkKU6kO9m/SRMh33zh/vMSakcU7Ayy6ppSdtkfZB4ba9Cu43gXTYue4sh7o
2QDijPslST0q1bTxe0bHyDLAtnffF7qpyUzjDUSmzEf7tsu+8pWZZZCKj6qHIwbyRh7XL1/YThRF
8nHqw/V4jJvs1bez3JguiDp6Y4upwetbzVuz6s4MlSmW5npSHuWKmuSt7gilV1yC6q5Y52KZVxD6
63yxUegpid208MmrF29QnSfcUIh2Z3K3PkhseUYka2/lyhRXXIqfim2TFOIuDFFsgVlDhH8KoUQH
C1n1vwQ4uXuLRzalsLAIm6LmR+VAb+a6RJbEezMnRXMyYVfpGo9eQLGWzEPIIbsmuGVVKL3Pr1zK
AIk+sQFnoRMKsTyOvgriofP0ozD/072Hk226efb0xR2XLukwVJ/gK1mO8JBOl+I/W4tz1xuSyR/H
VkO3VjuRXqPlg4e7negQ2Owzd5d1OHaD4rRbSB3ryZ2ahEcaXpJO2idBUoT+EjyEreYBf8sOpzqm
PnVrHhLqMdli2WaXGI6eW7F9+FP1H2EDKaorvu1LbI75+5ff5GFjjRkGaIh4zDcqxYwH4aBPnILG
RQf8J2yKg7l3OuW/7MsBKwTEpG1xUL0SOZDFeJnGVxW8VzTfT8f6BiPS9lllj70wCTax9K7U3byV
IyvTvdAZQJaZ591ICGM4lNC3ASFNpCkNUzBe9TZc7MSP/kgoKQ3v6DNhqtt1GXkLjC9oBXZC9y98
duY9lnsUVGYRpDbjOpHvmPjryPE/WqibSgpRbEJQb6Sss5OuDllJR73b+bjR0p9qxILNVAN5Xlqb
hbaVzNFHgWEij+UN1eQhuEzJYNzJifVfg51ExhRMu/Or5K+RIBqO3K2tijsnVFHRFhvYzo11WG5T
OwJoXagC1FBzymK5v1lVMCt6d9oIm1uB6nr/t1zHPDbkcR4h3nPv1dwl06+4j7gkTcU5EmnT8k+D
2GB1Z9F6lQDFCSLDnww6pZRhprUhcIjTEYT/woVPr1t0i1zW4crXP/bhPHuP+sjhVXjBv0FV5zkS
c+q9J6ypmlsg7HIEMHjUhp80yq+MmDK11NVvIYS+3jeBMaYsecY3O2CIVI7NqvusdSNgFJn1pE6A
s4tEazfzY44Tbag/yzxEu+aAzCpnkGzK+9AW6PhMdoASdmWfreiEh0Ze6Sf9JSF0iefjbKiblFDS
toG8NJ6PkPKMgQ6mpgP2LVAuUAdqhb3GkJuLCbRsF/edR0bxF3OZVodTGCjBbk6VktjxkHyTe0GJ
Q+LCnNbVeu93nLNFa+8eQiZ7/BVkPTR+1PZXvTMU67U8Uh9lGDVV4ASUiBny/0Er+GjSZsA8Od20
a40mbhpRfK23w9OihM+Nw7ibE4NzhM86KN//y6iE/JeoMhxouce0vRNDcZPF5bTTDW4gj6Utp8N3
T41ePd4iCD3eRIfXWHYNSTNIIPcV33tpqxe9YKS9MzoDnEV6/OctSORIbERHiGZoEHe89vinPmz1
Pl3kYJ7aHLWHqil2pkA/zebRtfk/IRHXSaC+bcdHPH8Xp9ESCRZpyX6Q4UYRfFxV3QlgAbFKGeDJ
mWORTTeGIJbjR652lvpigXhSPo7/okcCKcusSpXS0+iIps2BXXF75oOMjHfi1UVTZdWWVQP/AneC
+/cSjkpZFM71icFpZDcQea9zuJYDCrPlFJ3awg73LUwM6VZMkG+v6D05SjTuOsJbDwkZAUAEpl2r
/Mi8jLV2v8/D6BmL3b28ahnqKyGaLvHZjuzBnGqf/c6sRcS9ZKQ7LGGBW9E2qIGWEQPqrrAw+hjW
O7cf/nkTkDwccSX/T2oUzsk1vaC6UpjpneIW3jWQS/3GK4lrX4g1Lub0AiTmJ+2lTx0xu6wKyNOu
KXCgf3md+Oyx5mSK4Az1U3d/pih2FweumFSasqCVDPCmlJtRiGg05XTMl/JyAimg1jNDCpg/yigI
TSPEoNtLE0OYu05yzbWwYbf+vf24VmXpx3D/NEYXuwLgkeo1FdoDe6GzUesMy7RdX/aPJD6wq9+0
Vhiz4pE7QsZLlI2NjmMB1euHFw7Jy0MOvIkGIm6wCZFaA65+SnwQ+hjTkmU6ZyLreJeqIXHLxIKi
fK/SKRmkbXbVFXVGYJ2CbY26mcIr/M1Rho8WeI3qwgGgmyiV5iYHRRjSDvbLueROQNwLanoHGh4h
/OUKcyPa+nXcbxR7GKrc1NONXpOg5JD/7p+KecdtR/GhB1DSiVLgJtREj6sYb1NuhvEe+DmhHyR7
8MzTh8J8aGnDxPmyCUmNe9pUaKcK6AYraA7Ri+7pHJMF6lum/oF10O3em5xZlKglmEF5K9ME1KO6
0ZXpp3lEvrnTHnukiTR25daBlVYHudHze3jUNh7LMBLve+NhiGT9/rm2JJdnzXTL6V0tLNN3eVso
4cePrc322w8Wk/dOj3/jhfqKv2JzM4j0e/qJ3mWkkb168310weryPVXkarqPzStLE2ZFrijEleV1
LbF0+JuJssH9IaTIgaOWkw29gBuRadt7qYcT//ypxIMKCRKrNMICWpZEtYtNygrhsHD80UfIcaoX
BC+05Q3Kx0XFSsdDZ/8HZw0/JGIGYfCxz75YgrnDNmaFuivywHgtZX0Ad+3qiBLBHkqIp4rZFhE9
VVryAEbXO1MW8Ax9azmFS373SHR9XSbmBedpZeZ40Yf7czovdG2wNnoXNQ4T/aLwWdCCN4wu7c6Q
iboqaXmw17G/27VZNV8ZHdYN5XRgRuFOz40Vhi0aMYsaAbrRvjpQTntNXcFz9mY9iGrB1hh8ribs
tgxr64qjQF2V4RQ6BNx+pO32zCcy/Q4SRaLcqnRHaXgJ1Kj16JVfJ4fbKKN62n1bHWSddaDzWe7s
+wBd8b/tfoVzhq60D/D4kFebAOSWbfjT6LTC1YHPPtoKNid42lGy0aaDYjdzyHiAWJKyIYwOp8OX
bDKKCb0sVDJ+DfCdCKVoGKkEJjn0aESRLji13uERirQpkznrMkfB8Su9jIJUGcLOeNU8RzCWWB+E
I38fBkxpDRU0W3+xvfrDEy4l0DK7I6LwzFe+gURNkfeKFoA4dEFl8I0cUqNOVnyJTOkgNr4bQNHC
PXPRjAUaPCmEEusoRmo5TDYll1xCgsGsruBkMbBxmVA9hItFczTfPRZ34dH4mNSBegawdV530J0k
bDCHpzhs7wBL4uyn4mBBezuo7SeJBFY4mZ8FbdN+wPurSGlJYf6CkP5zYSD6xvxJHKeqmJJX7pDi
OXa4+oz8JCT4PGjyc26J6/o5gzKjdccl1U6oQjDABHbfJgOVIAamBCcMpGhGh3/iSOU1Mb+pnvje
zq/2cMQyjyrpH4Wq6rZ0NzDdefVTuUEQWWb7keyW0Z9pxGjh7UIJs72sAHpWj2N9Qj4gJQcEOsKW
tCL+ux1Ey1URGUOEL8sHrtDpux4inQE4jlpkwOtkh8Tzw2dSU6a8LdcgvIY4SEgLJV1Txaabkg3G
qL5f1HrNztByFoXhccQfObSeFK97yQeXn6MEZ7J9EEx4QL6BRl7NInapFcT4nbMq+KT9NpA9blCE
bOyFOLzaGezp4iv2ds9rummuBuaw0F+Nvpint+EWFS51ZUTNTLuBftYYpOx7300DFdC9FBcrw56E
ngYYgsIfhQK0TJ0/unA2TF3Ys9cXcUK5vfNuQAVUFGX6S3aHk3neRGO2RcMh/sFaKRmmq3P8D33w
zw7vjOa+918Sj9GuFlvU32RFwGCRpDWN44jIIa822YzmgJBCj8JZ4mMuIIWRzdPDT4Iu3l08Rrte
CKCYAG1pfKdBMBeul4pc2qglo6dJqGQ9Fd0UTkrz16LRBqrdFmbkyNYtaYiQYVyM77egH4uiy5Dw
ALlzR0ZH/yEUkJaZeg4oiRaC/xYr3bud4jAaWW8fP19pVqfGRL3TJJevYrfGx+G3Vu9sAVs8BM0v
FlNkgs9lDX7wxjXlceBLu7nmwsYyiajTlUMQWG7GW4LZG7GXSOqwbo0vHgXx36oDTX5uv7mu0CS5
mtNOKmqtVbbbcgbQ1Du3thdxtPy0Yf4JlJN6LyW28RbL0jo+GLcQqE2VM5qByAmCcERTBgxY0htW
PZfdTrPbBGtBF4a0VqkGM6z/NNIhx0CrHvQsHX85QDcRBKSAbl14Hj6zjKEJvwQMxZ7L4BdoYosd
xNlC2wxE1Ffv7MFD6dKHKgtYSnEl8I+FqdfLBeWfFHiXDmAHXfsgo29rCvqStH+tMeo08iUf7mkH
ZskfVN8CAJK5FI2kokBVpfyEjD+v8sd+03ZaYLukLFR/8uyV903eCt3/baVwym7uigGxRIEf57H+
QCI+oCm0X51oNwk8UI0hKrxw+eG8jgbnE6D42bPnDPgGeamkatLykN4aAnnA7C510alv8B2+kUIs
EHhWjerMOB/iyEUL6FwBKB4ZqjqkF/FsBMe1AX+e5UuwidjRBraFCjKVSLwyYkJF/Thrus1T07dV
ROg1G3nGvZtKW+FHhsEi96wlXAfl6ZFeo4tvkbkoypHF4r9opcer059OwvGaLp76nDCfftSHZ6Wq
JYvFy1lkSS1bU2kWzxJtJcQiIeVa4FO1UV49ylUVJKINJGH15dUlWcy0eqJxt6MbZqu6wtcoAflf
zlPRw9X26cQiuwmETLx03YHX75K0eGr6OTaqX0sDK+kg9Bt6bkN94zy1cey2KTBB2aNTNDgBjcet
4p9WnNVVmKKTTLrwRNm/29MBu4Jf0+OWEzPJKJ/rUnNgQR02tMdQN6yZvJ+8g/5X6nsZ9ies+azl
kTsWK/m53hK5YAkJQdrowDDMWoO4wWtmXmZARQ4Hb5/Ubygt9Y76KckSFOAL/J7RLhK2sjceqCGy
LFpHSMcGiuZEpzU8/cV5fCSM2eY3z0BqDgHYhuzBJCHkBFZ25DmV54F2CRnX/qn23nynTZuHdLdo
f3sZuLNftKm3NBUs4hs6ojUEQezH+KNdOWmTIPusxCasHiaXYF96K2MzMfujXn3L1d4bJV7vhn+T
MhfHaqDLpDcqjporZUc63KA22Pj2QRSktsqzvbu0kw/wmtK5Gp6l43CfxL8RSmWseAdPvF6DNtP1
5zknpEhqGZhPWdSSrUbXnVzjPbLgJelZb3XyPGdPiRbE3TxkUhxmD23HEVu05Rw2vqPAxaqfxk3k
vA6B/+1GovZP1QWWJbUCL8cNrxDm4Ych7sOSE3RR446EeOPgo1gMfmKpmXKtEblm6OGgQEh598uw
YyY3MIGX2Mcz0ocvcgwIYg5IAfavENfSMiefjJMsFllCYcxcIXKv02eoHpfs1IC2QHdLT86VMcAj
tFrFPjQxlcoNh8Bqr3YDKXp2kqp258EvEff2iwapnir4PK4atXlsVuhJBl1BbPr629/1mTayJ/5k
CC2XjDrYhUbFvAp5BkGpR8QSUHnvlZN4I5uMoRPdG+IyYcpX800zaZ/21rmC48DhCwZ0zM2ZO73V
lNeFKxbtrDNa1Lllz7NmqYMAa+6mkGMUrTgN27+mPx7jTWf7XEjDBZ/WJauhT1mkwsQ3GzF1MOm4
p8moi2ZJC4cGCh328ddKRMvOnoDFls5qieIaBo9GXy8EtIIxbE1LKs36Am7kzC+MvsAB1MkRdTHp
MSVGiCYEBnO9nlOW5M58KOhwlLdIEUb83j6s3ygBST//lfFHnNBDZA/wLluSA1oR+AISaGW830as
A0okJG/PoUwHoUoAkLKE416aaBWlfgvwaoNlIYYtVAkDI0RRMYjo8o1Gdgb+OppWKiix/Q/WV3KR
KazUma7cKybIcgw+1bzelbJ1PdY3oqcp6P6fI7iu3o0mtv7BbsKuqawt+tix31VAnlADcJRPgXon
vBqgKhhiMjG4p34Lf8i69uCY6e8qwKzV7RQZ/hkvamlqrLFbYoNcV9rH0kIJba7vwJUZhXvtFfZV
gNvC0CNRHaIiorDIxEua2It+DCqBAEyJrLulRNWKVhr1zm0oWS2QiYZ1PBfnmzjnm6ZBBjPEhIwO
a9V4yl4VvNmUUm6YdbaWXxiiDWlIOFO1THBVg53BJC9Dks645fsn2Z0T/aJGmbaYtYknz6LSkcvc
0I767svgDNgP+XFyvsY7EaYMnxMhfMwdh22D0SWP0nkJ7BNJmJxqUKRq63HfOACmNvLQKd1ZxVe4
g5uMVfgcaHA0B9GnKTbHSjZPz/pBX7nYtUzIRfN5o1VJZZdfOzBf0L7jZRUiXqgB7HzzbdKNwNO6
2JLapWY6zNkoq2cpocVYErpbxfcteEICKLAQQ3vpGzP6JaIMmosqhFqgaVzt9aDqRJuT3tw0vO+F
iGwUt0UvrrERWl6RNww+vuiPHsV9TwP2Bsi/H0u69GftNOg7jdlnEXm7hlU9uNiy1379AfmzzWWO
VXRdtg+VcqpyC0sBs2xtTbsNPy1F2a7u3ccA51Xkyf319SxZsQEVeZYCk4ZS4GevQXq+JZqSK/Kv
CuocjJuZDqTqhed520FKyvuEjM8wQ21LeH4i/aDmED/3BqaMhHKJsoBoLt+lK0uFdD0hxgBm8wik
TFgf9/vIjBijEN3tO8T0WRKv4F6+NpOlz3/uuS0dX2HpmatqrGHSKPQE3cqzDFPvib6ThXCq3pfI
SebKQes6i75TBbDoRdAMURkhytFQ4Nyp/1/oOdwUPiq76f8+du9L/XXxnFE0IW7cD/QuOT0l4y/Y
YJCynnD6J0gI/nD0WbatVR4glSF/hMczg2uU8bdDvGJeVUkBR7jVr0XLew9h5fBsjY46sP/EJ1oG
NfevaI4kHp8lHIMwMh0WSdRfBVfiS0BuCQxSK1QtvZr0QVXMgy/582Ly52qDT2YEsALthqoyyPUy
i14oLRbBEL3eG0n/NrMeT5lxXq5gTYmio+cLVGumrR4KL7kQtTd+kEZXlcqUBtggv0zf4QyLtisa
VeXrmhuZxbGUZMAX5MtrDv3RBjYy20BUMmnK0EcFhpldRfsHik5LuzBy674u87jYl/fQUDhBtnhW
XGs5h9uYmRRb7+5KDmlGBYJCoyvOkZG8nmQlYUTNQCDYHyImiyPdMEelRGGU2INMbwB+Gzieu93K
i+Ki4An2r+3CEZ9BdRIEqurpbnBUmYZESuW0rj9Hz7Lx6YcOKOofSX0RHIKzDF74kTzCsyceKr0M
b8IFowggKzP+Cu02BnU7gUZIrkSlZ2kNeXGlzwTX1cAOv8jV6pBD+9hnk/MpRk2Wj6tijAf1K0Gb
7dW9QrVhOByWRbNRF6OVVYQDNlCo7wGFWlYUkXQp62emuu8WWUQNI0VJqAERDGUqDh8HpMtNWkqK
wQBpE4vpLNMQUKr0mUn1jZ1imc/eOJ+lCt+opqwlYGH34aiIwd+SiK9LSIVCr867V7F6mMPNhIDW
s9mDIEw8xjbcAO/ERXO2nZT1KcmJ6+aJaywUnXLly3FWkMKH1PRsv69GpNSo5/ym60lBxJoJf2ut
t9LguaR96wiLk/Rk5msW/8SEECwZvhz3oNeUy7AnKmwXsLu+rb1eIcNqJqGyE3rEDwVaa8MBHZiT
gAWbOmfmM3KBYmHpMGooXnwsIM12VizNAPr/P/bVNmFFGMritawisY4lKbk4BtqSA76cW/lu/ZMf
DZ+vF6cAb2spd+Y0/4jLUHiG/pe4WjYqBNoqY7TBgkuNoZ7qlmPWRtQO+8qtc3psGYZZ5fE2QATP
JOMyAutsORXFy2PcgCXLgZYA8CQg1LCPxIpvA+DCwCXdgSVafSx0/KyhRG625cxwyyDJp0MyLtLa
QognKoFBnNbXhMCaEGCAR9+87j2tq0Bqx/ykwEmUXRVUO2C72vgRG02ocXxwplmcTv5/8+C7O+f6
IGSgwhEYzwAZKiSqUj3cW7Z070kDd0rEKapsowSrm39I8iWMPVXBKZ9prv59TWRg2cKsI1hslaOF
gHiiOk+D5zXsUNr23x9Rj7KQpxpbsXDJPo84UWHJ6Hkk4pyqJLFVX7gJMjmlEyIRwSlmA4XufpLh
GlqFaj+6LC/ex9KMXJXWZ1DmSkYvYUwrOedog2pfLxL/kMrDuHBfH7eZPzF0+n9wwbVPJ6LMzORU
0M2sbJFiAJKPPl84fJDUlQJIarS4WHYJFXy83032dezJNa4MRMX13qiCWxxJccobSmOxc2xzAJaG
3ZJxjE8U9EwQwYabzWTA6NDpBLyWF5bywydWohXHZC1cFoecmeiDSwXqD/tcouqiBMUlTUf0Vm5T
CRDz3ctpnk9seNSzY+Vj7FhVrV59Ep2AggIDwMJA1qvlZKKYGncy2qR/CCRCjKkxlaLULQyQrwIO
19F/NQkrY/PAc3xa6KLLB9kbTewrWy0PFWvDSu6r/AcJcLFhfGYal4uK8IvUuPc49n3ZirvIPjq2
dRMOzlFFDKBEyBcXhYjzCGm9hm/ButXp7Tg9OFaQff/7LVdOKCoLC2xl4XTZDaFa6alCiAE2qX97
b6CW+faRT2cTT21avuYTbdGaDfZExBxeaVyjcIs1M1bAgYhpoztNuhGXCKP15aI6sWnQIoa9E/es
05/dnrUNixYcIFjjWcwmFvrGOxWwbKa5w+yLTEb0bV1PyihfZHsZ6jF6OK33iGmG4i1kI9lPb8Cf
vTlh7UhKC/piXTYdZmM/h5mLyHUuquTUMAqA/FZWjBzFtTeq+7SuLEPmR+HoZqjyHM8qfMeRH/nf
GjPhqRxMz4ozZINkUd6+GufbPgEbs7yfTUpriiSl06o915XOrMpOY6BcJVzQdCOwmJSMXtaGxflU
sMn7XYAbVBd4yu+ebXGzgjApcNIBxPLrxOfJHUapSjfLjIZSgzetC8oOkjVWRQdgCz9cmhwiKxY2
m/bpFIKbakW1cvB9Ufk04HFtT516e4ur7+1NhGdO7h6pVCTXCifLZJWQOF0HnBlsmaKKiMtaTF/+
ZB1RDDB43aFfnTJcvM8Ch0k41GKGuETBRXJks8S/3MzN4OhG9xN6jT1+EPYtP+4y0NALTHYm5SaH
AdAWtG6k31EGB1K1gCtWHnOWjq73VJytKI7pZKHJ+ejeBNFIRm15RFSrYyAkCIIHazD74UuJnhFL
qU5QYu3q36FACg/FoDnnZ+uNFBfCepK8T+ZFOGnqd6omONf20naCGXkdPrAq8CiUyrXyjZFdmavV
rX9f0GMUb+wH4d9L9bCWvbSLt6OACJICOnsQNb3N/KtWYW4sR7rgoJlupKse/GEljHpkzGSRKXvD
0DgIg9IzI4yqCMftyj1IiukZqsggx2bXss8R05xgdPyGErt2zoCXqgxKazj57KLmkPLn0IDtMx+M
HXcCdaIrKsNgxh1So/LCJ5MJt7d+7/p1UlQE0cc/afx5rbFmtxz/3i/4PeKEe45WF+9J2mdLdYOu
vxCtGd0tlCbL0/ubKCO6dh3UJ1xEnhK4imVaotGW5rJalnYuPMaqwQ8d1Abonv5fWEg5xx7uaYOm
NyEXLbKj1EdXr4krxIRVhtwJgfo6aGiFQBuv7CJqMet7WCzggtqY28oz/pMY8fjIB8qwc3O7YoH4
tJKj00E/sdr0TmaY+yy31Zi1DaZs1tzgIXext1nIbtb5kbhSP3LdmRcZCm73qXaPJo38Zwrky+gn
mcwwtUC5OlmEkphRRbH0Q3ckE7G2lbnwxPtjF8+9wfvmVQAeXtvVzLlRgHB/bPYTckLP9LeWX1q3
ZTlmqk6Wvpi/BiTkz+F5V9rdMmv4K5NEV41TesxT7vinI9yVq81QVGZjJ5F9ZPe3eUTZNkuA2Rs7
ih0vTuklusjXq4lyybanFlEXsB/2qnuzmAX12Azm89x+Mbz++g7UF9ql2D/NI+PNscZkNLvdXmJQ
XbZX6RCfQgWRmkScVnJsnIy1USiLt1myJOn6CQ0ZFV6fHAIvPCbL1ey/159jzfYZn0aaOhPcjL3H
Fcs17OGvvFWKO8Zys91uIGfyIUtdU+4neW1KUAJxol7CBU6N1/tizjsbxpcRYbHdTF/c85R7hhB8
8aivw98inr2BGTKczQXelvaKcdssckGVYUu3lNh6qNPTv5DjjrLr/MDeYtkMZI3Hc0/qNngdRQX9
JxlBgVm7+6CsU4HzpEDdfNxK7HJv5Lf1jbpXxdP6YBgr3slk+bPHGzDnjHmk6+aRMqHe7QKAcYhS
uWTBP/ZYx/zJtrhcMhD7WF1BCipazQCxlJk3oHcZEXBdMRVx/XvHLAV3YFnPpmO9pXWmp9NXFAXH
DEtYouqYBA+xWFA9q+clGXVjMsU62ssRTJ4AwCayVU8nuLzTmwPo4uWpsTP6QphfirwDkvSU+Q3W
wJSTS93tVbeywGTq5UNOB6F8iUiCP6UfzVDl+1sTTt+GzBLGjYUUKRQ3dJKUTKNhpupUfoPvjq/b
z3LWe6F0ooJt/J3qPSNv3fq9bF1J6msMLTutGK4grii+2m+TCeUrKIh9Y88yiCE89lUCzbXmkXOd
inatUkkekQKpD9hSDnXC4eqLOV8betjVekVwx01vQQM/1E1f/MbIN5F0FpRxUF+O6mPlSngabUhX
HngmjrrUWG7k5FoMZUFYOQko4FbKlNtiHe+4MjVN4GEKl0TJQ5lj7Fo8gy3zMx5wlTIWfafXNOCL
7hU4QXRO3q1HsXi430Rsqbh4PmU+qW2HEBk7EhnxVFxhyn/88FlkG3rt7qFp9BMmpA7ou+mbijSt
Pi7GwDo2nuWaZ8XBbIej2I334FPLpXAT/16AyEulzYoOdLJofY/IdPiSeTlcE1yHX2uDUxjfEYxd
unck48jY7cZTWx2VDc1xKwJhr+NV5zr7fmiEDJ9M9gfkH2QN+kL5txJqQSNHtgrY2g1uvpQE9I2f
yXCAHRRe2YPFpVvNZ1VCNGjVNEZcd+O2JonEtsGJ7heccfFlGXRnEhgwPFj5b3NheoxbvNrHgxqj
C8uVUxuLfNYaH8jKIdLAMYVblkrkP4B/ABUyU7+KaTMMzeduQMLJAJUCf2xNmUCil3UefPpowk7R
8+ETDeakJrlcap6Wgz9GtFJhKPk+b8vI7ENzqTwmmtfq96uXfxFzZacbAcULTKAAxPpL4ws6lCMI
Oio9gQgm9hXMDmkKGoO9qoMsJUI+o8XPiema5HX8g9/41ifvmZ77FzN8gSdsWOWmsJGM0c3Hxw08
OiriYCalFanxZ2ODPMvuT2VLHCjnPEUCbWO1z69Zaugfpl425OSZEtxHtk3duaU1Smq80OHosldV
Z+SdlmkVTUtloXRCRLo8oYQZZGI983ta194JbJjkXF1kbM6FAlMDneH3xWTpuUtFbh1ku4ZyZDCG
jcNQwgU4QNHNWVOu6zgOBAC7EfCBwG4N/zVuNdkaaVgQqaksIRyAvfWAN5r4MVigBlL9UjzwLZYp
wi4J9LJuPQ2l998X3rFQo1u4B6jRrUgB2YT9jaDWn/5F4u5EIyxO7zUHkP3wuyV6RiKNkG1bj7nn
Pv8V8mIjgLsVVCnGlJqI0+lWprpnQLqgyK5AlsNuj5SOd59VKeaTpe0dmVPuIWoJswa+J4Oht+ge
nib3E8fa4/8UUOTXHdFcE1Ggl3bdToy/WL65cbkhJ8j7GPa37FVp/zvPAhoBwoU9z4I6dKAWb1jd
J7EJnnVuSjBzinjr91d7OZclt/ATCXqmAhKtM/oe3ta7X2JPns4r4RsiXurhf8ld8hUx64FpOtGE
muVPjsEHTEIUYOsxmgPCK6qQdBkwUgc3TTQ3/5K8r6mC723HJvIlVIylhoQoKp7Gq0Y0iJa2+eU5
FvAHNigXduqMpyR5nMEZCx47a/W9zFwl5Urs/efF+0QTtiXTsJbcH3OweTEopO7TOETlfK6yCJLs
DkoHUVV06lwSWUMoH9oOGoyi2lmjcoe3uVYTJ2Sfmt+zYZo69bMmgQhcBkB/3OqMcT2DR4r9WZqT
T4Ee28hLfmct1lwXIOz7PoHH78bMysMlqtrFTSALpSlVjj+ywfSkJjSt3ZhrEdWP+91aUbmCAq2f
oFYV90cbJ98hK/DtJh77Ye4HyGBVSfOCi4Ol9oxI0rRw8lnCnXLzD90dKUdVXJJt0ZQPa1vXZYdT
VSr39cOCuX9I0izqTxCQxKzGJz5PDeWNyNsdKUv1GGFPqTMljb7zCquK2HirN28q47QefyGB9NWx
qyWtp5mNNlAZ1gQ5tWG53sdg8onzdLkFslNWYAeP0u2/iPZJovcF1xrNHkQYigBFmp+hibdRFYKv
OywWvtoEDN2yLHkfuC/K92A5cGxYpteSH9HyStA2+GN1oIL1T/PqRCC5EPXVjrr3TwwX3uuPJmCP
wtDoeKbP+jXBsvuHQNfC1PZNTmrF+kGKjcltXEkRzobPnYLdWs6ejlz1Z3cYpAxPtycd61viSot6
vwUS7OzMrl+65KNg5L3/MFeWWdvqFEqarOSz2vRcP5xleT9iObmAdjf5xBi0qoCx/cguS3AqhDmZ
sJfVqlxd7hQMx3J8S4N1hj6UdG5FGV3X8MtpBZeSI6jzSC0oHxjW/j2tk4W/tH7bWZrBfMMpXXyf
zSRmPx9SHdoVhxBx2uySBjpx1YWTBnefz8nJ9pn1ws1ukR+fofzw+sYF0hBdTWQr5PPpnJoTwFkK
cs3g2s6KZVYh4YVJ2BZZeTUuHqi/Yk00g4Tsvwa1WdwaWSkKcJYtGe5n2StmUkJmIJZQbBwx3XeC
rh4igtOfdYto97i0YJe57JclmbGwiXAUjFySE6hN3iNMHdXcd7YZsYjzCaXQ+pIoD+peoh0giHJ5
LCn7IdfedJ2JsbskjcHoxFlPlOqlI3GNu+Q4OefVBBdxR7tjRWUZ5UGq+NGine/SU1PeHSKP2DDb
Ws/kkCIIWTYqb5Z+/7unbjscyoPZD6XCVkkrFhxgMSUe0/ca/exlR9wqKaPoJMLr86dUg2jkHwYJ
n7qs4Vhcez35mRfiVFellYGWd50EBzXGdCOY9sfcL0fW231sLsnHp/LQYFzLO7BNTejdiLTWK0VR
o2rInl+b55qbsBe5q6Fcrhr2NdmLO+NocT8mxF1vq5vtOpd5yFlMu0FnvuWlUoILw+oitvHt3brX
IMIQ0MccT5GVjPDaX6LV3J/wn4Jn/b+axbbJeBQpXcLMtT3lW3jFWISeNnNYAXH0WiEnV/ML9+Nk
1flTfePGBdtfVtzJiiMg6KlQ2XogQqZDNu75J58Gf3IgGUaOCK5NP0d6g0Vaho2vw/eLpoMUBsiU
T7reaHHwFnLdXSXqnw3f+7PY5xLZEnk3/ZIHyg5XwZPvr6T8ehp7n7W+j53CMSrqVL0/fg119OsL
odkxIc6c2OiONo2/kDmZ28whCoFmHARa33q7AqRU5gRlUK0F12I+lNaXUmRYIPOlQaAbicM+Ogql
S16VhikHYAdthfbtkgka7GudClG3MXWT9+U/UmhPewobrHegRIc0IkSMx283rc2ihzEvStIeRxmn
7dnP3D+C6cYjsev0nvD8OwX7yzBhLyfGLCjSOJ4yt1GJGchwarS++cB261IChsgh9tzdReS3AjPR
jiWfYjgHCfVsVTmhyDkXIPYJZ2rZxzY0FIQ22p43jaus5PFQhY0A7ofsaaSnt+yc2rrp3t+uGTuv
dwsVQJs+frSWw/obHS7hYCxp9C28Gkis0K65p8mXI+XLqbMUEuP939Kruu5a7t2yvc4ZNgoDLp0g
H3zcG1iKmhrViL1QRnZY+7/GTjIod6sTN8l8/npm1q5vS/q33Lp1UnjkhhRoFlG5Qv9IBvQsZcqP
TAuXjU5wHMLQT4M12x7c4woVWn1SyFWGtXXvPoYuw8Kr3ELx/eKvGFczbmku7oQiVLW8Z7oXrNHt
EIYxSd/9VcDewzHekwo2KBS36b9+CQVCPbe2HtpfIEMAOAUmjpjpN7a7It9241JfMZ/JiRTbbkZH
JVYodA2vh97LuJrfI3Z7Io25nhChKmynilVcon2oJfdR5XkTPZVEWcH0EGY2QShFBDIYBDpMC1MD
4oO+fNdvEyPOoF796//iN/svBbKQURmKzdEDtQ+FSe2QblCRgE44FIX1ZTkt//20n6Nm4eChcNkU
z0g57FGoK7g5p99ehjPpuFnCLZyTMphQ8/00PdpTCvw20iuIITK/aXzxjQaNyX/1PwyoSl1/LYDO
t4bMMbZ7hbT5DiWWAhw2nmjhZ3rxtTvwmmFhI0Vac6b/Z6gCRj+/AO0qlm3Jzk8CRWLyvxcCew5R
Aa0lLsOye+aTnPtLmwRkFkn2el2Fs2m0kg/ToLswWvFEnplu0JOfAoWpoLFXaItfAsZZw6fTa/+H
iHdAyLwfYjGASk+t2l5IBh6pBExXKZojcFzcdiWlGnQXoZPgQF508qAySqsxlr05r5ws3gWDQ3nW
Qq7k7tWemZzSUJQHqxSa1XLsYWYTi3YXpS6W+4ucoU+XsI7TRocYQEzVUQIrXVscQ1FneJwviErj
b2dlMRIbwJYRXJ06kvuzIKLEVGoir+Cgef9hsLT8hVX2mD/bKEoDTsmTpcQcyKqOkNFiIYTUAXSA
t09q4xitmzEvh9/Oy34Vwh9Bd50m3+TFXqpARsUxNhZSQ1DMvAGYtYE9xsoez1P06KKjZ1+o6doc
8akFNODWf6YgqqmT1+DXfxWeFjBhcLGkrEUjrCRlU5J71yok70JJ2ZR2NuxK9HFZpNzlAnZuQnUh
+wCNdhYPcUPPBev7FkjUgx9hD792y4eRE3/VmGLo42+4D9bb668L0jsROVD3F9rxHCaTBbpwsyNY
T252i/NFY2Jm3nWzxpH8KqnCLA/guNwqpR2/3wsYaDbcYq0gltLgoD1H1BKEZvU8LycUevy0QFn1
sT8oiMvWOOLE7fONMSzP/1870yKV1XKHzaSBnoYCGMwZFyQqF+PEXR5xaS1ddbnJaR2W0MDO7IuG
Jd/cF2QOjAUALnELGE/aiupKeqcKNvCFbRuAn0+JzQg4shSLlcp/mWLu8LV8gJw8r+HrwK9aFIVq
ljKwMJNi0+q2YIKUIPNOOSDEK3VoY27FVGYP5yy+YZ2xcE2aDVc/DKD8M9EYGlw0LkRs9L90Qy4+
d0MyQBA3+6DTLbH3XGTntWsU5ht3yDCXKEZuzvsQ6DmpGwe97DKgUvuBgUwzCgvGZgTBMroxcYdV
wzZoiKyYYg+gJyJpHGnfzR24kcBLJTe3oDwYyUxdo/kJaNmjz/TBZXltfZ4RffzOveoZc/c/croF
OIc5kU0VFfLg14m7qXPyidrZ8quwfwYL1ntORyRXaPJrat1RNbFBUtphEGGxFtkqkB3qWdnVhCTa
H4NE42Cff4tTY3ZhmcBqpxJ83G4zePBuico6eAir56iq3wSGnFaN2TkNWZltMQTIAXCiiZSA36nS
1eOdbK9+csk2xrgG0ecbkXNh1yElt+g38wu1J3os4Arh5dg8P1+6l4ll0/irCoEYGzIwBtgBO/ip
uZAbdpeYiEhYx9KXgVqN2kOVsKeWONCJgnqyB/HMmhuMoCN84MXxdrNOupNE8GWUCy1pe758q74K
R7+W/MkmFOayuFzr8rA1IbHK7yQEO10J5bsd0DAOrj316tJxMwhs5ONSiUCx6mvKVyIX1dB/JT76
ALeYkU/i9+79hw9AvcjpUiZcQSC98Jl/qAAJ0r2/A5tc6pyObsPxBCT3OLim9B1eQZqZ/BMHLOqc
FR3vrxoJytlNmmiN5ypI1oRJuQasxXhHSPwaatyNlwra2sme1DydX4wsasl8npkdGLo9rJslstUs
f1GnFKW3pPKOD4Z6nqxHtoujkhI/aK79mvq9xy7hEqO+bdToW0j32P98jIv83hK5VMDJQokXmW2O
6s8Nop7LKizxAxY26Vq79MCeAhJHd8r5GeOdForiSNcvxZNIBRov1bzKXCQo3bY077I/xA4IT92Z
06EbhqO2mhIKdEtwvEcJxVuhKrq+j5ZhFeEYq9G4CFEv5qMX5tx2bmZrSjvM5nKbpdM3jfXuTThT
lOWq1x+e723SHDdPaZ5BXR2jH5E44THoL176n48bTIQ8PhpQhk9od1ngsmx21HXYkiuWJUhOgt1s
HJy2WocjN/JI5aobD5bOF2Pf4YJPh0yKeueGgKo7xv2YuCF1U8jplqiPC/P4GhnRplcHW04XH1tU
0G0oGQcB+IBqPJxJZCv2eKWtrJ5YtlCau6Ip2i7/4LPui3qGIoW042yKm6ipOcSI8nzpVzWNbvAR
8ROxvpYX/PRjW3wQkyn0ZtBajE4gNi75xOhz2kqBP1UgxEC7QoVGSlIawbkKxul3BhZMPCz8ZxTV
Rf+T3/wlv5GDBgNjUytae4W+fhtGXlirmPm4DsMJ1s8gAjguCsGEXop21GI4MVDm/iNmPSq6dfHA
eQOaMDTF2UPEmeFD17cMjMe6pxIqgdS3rPSRFvCMRkr3/f7yhtPOUKzZqqERRODsPqCf2wVIzEq/
p/GNrivURVLgDm96GyaDe3BB7+I0SZgNAVnUWsKBP0YOqgg8DwjLYig2wHAdIIbBfihVMtwVfeTV
fash4Nf0iRmRdOqf+7emPX6uqVp6i24cO+bZRmAoLWJxcC65fuqvCsptgLysIC7+kk1QKtspHj/Q
uM9FyQv7oqggQZMOQldo9vzKVY1/cvrGRvZEJTFCvSCceFisX0n6lDVnWfRcbSccCOvr2nKS9p9Q
CvEf9TrSCubTmST06aWeUkYqonCh2h923c4ARWeabMYuf9ae7QEk6CS4DB6HRLOex8m+TdbWeV8G
BEDAQDAlnqs3LZ3Mu8ldsq+U1bRi4QeVKz0TeqPD2wEgGMZMQyRm3KYWr41DzsTSagUu+XdhWkRy
rQYMZU6z4A/BvTGb9iv+b/nsEEBv/r+3sa3ej0tToYc30Avc2pbc/DhHDLLeoEQQLT4litdPIJfr
inQ+QCVGT8wZ4RI2eNVcwi98pjOmohWn8M2DkWDaRPSYb3Ee9Y4utN6io6YAplvLEcRAh3tB7shV
Bd73PZw9S1A2iBQ9eyEyBZmlocJXyrwCoAgW90dIqM0N1Bj+UR/RRbMX6RmdErGX6pMDzNki5af5
lUSRF+pPC9iXKv2rtsV13VCTG7P6L+i1QMXsbWgIzpkOq0RcxpBOXes2djnvMecjUw0UFbs5m8zE
rceTi8IiJgx5GExPV+FDnyr+6i1D/LVSIDZ9S+cLm7+Anbfy70YIJsT3pTN/vi3o2NcIcAPyWU3X
M2MGKYJtXCRciMLTREQJpIpLSYzNNkl+iYGY3XuHsqUDAhx+ctXU7A15aQPd5tBDNcnzUTubLOM1
9ccPbtNPaZxHKiz/iW1irBnVkO26nZsK9x7Blh74O53aJYJSbKyy8rd9DgFpb0drkmXelIBonxVc
y1CI0VkRF9dMHkDIQ6A7LzbjvVOyCxJEVFK/c3zivjxjfOgCCVqihgdKJzkWC7AtD7F8RIr3Qj7r
3RwQ1g0tgS0PCPAspqLGF9BODP7WdUNPF+Mcs2QkzOMd0JyDf90kssIQNc7B0bRkGnI1kSZv149a
9Gq4aE7Y3zbmfTpLmT8C5KYC8UfePdWkIfkPkBItZIahaNI81iupO6f9lcwaSxDU2LoEjSlR6SKY
u+a0BRkz5BVCtynobPYpJxVGXQ+0rS3iKs1b79Zzejd6Y7r4wNrgI0pny+jhaA3k60+wRFQwNoz6
EXEeoNyYaP0gpJ5rmNBQy5Rykzien9Inacpte26WPF64eGxdgZ42gtMU4BzedvdvFSwH4G+SwCd9
6mMyU2uUE3najwGZpVTzP381vYYPhk4A3SpvEwLokEYUCbAshqjnPSKPZCOjT2UOtZd02zq/qRPD
oSpBMhovMlcK8WlxVi8Pe/a4+tXc95C3xlPAzUp6USvrUp8JfGlg4ufi3NcLLXKpm7Iy5byfDfmr
pr31UmSGHuCyaqS7FC0D54vKXg3OWKeiO4XW+Kz6OrUTQlQ+Lm+qimmqVtJfWwztXYGP59gPvQRZ
DpAxY1/TeVuHSe+i25nwkbtqjAr76Hb3lMZVt8rzUhTQCZ5pqyIvD47K4Lr321EByEO1oBjICuJb
u02x6DhMI7E+hZMHVZsTetTk7xBZBlxmTAnLN4GfSsQL/p7A55s5LxTZxW8hIok+KhAW6dI9o6X7
ekpuqrZiTWXZToHdIrehpQKKAh/iBxqNMX9KmvYRfA2/tTmiLp8Zr/PFioKdmCvw1X3vnD6Us9JA
XrQX2jjRzfszM4Yo1QmcmkDGZ4lttnXe4IdAiyyF+f34SHF3EVTd/hQWt4ny+mxg9/ksDTfaczv6
vRD5Qu280B3KkFJVbWNULPHXM1U4SY+aZviqTestPg71VI4A5X727EtsQ2Op1emqDH5N9co3YxQS
onhbw4AFttiD/reBrFVJRRe3ReqceHVRfyt3Zbhv+bclysLn3ktPA9DXFRIs23aIThXysscBr49E
XfbOILbLjCM/jguWBg44DwLuPWCniM9jPXq3wkX1XWAGTLWnQMcnvwSRFQLNROedtdl2DWnMA0zV
n1UcP/nebt0lZO4vcPPJERLxJE9UkFj0u21UpTJ7YlKWiQi8uqOqrFcSNmZnoV/m5zyA5ltPTDG9
xF1CVLzl11tuVSkuHdUA58ykGrnppaZ/vPMjZU4OICmPITqhxhkUzYci1Jkt8GV61TDE/NODDfmZ
HZtym43pVA51qaObI3EDdse13GxOCVsXNS3dtSOMWXEm/xHw/USYh03UYDlYJYSEPxiGP4jFIbvg
vqERu5wsjKfKwvQ/+n/nsvLeiAiw2adm0pp+62hZJV8AksxBmEq729sgpGPE/BGj6kyZqb0rjIHr
nr86OyWuhE7bjXVlQH4WlgQ1zhSLnjiDnvWmGYtGV/1J0l8pAoAGq87hHV+IFq/vy1R9jP0oI6kF
lwPlkjRWAHtYAbD59PyCFIt10Xyy3N6cdG6QAYovDZ2tXAirXOE/BLlY8Fj3Acf/XLlvvNepL1Ia
xW18+TjrMOV0tqnonqQCt3yRF09pXKoqmqKgJIXwSw+3VdNy4PBkaldS4iX/qyXDSaUejWrz+Pc0
20aCdqq3qq18fdJbTYpqjM9ldIdrCAfVg+4ihww7VAZQUyJEkKa4PLo6FgsgccgcYDvjOv6KKCm8
JmL2aPwbqJDf2itmtiESZjZBhKV/qIG6PJBAFoPkpO2g8pLZQmPOVYJjU2zSL4qYL8LoKy+kJDIh
4PqeLoqrrhQ+pZbw+SIbl9X2KSzrj9qXtiV0NDr+aVtHWMsSWtaCiyvvMJKTyjmHIcyJ782K3ggJ
rxi5kb+V7IuJHwr5C+zVOiZ3d/3Wa2Ya/u6Nq9XyOOLU/whXwAPX3pAAsIj9krS4ehE+v+5zqwxs
JE+P7fU65rdm6r3OquchYIQ/9dNluyqfYD396Rsqynks09om+/YQaeNc1vWJzsuSDc+wqZ6azIbl
OV3OGxF/oJ0ogffiBTV2Rmcdu9sMRYsbMpmkWMGfgfUvV+CCRPAt9attmkFyuDN7GA7YuaXTMn+o
h2E1BhmLWIsCNMSmMBLIZPic3JaMoMGTOs+Fir1c3B1IgLIfQ6TB9rjKf1o7wGBS56WZGMY9VU+o
ghzkU2X56EIazfepRYFKVFy+X2p/HILF833kue3KsnJdX+vDRTKBFra7lJ+Y/3vUI7WjUVFMmeej
xPCKx+3zFAmWf8Z2qENm2Jy5rBuKxIANPv4UnCjauVhgDmtLd41n9Pfw0tV4O9/CE2MWDuK7zYwj
Xzext0lY2IcmIlVddtkyt1mE8eveB6dQBq/j7gKdSUB+cz8XromFfcijQOGRTAKP0A7CoUvkCNLR
/KsyuC1KfwKR+30mwUZJU7cMZPdr+KJWmrJR+TUvtMcIamgFBotrR3Hu2Kxb0bxFNqNj64paRIu7
3aWn8HdSnAy2WM1nSIuBQ6RyT/kduyOaV8ik68WAFPFTP+I04tKqp6wrKhIXlgZZ4QC4KLI9+pVl
CWx6+VySr3SOfY4cycMKWLnUz8QnaY97KCCV08D8k1yK1edBpy/2Z5DzdSBJm2HPDVXQmo70HKQT
FpTZ0AxCWIxAFUX2XPfXVka/yyTizvM0vHpWZUomP+L1Dd68iQWYjua4nnA+XcFOkkrrSs5gKGaL
QSMFVqVrXvEaj46SzqKNHiPQZbENJg9Qhgcy6LmF3343lO0gIuet8Y5+jwTCLhOTLZOz9zqBu8Cc
7cx/8ewBSYEDORSj5mLTl4Rpvr1fHFpv6VYUS3mDnMbevASrftm0CKBs7/PoQSZDFSTSsS35Dek3
M8aRzE5H65e7kp1QYfNsyTO1vMYqCI1Eg0BnjfGn2F5JF20F6FOnutwhkxA1XtUfL82U7JybjFOL
eFHivHkPnKvpgIgtruHFPlvdZYXbcMKC3moU9D+xIheAN/UupdbcSnXOj7cYKIq29iRViQL0rIPe
+qF4cnypCmgLPlhv6tFVBHy74aSREtk+Ip8E6Hz2RIkhijJ75LnQUFK5HazyEv8xqvBajEb7aJbZ
lnh1O9b8r+Jal7OvSaCzv4P0Iqzy9be1KynA/lSU22uS8sUabwUbPbN2T1/lIwoELbOYgS+/gIly
CQeZqaYEEtgmGy4ylX8tiMGyPmLC9FUaN4nKXZfXwpuaqufGNGE5HE73gX6xOWpeb6NfT0dKkAAK
L5oQ2wInn4cDF2wxE1ccR3aWUj9LughzyLJnbZMz+Jay88DcbHqN0gMuUxCNGVgiEPa6jgfS8hja
x3BYcMyCsBnodOIbTDzcZ7prpYw74fwaMIScCChwNhinYcV94Py42Sk1CpC6f58jvCk1+PUAMYF5
QDfNqW1Y0Fd/d7rvKVQZp6614Gnpaj+hBji/eKQU9cuV8/BrPNp4cd4NY0vLc2U3iLhaSSgQ0JF9
EmLxG2G9sUPFxAQb9nxm9JJGWOKrVxRPgfN+vNS+v9NRICxshxF0E+g+0grqdoXETKGyehZder2q
otPvlTPhoMOVADNXAo8d6qJ9zxml7LuU/E8hM4iYZo8n9fZjFf5ovKWu8/9gCTEpvFohj7+DDhvQ
GwnJKUOSiOERh7bI0JKOcR/2KqUjlp92ZysJE29WnKWN7hNhKOOtNfEDcBH42cq/K4OTP1BrMauP
YAmUiBjpDWbsR8lteQTGLdGHURBAdqbgHRDACj9+PchmV7Kx09m4t2mRdo4js+vnKFqwCTBqM5LU
JAffeWcJ4CC3JRqXqEiLeKqN065oZU2A53+FNNOXVxpvrngTC5mM4TksjezFc54qsBY19MpwdRS8
LAhrsRhmFSIc3sWQaYuTE1chHPR/QR1cgohyzDuM707cqEbtrBaSlYiRU3Q+34xgJXo96k7Af9s6
VPRaaug+mRRkMz6ZO1BR6HVBJQBhcFkom1OkvoXXsW1xdw4gWhQaCLO49UVvuf+HZuSQt1fxmhlS
9z0lLZUbXT6r+EV84WJsltyhVY9SY9N74uMmpuJVG+n7GLHKHAfT6PO/V2yYolywfYza+7F8r42f
Lqt4uW63SQCBqNLyZSVQDf8tW8Eh8HfRkTXVFjNXh8xqBcNYBmYTmKxrHN6KPdAf9XkzVOU9dy4r
sGsPCZRCTiBwxDsQJwUu+ZCnw4nVLU5Kz9KXJYua0syK3tmbRrLpohPLpIDadOPs57LyIypuxhyz
K7GtjyPmOzxOXmd0A3OHwHhWYETSJAjgkMIG0IzsgiPpVKKY7TiNTgoXs+Y7ASbBiDb46z4dY3C0
Ol+Sep7ZZeDIIdPX6w3sVIokzXXwgFHCjM6AiKU0PfqXK2fhSa2FvuektvmVl9d7IOqYgcetRdEL
3SXpaiZEmhxPmEGSMHwYGbqcYMVmsWIgDLkG9eNhXFSIHChV/Qr+ugixQSOyJmV7vXznDr9fZj7E
LbSZBrue+oID6/Tpqha3T96eLZ6VjL6XGg+J8zoXjzMWUKvphkD8JG57XlgAo066Ho3OS/8dbAyu
ak8FgS3GaCjobUu0f1udSb4P2XJ0b0Wk73RQAfwKomwCJNZO7jxHD8TZfsVSGWas3wF32bSv/Skr
3SR73jnnxeRnuAt19SnCgs7IHZlVKRUtW8GQaVoWSW2I23/GL7yJk0fHNsKPXZfWfqkEoO1JcgmM
nNMM8vVUXx7EYCLDjWzdK8Rwoz5dDNE/dv81XzVQ9u4K7KLa2l+AuPTQzWkMo34aoMlTPxq0h187
qf9lRxiod4xIo4wl6Oiu5jFfIcvtpPlGe3qSp/mcHyTCyCNoKSsytksEkeRObQlaFvACjkTYQUpb
G9HdzYGbzDpadL93Ealvl7Kq0xvP5WDhwYq+isggvIzlki7iRqI5idw/f1wsSUh5nUnaJ7i7fv0C
+p9ArYMCX/U6fZ3ET8CHtJlR5ZLDwdUVagY2ornFsbu94NYi8o5XpR5EQIuexQyX2q4Tge3YgOtW
b63nAfrKERA9SGOSUuR1BLR3VwgixQG5xfJ3aa7nA3Tplo/yDJHtwkLoPKA82I8zbi+/pFRbz3wL
x3hfanajE6CnCVPYe3+Yikfyp40C8/Np6ssJox6m5ENflhOXvHxLsZciU+dI8NURMPBtp7rXuCWT
ORCk7slZj4Mlruarn+y/X5No8aLNfPKcd4AtNvHbWnjb5KRi7xeip6hCe5iKiH6THZTrqV6zJ71l
nFN1p/nLvh6A6JACrl3sw658iVBPA9Dguap0Xhhx0rV9Eic1PiOn2YPp2W3wq9E1AqWWkVOdB9L1
jU/6jYqSmKj7P6Mm5P6jwuFDXsDu+1KJx/QoFfIAMKuxHpSKH6SNObUhGk9E4pqDOPAxKb4zNkUO
p/7Yf3VP9ydFLh8Ir8AOJRWkVDUZvEj1Sve1y2aoSYF4R95knoo1Uiw6XaczysmShFyV5B9y4Oc/
MzhbG/rHbg3gV79vviWxqMZa7f7npU54yL49gtIeGDQPWDwoNF1a6Az+Tl777uYhkFlMKNMCqs1/
T9ay9fedBmSp19wcGKXUEM16t878Lc/TCilnzPahb5yzxBKZHM9+yT56QLXT42ti8VRZxUVGqtaQ
VeF+4YZeAy2nxVe5Mfjej86SIcLm7lFmAz1aUsTK4yCj7YqNvFFN5+TKYNVXrm3/YtX7kcEQvsxk
79Pfp6lDpaubw+YJdjGoRY9LkIyBZOyc9fe95K6e+HlaubkAD9Kid9ir4IjkKm6RUUfu1xXfyUjb
9fEKdCiN5DUBIERmkuynUwNATwdmTWd5JH839opLQLx7wC0alrX5KzgM1aVBjTzQEZ5yTDjNEzqP
eW+3YDew/zpINW4K57WJeF7QPDhM6javVYOIootSdLDjAO18w37q+do+sFjCoIvMbw20Y7oBMZeC
zN4aZci7lfSCtt0kv7c7k4ig9BqTqOwJ25doI1mKXAd+5IrNm8YpGnZcFWOm/YPsvTsaASVO0io9
sZTZMH62zUDp+0+OJqr8XdI4SxhNBLbXZ5qbcqswDj3qAcWC9fXw1xzSzy+oStiKBfgRoCM3ZSOb
XQ+7KGMv4YEmmpU92fh573FceHQB4EWC7ZaimaOIxxCJ95sV+M+sP7hDiyTlzQeOr5QC0pd9sCCy
bIS0GGWpDt5ZIkkMDf70ktVyfpQC9D3bw6hM10IMpVC4XdXYU5qI125zR41tfcF6L9qn3MPIo0im
4TknBJhpQA/l6AJcWaoEsQMYFgHmYRXpA4b/ashJuAHj6KGS9tWD13G0FLshQ7pPcU1Nlt5kj6/G
EFdGdBBv8TrlBHch1c1LD329bTE06oNLpfj0ag1oIMG58YmNS77QImxtEWlKiqj/q0791umnOFci
HUeKbjymaZcWuVtPERFufpnAWH3QXteZbZFz9okYLf9bxY+VdDfk6h1PZcmM7kiPhgRyFICJ9/Z3
oH3GvaOcGU5I72GrYt5GAnm8Mkg2pmVYcVidPPQKeJVGNi76S9aF4XTHoXkhOV6eL4UW5JaHmJxL
dzBalYEZzBBogNnDplRaGzjXjZkzONLIy+Dsp5c5AIXfdSXZr0TczPe0Fi97slfOvJKi1+h6fXO4
g0Ucmau1Vylyik3rBTLvd9wKSWv4gFSlfrUXFBNujZqotE68U8Mxc9KrH+nxX1YZCfYMS83CkE6v
qepKxdLAN3az6xMZBSuLZR2ZDimQO5TzkVDRAh1qcVDWuSw3uIcdiHMI4yaWbhGu3RnSH9LVSs4j
EpzJml4KfObhkvcM2F6+CywPw4VfkWnwOYUYPjZbI4UEdiVvRyGvzfcIpW21/ipI8Uxr9/GdXlwo
/VwvXYTr+6yw9FrSmmVGlXYb+86svcYY60ggrfngk7aa5KqqmtrQFY8dXAs19ge4BZuEbL0SOZK8
EAwoc2OC4AdZvPuGg9qyf0GiXhGhv6md4+chndFHb8VeqWQI8zrXdzb5UvPOmCM81ZMuP6GtYPwH
rW2QnhKJDGEivGp2QrAsIqPStmbDcY95aWG8U7udTd4xvTZCruWUO1J4DzcHT6OIpC53jokwrhbZ
uQX6jcAr8xk7N0u//zTcLwN+OqkfGQclNdF2YmMKLTjPbd6hUm9YNOL9oGKtqaN4XKmKMlpSDeR1
XsecL/WoOmacDf2PwC1G7kzOtfhpCkEeOE8M4MJ7q4xIEhQKih01eal9y9OaWCt3CgNmHoGeoWMY
oi/xCd8rrXNwAsgik+k6nkEnvIYZEb8WLRpANvD/Efe6C1kNp1XrXGwoDxM/uST2cIkrktsDfUuI
dJV871EK5jB6COK7XwSf1BICxFdei7+a7KyZLXb5ULcX4bhlvYm998wwfv5sFUH5DxRhFF243DLT
09BvXmtoBwMP6xcmVhyoZTfd4E1v6c25yhGlYAYBL5XsSTDH10KuKdStUnQe0CA71Hm2Uxokey+d
vPAGvJxwi8ytK7hIA7p9AvL9o9bAvno/kgEXomScD7LWa/skaFXRH8YNnMYn/X1r5KMx7sZ13GII
98a/L9ldD+K5FVuwSHz8l9hu7x7In5JlSqsielH0MPO9QfXbKId9UkY3cIxZlauU7/MvCiYPOTXJ
Ne7qWHsl1ihOdeYmo6g7CV+RYHtcJR/pbs5kg8XJgjpkDUilZxAWL/9L8wWGveisSEy91J3zdSMj
i3G+Y/t+FmrgVVtukhL6gaGNw+qLPwM1aYotCM3kedreEIYbl4AuPqYTceOmZPxOZuoFkmMoqUpK
GpJikykDZZhl4cFlrqHHcbHnke4ZoYy43z2dTiU8qnFg5aAyWQdfF1SO4Cz61KkH21KxVHLULJtj
Ua77qiXlc1G4hhZK7sZdgRvGdCNEVamRp1MzbrlDRT6JZgsd3pcPPn8ek28dNeEvEMrrk8rodjO2
rSly53mQLzj8ePTCDb2oxQtQKaS9qfbPzkfpbXVAT6dLAgxiT6ATD6fyMni2X8Llp1/1LWursNb7
2G2hqN+M5NW0GGkqVoTdURnrHCZGCkI08GuC4ZiSRvvzw7EDiA8DML6q2NYmcsOFu0ALTmoL2fig
klZJ5E/fcp9mIBZgNrQScPcBSylAgC50yUPZaJQbhzT+UwEMZjCz2Lxl+P1k/SIi80Zsu1IfoYnf
/sMmRujKLsz8DGRhuR8KrvGH3bBVl8SGHlKGED9VrfnzNE4WDirdgrTWc/wgn6rpFr8fn2vGruvl
NnUxKQGUnB5i7TS7c6C9aRPZer96cZPvEr6yC5KFtR3CXn54Nl3Xo7h+QVpYldu1RVzPOHAnz3rr
wXTJzfdXncJgknpLdlXa8ytaI9sskc488gDI1cO+lrQu5ruyN6SfucrLhR6DM4Yie4mzBE9edtGV
qbLRn/5V65MlVTxl/vLSfReoU4jUwgycOelIl+8F4Xymby30PYiqh+aEc2e9qOFontxXUiHl6/Xy
0G9qop2ek/bvGsBHjDSZE2lFiYdy3gZyB6bwyJXE239oGIhaf+K0UPe9H+rQalX5Uh5evc+IK4J0
B7zetLuCu11kr8ULbqoTID8LMmI6E7pbiklwN+cO7p2KDyFBdrkb7UMvRHsd3z7g/MBxcpebUtTt
/UHLGds7b4CjLCst4TR/vzPOkRg1bILg+HmZ4u3khEJbXo7AuIz07uQNLmLs+xcfnJkTY9TAN88e
Sf6rI8vgVgfxXsrSfxNuWed9/bF3qdGGUZkxv0zRPdcSNqGobSFG1wnpwWOk6VyO74phB85j7g8G
DoNGHFElehpd8Rh+gLiEFj0b6NAuEY287O3DEqrmI3tD+rzPLkOI63Ukn3dQY86jRL2fOJX6S2mX
kH5jv8UDBdHkhdb5AaNyQVfW5fxEZl7eB48SNnDf3YIpbd9Q+5ty3vEPaekS8e8g3UY5K52yB/SZ
iuUh7BYWymt1BNBRAu/2jUowrXZSgzzCYP2xQ81uyI6kSJB8ID662plkbywZ25h28mqoGQ81ifNh
tL0F//3Rx2YB08DEqDDIBlKAaqfuEoU66bB8wK61hvIzaf+Sf8uGBSv39IcsJyvSDng1+jSTvGic
NTLg1QG6wVNQvmBh5DhBQPWW5dt0SDpYFq3G08O06e4duuE2LhAki47LmQW9BBWtxNQ4cBYJ1rVh
hLjtNkFEuAh3TRx5Dv+C3Vbsev2xXN7rWg6ykfoI3iW4i5jnbCCOv5tgVw3NsY8pr/X9EAD4KS49
pG6sZ803ts6rwOgCAcAhUuTPf1n8JQOeJwT8C+/pb6Rn9c7/g/M2tWMc9I+ce+qm8LwdBmaGQscu
XEvtqgirJF9rIhlxPFapfkucGZSf/fNTD93vtKlMfsMEkF38cd23VExG0D+ZZDco4FYjfBMCf0h+
xvM3ekN3BXXfPzSITojGkY2ZaLIOxXRjYPVzzx9f77TWXJ23WCFzlghh+IJk4vqr+v9tGms+pW7e
vXyGqDo6GYImGyHFvdlj7pd1q1i2roTnhEVVtx167KWYTJB9K+s7WMJp4YwlNCRQVCy00GXhZe4H
hJmLvvqJQLGHLkxP/w0OHWbgwLzXW2KCciEGvmIIxru0I+VIKbG6mOzc7qhYlaVYsBefy69cZaF5
Lt3uz4l0DMH+gi+DnqrL2XMBXzahvRvKZQHcuUFgTU8hkhLe+umVzZvfqq1NK0uGoQrRI4AdXjLT
DvfGw4DSvXHnu107RqFkfvrGpNpCWYgr/AQcZkJiYF0ZdujWkhpJNhXPwBSQpshUTQYcygM3miYQ
q4QMpn7CzfoAbS6cl1Mp4kA9OECbm0uhgO1Uk/L5osMcUaFJYjHKASzFsRZdLHXvZLoXbl480sxB
65Uh4oyTZamI61I36JmoHgEpGo3wefVsUgFyLl8lbnlRgDHpPsT93oi5O2P/DvFbKIgtV8ATq7l/
rVsB/rrrfQIp7JMw8Ri7XHLBzfU0MZH7r+YW3VLzvmFfaAiZjp2EO9WAjXJbptmFYjEpbfeMQlBj
DFvkey1OfcFVMKvr+h4VJWmn5bhEkL39VuVDB0VYEcJFpoNrRvomcxOm/umBFKu9oVriLwATTsFH
h3K5ySj6qu74zhm8VQf3kk3ICNv94Y4N9pd/rpoRwk54H7KVGmjtdA3m3/ls9LmscK5bVDXMVgvT
3IY6mSq12s/SJ8pcOn11e84t/OmDjqwzqIGjVGCtx5Oe8FJd8ugOvKEi582DBFzo5HqZKC+jlMD5
3NgbYOU+dQiJ60PO4XOnqw51v3uVSBA3Zu1T5q1OHQ/AHV+Xvfb8FEq/Hch7nZKV4jN+CWbLwEx3
T3Zj15nyFIHrN93yijuf7kBgBjxZv23Q+5xPrWj4LOoB+7Ya7hmYQ1k0Q/4WDz81Uisl3QgcvXYT
Zo6ooM6shsCCZ58/69ZlY+9Yor3dnSBWzJVDG13x2dA6o6N1Y/2jr3maI+ZdTGfO8km6e01CCAuL
PfD4l6jQPtebYkxQxbXMbma0dCAynzs4+Zw2+CUirVMnd7H823Ir7XGWJbjQwojtEGgzEkK2kj+o
ryonxUMOcg4gCoL+bPh0OGcBhc0Z95p5oCUxgm1Xx/Xpcsk/FxQRLM3XZ6l7Q4K/1QRa8SHZoR3b
PnvKPpl2fPVk0NXJJX0kaL9Lsel4WxPBXJJr0HUVOYJKv/CpqE5PqNefAZV78AbFk2v33k0nYjky
88dZlYr0+4BH+0JdfpeE3CgfjvwscSLOuAXVZ980FhdHSWlhkpy7NybzV6AOTK/Cz0oX9f39zVSg
BKD5bSSb+bb/U1q3VMzHnGy3Fn2ii0kVYdUKjPHepwzYD4ViE8MA4PnYrtfzqg1YX6/WHKTPc3kr
qUTTxDcPkxotlyde9+FYRRqMSc6hap0T0CDxp40luBan3YDl51GB6yYVGcW8Fd4FExIH6+DakrOI
dGFm8pzrThlq9lqGAglD7kYGlX4pbtvUvUXJqHWGr5BfqMEsR/R3PDqs5mlnGHz5WTTkyX1XVtBX
NA6EF9/SrsdhJdRQna+H82ugvUEclfYM6z5+BD8dHRdTkE2cQyHsrulVFgX7sdxMHz1fpSOW3FgM
jgoY2GmsZ6zx1QU5dhk+lvXRLACrwDRtMj8HaggzRKiq1L9IIhaacXMSYPCg2hxiom6U2/pDzuVP
cmCabUopjBIehwV8m3+ltWvDdV13dqOXtMRlGwMsg6mmcD8kfLnoto2plML360HxicY4yV/945mA
RW5nOR/vRUFLE9WQn7YHsfxZdoTIhEMC0mN52MCYQeG8mkaIG2nRDy9YCqZQK40dhX9xS7YUYasI
6kkLyRANfRNvKRioYuHQhYpdDGkTUmFKxHKX21MvGme+xQ2ZYYRsd3LR7HdhJs0xkAznoikk/UVx
CWVUlE1+5Lix8EPYIY2ZkmlNbM9HvRhJmOVeF/8OtMR+toe7Y2nzGbju5uZfYdmvPn7UYSB+h80U
S9s4AM04nBfGFei4DvSP9rf8M4oJQhjA0x7zx0bkIAhDjd91sIB2vR3zJNVtbaRSkSl6CccqHlKK
YENdInpZVZCpQrswSpcFUBxfCLvQSjpJ0cTt7VQY6zUpIFwtj8GTHLk74r/dbK1qLDf5BzggJmqv
Un+M0/HKucYea0yI14ugN1ry47qPMPZUuL1u+tZdEjoMxb/b1RGlybx4/MclRlGofiaibOcbIq2F
/XsLY7UhYZ7ny994chQP/7Z+ZbF229RJV/do8zVgM7TYtSBguIxn8tEljxhBRTUoU4TvxeNt+y0t
kHJnwUFvFvY4G5YLQKeanN1gLFdrfahCouO5K9jpfmI8TKfZ0D0YUPDcAfNsHWBlAqVmiaketT2n
7k3ILdmGLTiNUPeMbtiJ8k/bQnqy7wbThw6swlsy0GB2xg1/84YVzRKuIBKSTeGKy0L93gNmmb32
WMlfF/hv8uq6+x8YDxMZaA2+ymwsA7dlhb9sBlX2vQ2Ni4eOQNET9Pnelgk/rwu8ca+sxatoy2dV
gx7w6OHd43bHPB8nAw8hUXJ/5QzWTmEce6q3t9rbOhEI+AHvteL5pExorpepDIdkFzz8Rt+E7+W4
GDEvYjMDaVCfmulVzsvwUWAX11gUETEx1a9Ify+z8NmrnYJiU+utyE0bFHK26cfxCvFJojW8HbNM
IILzXKX798910H558HIjmF2q0NolHWqgE09Iw6AAqsj3YF2NfneY1lKYqp9h4TYDqLkYeNmrRClL
vG/W/Y3NI+4xnbd46O+DPf6Oi35CJ6C2sg/IpkR8e2sU1raXGfaLIniSK24V9mU8MZsmOXxDxpLE
1FPRLQrMTs8enP/PiWiXCElCI7zsuPvXAC0q7J8vkEW8b8wcpMZu7z5yZu4JGpRlNtPoEiU+mecn
Dnl4CtQT4T3E2DbqIo/d3rCOTWV/NXNd5+99cvLhwHKicUUlO5v03LAFdHPZ36xLK9vGadjJRvA8
yZd/wb5NIFV9kkKitohSY1iUNCwvPBzIf7OXD8goUcpvWv0IG3ybRAo4NjrgzswpSCpdzHJSDPiE
RR5bYYJ0PLadewlvVpPnEOajpXKWGzUo4eaffKB/F+4cg3EtmVDC9dIIn/gUrqscaAzMk+QR3nGR
vQnul/vg8vRRDgqD3TloI8wdTgtrhc2tBeRipbHo/SNqfU1Hxe6o0Vs1Iz7Qjq9aNSO8vzhA9wP2
0ErGUFroqkg8JpOJk1HpHC30jcat1NoNPRviweXeFyutVTB7R+TgjVHz5Vs2ic/VJxXzyE5dkWns
xBKBCPOigbbOA871o7+hkpKPEyC5V5zapiG7+Awo2YiPlhMFFDu34TglQ8j0WUPbQiMR+Q5QuTGU
N16R0hy4Qm1BPt0sOhrokNh0gUKQAvwr25L42c8MlVe1tuJPJWfyzz7+Dj6Nn2EksWlPEpliFthF
6ZX2H7VllBcI0FuZN4R5Z+M7Uk4eNvIz7K41sCa+SbEVyK2pCwFxfgPBaSSU5vj/ol/8nm6eRqX5
mXgPB7DzACEn6og5MYPgajRkp+dkjVDqiJ9aL27oHWkkTU22UrG0poX8rGp879/XzYgDxL/mtlqb
l6Kar7RJ/Z4iB4/KvTcGg4de3HfTBSAhbbuRxLwtpW4WKnFcxpb3UfkJ6uSwKwMgbPedWq3TOFcc
/8VTHswz29b27BSCDJM0e5hgU4nLHVxBvJtrm2gJpetKt3VC4igy4w/jf9oN50KEl/iMOYLHFFfr
IuPG85pMO1rLu1kk48zy1C5s0cITMrmPeUd5MN0yUucIHhM8hytu2vLCvj3UXaNrNnhh76v4IcjD
EpXMc7EYA0R2PacypxIPe/HzZLBx60H8o4MC1yh8audbjVXYJKvQ7UiD+/ONZdE2JvVfEDFIdRNH
T7EY98n+qYgcPCpE5cZZE/+BP5wG35tcsk0F+iz5nvLSJzXjWHAKOJoSPbqf9vwvO0shUe8GhCIj
XQEjwK0ir6n7s6L5vkKSY4Z7Z9uw18YhtsGQ8bTeECwBTZu7ca+zMCr7wQ1tTMHcFyyojVBM92kg
LsZktSNqtaBEQT1CjToDq52Q5T3IXZqW261sLVSNDZ6lj9ykyjxA8bRsbgKGDpV1I3p/BiYAahkW
YJ6OZsRsY5pdWeeglvb1Q0ldxIBCOrLz9BRjTKDVroKe6pI/4RLKtRY4JRQLygfmAnKdbjZq0il4
rRTG7EKruFxW5yZCOyHJoFDgbDeupH+RpJ9JdBDTjx29JPOQlSD3l+nS9CAiIRNwoGQbhhp0VIYz
LIuZ/FVIUKU2SlYT2lOCqG5w42F1+vUP71AQ7mg+4qafPod/Fg7JyezdwPN+9fxYIhRoC8+FhR9t
Yy7dCC1VqI+LMod72tBhktEE9reDvilwQdVbRBCg1+B0k5j1d2O2YIT3AG+DERcyuVHVwtDwAC6Y
jXoweyBWO25x8XABVA+kqdQZVFH+opY7TFUKgqLHSfUVuX8EeRxPvrLtESaA4gtfcIL5yN4g1MKy
+Wn3GXA+B7qS8zaBynrUoHDqngRRhwoDbRwN/yAfOIHRZaWd8bxf3CZn677e140EM1ie70fP+Sze
XYQXcWT7wSWEHeaHfGmHdqE1C2yYyq+l+YMq2mPHwZvQtL8PjF4JgIWHnzxxsJLd8+lrWRf+dify
KDjWRTam6HfomPgGMtcEj+JeOjoHuEpPBj+svCBziOfN/v+Gv/GAzm1lL8MGE3ccN9VhW+JnPhPH
wDtWyRBesWrioWVOsI/u9xfrVVncDxDpt6ZtZUvceb2x2pl8ykOBeKWdKMuUZmRPMeXGXaI1FowG
ZCJiBYiJTHRQGe7WpdAaTl+okEDvWcUsFMkGRjhgDuaL14QA/tHwhGonSbCkZbbeW9XOzJT7wvdN
0SxU55cvLv310jVQsKLAzcm6gZ3GRseexqIi0CkAON7895fp877kNN+OJVOuR8lKJThDZ5nlTUAL
XQtT7d1nTmZmTB0CYYnK7CTsKbCvCsvGJZ/YidVZgGnVUdj65bH6A0yTaNzp2v+cTnkcdz7aXTg7
PpuB+azu2QPzw8NgwRj2Br23KLX8LQ/OYxfJv7Q+1ObDG5Ku5HXbNQgsBXSJrqmbj1wwc6OQ8ppD
GAtXHLVED3jF5V+pSGPTxhRujGcjHQHf93QKOfqoR62G+4vr3MHDs5j8WtB1u9hxf7RbP8rDw0pL
4fcXLTwH9CA8ERhfxd/yxrsCLHcctfKdyt/1scCCcBmySuvOXgtmm0/wK7QxfvT9rVI0oyAMXrjX
RKHAgn+MP8ciEoMgUprB8P+Lgl8KT6n9WzceKP7F6QVJjAJNq+b6ltWOhzaPvxboVIqTD5Ptn2FW
G/fbN83gpxipiv9Rq4Iuf41xIBOJxe3RMj0MnvoDHAYUqys4H8rmWcULl11+wye7M8QyShZFGDBT
yWlD8LkgYHVVFOurbONiwGo10kAdWW10XtJfsG5QPsfb/izlTxiEKiWd57z98TG2h+oos6QS3N2C
aGI6XtyWVxLAZuLU3LG6khtgrbPrQNe8ZkhYHXwf1HlCjEIRXwnHlfi2kNyrDm6YpuR8HWBVY8MZ
Fcn8RRVIsxhKAWB28QSBvO/Rl+xG2MLoKuv+f0UVOm/wvxJcuOae93eXyO3uf5PTQK+ZT2nXp1r5
KLqaIy1B9yM8bCg7qeol8LS8eeg1DiX/JhKTn0Kg570fBQqGpwcVQL8mWs2ZIDqaZtPwfPsIw99/
AiFXEQEtob38atm5zHI5LfvwEiA2wMUzDhzukxA57lpH7vYHJmhnA7/YSfETFyQBoWt5IdAGsJlB
uTuoTkBnVPWuY1ixQZjOZ4NOnIv5SuU9wK1s9O82Mu8BloX0Ncd7PD2rm37lz0equ3z/ebaPt+i7
v/oGECk92hPKihDLydzUtkGKYj3gC/rIwDq9H0wnr09EhJwke1McbdzT5BpxbOBrypSMnhVTEUcY
yvd8FxNl242SLduql191jDCGsvy8NC2iv9ro/iDN1XMM/Co0L0eWZW2ol5yem2GycK3RQ5ro8kNT
58NpQppNH7lJYp42/Wp5GJSRIS1exuXgZHkw3jT7GxoreIrakXKbkFO1zftAq3nHYaTMjFIBxl1k
GLLzamKaeu+ZPYSMIO+2I7DCKYzqZQZFviuM0GJnmXagtN/5M045IKhpK7nGrgMKQW7g7mbGmPwj
mY1DxWAP+Ah6LwZwqoLUybPOsFYXk0z9a1Zy/shFFNPpuVSAWCWiJtXZNmC7SoJ+MItoqE3SdSGl
1tyNnVT0kIAbYvWeqeEM2bqNJfod6H6fM/5DW2Ke6VIGMtJfqunGKdUJ6URLN+5xVwzEyOPDVDBt
51R2DJgHmq1bpQzCDMQoL+smDE3Z52+qqiIG3RjAZguJYy+i1wOBY+oBdSPEIPw+T4mRkkQkw3YQ
kLLjfmzJtUa06KZDyPVang5ht0NFpa3374fs1LIiAAsiRRGWuyR/WTqiwA8jzf61/uYo1q2INTCr
rRRjKuWkaQtMGHVFPTll7H2owcEVM/Mq3GM5XBN6XJ6KbkJseJk3LYuw05vULInPyQy8lPc3NJBK
OKxKUP2KxiP1ENscGST0iKydVCt5/JGG3jwtP4uMYaYpY90A8gtbXt7F/xLuDVASXQU7k2bjP/i6
m30YnIV3QFTiDdibU6Muv1U9/tV48PEGhv5xcluiZ90eh/bNY4Tnpq82RU4MLdtKUM8AelBr1G3W
uKWrnfnkMyx1TjElp0tYVyRfqs2owf3W24vkL+4AZgr9j8p+LutToK7/mbLnVKOiSDNvfTXEesCU
lA3ijl2Ak0mJHz1R2nadl6iywsYHAKWtNZBxckGWq4eye1gzkGf0r3TetJFsHebpUqYCeuzzAMrR
kcpoQXXno3Ffz19XIBv+k8vUmLo85zkMGckeiDgOrxJAADe6OopXQQX8wHR2mhrF3AnM/vdTs41/
nzew3p7Jxd1c8SMzwbunlVC56Ur303ezddUY9aq5otjwlZFYSFmyhMbDdjQhPpvTHxGGP4yxuaGG
mXkE8VMrdE2EKByDnH8iUY5zsKJKJ2F/xDDiJF04jYR5qthTRlPqExZGHHOzl7RHBIAEV0CqSrHm
/SIciSONWO3s0VnW5pSbq1U5BUybhxvzt8WLXM1LVBPBjkZVh/mWML7lTc+PTEXV9eVYIDfwvjmK
viTbEP58f0r3NzeP/XjB46O1yxhk4znano/7Bahzw44L+oBKbsZ93B2T4SoEtphbpzC8pGf1PvhD
Gl0ZpG23P4XY+ZltDsDHU1JAsDgSpsIYVN7RfxmumxQj2/jMvFF9AUFqkn5c51MINSjlgWGlo6ym
g7AZ7wvTUx8DKY0Re59g9lyDpjhKe/asBCXod1yh05b7fpLou0/vTFX/vcCrAxo+jBORYwMo85sp
pMof93VLBJHnLLRBRvmbJQ/ffUoEiTgW+uZlMMeNivfXnu3fwcmmMjedvFxNH+EqjKWG9FwyllVW
5trMJp1X7tkRFCvPnvxGoZKGpBTAZMs62ZV9reZPF5q3igB2aq2K+tTY43BfIbcw/xw3YnbbiJeM
raCDLUDQqspYzovEpFkBASRRmILN31IeTauK4q6BzNHicKGFpx6Lxa/3WB7eLaffe+LPnGGDxxkH
xxm7iwEg8Sqx9IFsRsgbicmjgUnVmztqFM76RV0M59Ulw6bZQLytGOTXJMujOBJ8PBzCbgvdf4hU
rA4qh8vIAxzpyZiWXLmpS9eNl7SpgQbLt3K4Cd+NbjwViTjnfbJkbQnUJyV63vI/868kRyrsxuTT
ybg74YguOEhvpPlRFsQ1R0OFlBwOOlT0YaExHbIvnt0/JtjY6OYRFJZX9ATpaquMRWnf+PtnVmiO
nhc34XPkLvMqdo3B+fiJI8UMs99lO4xt1Ffan+SHFdF/eMQ3dubWtM8noNmYNyHtvfJrMO+uO8qa
jxEmqG7y9k3ecAQxVtgoqPHKYgLsbSS1rzgxL9mjqjDzh+oUvixxEjIIgkgFtQmNtVVKn9Dmsh25
YGki9R5Ud3kf6m3rAtU5ludbVS3gQxVhOouDTUtgemrKsw/REZ72qm0YAxeGSdwuKS/WVqTNubU5
cTfzgz2fhhvS6ljwbgnT4lZB3+bXEIhpZExo+mE2WtVbl+OgK19ehJB6QcpYmOfKl94aC1nYIqJ+
zYSfgrd0+bNgArGW8w4YZxibE5SW4IOPPUAep1LhGj0+2JCBzpwpFR/xTUe7BXV28pDj/94kV0Pd
shsUpTQbn4897c6NmV440lTFBrVJO6UqSXLKAXslZGEmUBaWsu665Yw6NhaXtkaHmqOhzFCim9vn
u4yy55GlhtPIZ4IoQYRbMoYGsyWBfz2qyM2N3ql68Monq3ljb+FXV/kW32R+HcbDz77iPc8Hn9s7
IeH3GbdDrOE/goDZWQ+oKDlbyFs19r4KVlpngqfvS1HKDVUlCwj8F61F2UQr8EUsQO3kqeZxbM5i
qC+MpPcU42KEF54fUOmk5qoEEKqLutFyJXHXVZ9kCtj+Km4hdrCRIoFYZkUV3PlgyMl1yHJcmCDj
CfGmztbozvEmmwLITlcFzcVkxEffSwDLS0f5qqDNjH9maKrti4hk3vl1BdjB+nnDhrh4KkVxHGWg
1/px3wOuabVvSiSmKtBteXC0ncOkgeZA/nFGOm8jbupcjWp2Bn2ZvcxfT4VWRAu1VNrHopWhPugP
BQv1Pb76Z0pU48zSdY2AcnRyYjwqcP5M7yhrCl16COEJeNyXpXr/Dz1ohSqeQ/1C5B3OD11QqtxS
kZ3vmNqHkVxrYRkOJoGkE7gg1qR7nMVrCKFNfZzZbYCj4lz5e54Xc9/GWSSoJL+yWeAj0+KQV5BF
sQfcw2Zv86SlkKzakYQb1mlmNzSZbfhYiV0RTmYsXtVnhjPSfDqmcZBojPkfU/+olRhkww9dYNJu
GuZ1FyQG1lWG3XW79g7yh4VSPKp0ycpyldoSTqCKhA1yZU5PDEzEfoRpeL3okvWeC15/T76n0FtY
XAAnZ+Lm1FrEMiUeA2NdMYuV8fZHHwWUwcX0loiO0ulf/J7PO+S9WnOd4lLwp2ZAb/qco1c7rPsL
7a8sBpTyyD8hkXbHaU6HaRpIWTgv/zmgetN13F2dcVCTWnSS8ajnQnXt+woV4sWVDkVkn/grTfaK
63nO6Ujn76mNilBPnEXZzFYt4QDjce38jRWS2KJFWBxkanvIBmMamwz+0yPJynM2xIQjKIfLt00e
mUmt1Bw4ngaHJNleK5JG5RzB6SJ8rmdHON+1zKnkkCD8olRWRCWsIb5IaSYbLRiHy4pDZiheD4XO
XXtEr+ugXl/Udp2Rk7HNuSeMdMZtQ7yDiKGILmfk6sXRdwNAr5YoDgyEpZQ+Th5v1vTWYo0300UW
CYDXes6ZbZBDN8PYPaCsZe4ySMIts/wIv+iNR02uszn13occTTuY22pxPvTFZq40aalivDv6BhxL
IH2DSKKNAuFejKgzEmA0sl7ULJJ7IfrTKsJWiJWE3ocfaRMMwEhh6pGF9i2vcAypAM6HkCNkLlhu
f0RZOUebG25RnDhOOqFwg/me3q15/v3X84b+ah/XbKGbYBP4C6FSn/KhFHt+QIIejQ7eVaZho2mu
TcHYnNFdJHRxszEbhzL80CuMMMKUrI/RCkR3xShgoSss/Qb0Ch4SoN6KoqRIilUA4sYAw6EqO9fO
2i/ooAc48z7VeUEiiucnye19i57j9MGPyHfpbd2Lc5jbLk9q+lp33/xvkKme3UTvjhz6+dlMSe5M
y/KaWjIwwogw2dNcL7zgdyER+/pceo0iB8r7+kY+O1ApJZakGm0Ct5SA36HTTP34E3uatCJdlQah
D9qYfChWwiwVqKO/cZH7tuKGsJio3NzYKtPFA3kf1psjipPXb8tymwqaXf/OYfqfw3KBMOkrNElR
IjUTIar0b/vvmxCGq9YZPskZamJJNktnsXVDuMibXN70pI8G41xZY7k2ud02IYS/tH64yDFtCD5+
YsKdkcRhNFuPUlgjrRHpRdMrn45yDQdKopxqnCDpGMs6wX+f/R5/3ocCetp3a7OawMeJbG8LvuGf
/TPlS2vh7e/4ivPOpN5YPX1OfFj1DPniEd2s2+tTdxAUoU6ocs4rG2RIxCxVqyo0wH5lWrKOoWXb
MtTwMV30ps3Kx4abJVbaPLWpYqWR3u+ouZhbAHc4SPLPGC+7gyBXbOv9+jeV5xuuJaO/hs5g9REQ
8mnD8kCH9GDz0SPRvX2Gzio4rDL1DsOq2A0pP07yCTdWlfyCPcjAr5radKweTtaVdBv3lkzA+JS3
5zqWg9CpPd0+05KkLU/zgU8wL3N/ftbK8NnCkkQRWvTqgN5bGrS2gs8VgWcMagn1QovC8svmdc5o
7q47IKeH8ziHccJGdXkNvVt1NnhBTuKxk3VFCb48bS+Ict0I2wWwYSiuiRaZbkYoONG9dmGJj3xs
Ph0BkE8mAo+0bRHKGQLpRBgXDMfHMlr7f0iUdJThVAu5ifj3lSiIc7Mo0i8qmp+/LhAk7u6rLUDB
hGiYosU3rtdloh4/nj6XGmT3F5i/OWfmTQKjGaX9BnJvrlKM1rtlHo39cM3bofK43RKYNYAayyCu
i6a3aAGVJR3OMc0xN6AnMre6zw5ygh5vheXuPuPl41zzizDVraSD131A+o/CGmDWvH0xpy4H5B02
koi0tkADsz+fQU/FTJoCXOj6fQpWkKXslso7L1hUnsMDtWWzCbQLv1vMnxZtu18fL4AbOgMz/x9o
PNxHzbLbXe0q//i+OMHKWN16/rYl66llL8VJF6k58aA4M0QDj9Jx6f7vXeeZFXS7aD5GoBK+fM71
CJGUMTB8DWbCP8C55pyTXL+e7GBJmMscdOrp1T4nN2/xE0tvaTFljpbtD8/VwoAY/wM0jUOkxMan
IuUdcwwEiDjCgtOjmx8kQfTrR3upnborJeMS5sbE6Z9fJi0leyeH3SReAxNeC54IanNaqg5GGsNm
4JgeeBh/Z1asBAvfoqH7136fc7JdLE3UBCYn9FHkJwkrTQh4oi0J55vLQKKi0xkUJuaCqgBYZjT8
19oawusXQRgMPKAH+SwOHDozqUccNtH508R5UHBe1hXwpj5ocxW3su2G6f/iNgZFqnVVg7Fn1pdY
j/tONVnBwPSKpD6EcJQ+8mXx/8IEeoA2vCWmKfXhM3MJsxRD4QrNmars8DjpmlXFu9BoOvdoxCSA
A8cdel15faaIyQCQst9qinAR2dk0esnY7LmK3WOYueRn1oQNz5E0ynwMl3HlXy99wej8Ajg9Rq/V
ZqqLPBll1XSmA+z1d1m2CubzvtgA0wjliPsIylo2P8EFssHYX7dR2zWO4dBC8BuQNNkpjXFzkM2Y
Y2uz5P92+7ZwsB1ErvWrgB/7Vgql6MtEi3pQlaq9sbAJrhZ9OoR+g1JX5oJXfXGnAsSGjcRgtaI4
EKNRSpMUgV8WdodQqKOvtJfHwzSHdw+AJqNVtcE1PLkrjb7FMkRRVcy4rp7zGHMbpe+UJ7XQasFX
v9jYTBLiuKHO/akE25xHp9I1V9ZC1uNwwugSPUsMpEnOdJjcjJoXO3BFu6KQMfWdpjwHaKSqTNg/
iNcaakfkT7Tl0VAbfHo3vg2glGVwUym2yUbgI5NE9BrTVAV1UDuU7AshKeCAAvz7FYOsQFmjPzm3
aFYkjOSIyFdTP01UYt0DmpgnvuFiGpkOfQqkgrfEZsvLf9OeOYgW0riyHHx+HGkt1Xc+e9Kyn2no
9IVt+8fWLhKNNAtMDOtPGX8ZUpUiWaDaYtmWfYzNLD6KWeTqYyBSRMRd80d6M0f3XszB0EIB2Emg
AAFIrYMK6cmIUXZWkXNSyQRWm5+AKCH89a+e/D8X5heVScoGNq9ACGgxHIHM7skgq0gswUWsGHgO
N4T81KRqUG/IWASqIZi5TBt31JJutbTtXOQ/tGEp28bZY9489d7gfjVgwppGW6J0V5AUGijn8GwX
MHACdO5UFjUJocrDMxfuLMQK5v3A0PgcKoWiliyuvH11EBrjyLsom/KqZx4X6r942mWJY/SvNukA
rjYkrt0EDPhvDJ9FvTjo9vRFZO/jIRECRIEBq0IW6R51o/GM48WyhHujvrDHTTvPX+7fKLiqBoVU
g/TncK91u+HoTg1QKWwN02+EOPbJYXhlcqmIPcVA7O0vF3GrWot6PQXw+fDhaRk/hNinqtNN3Qky
lvcNodAfv5lq9TY7dnSVOvEs5AfXQeV04aHRizITN2IyVa6d8p9/5LIF5TV9WAShBe8nQb2Fut7g
Bf2vrapVQraOJ+WKtN2KVSwBYYSaRP5tOMgAFRQxHrtmyV6+AXeVv7of41Fl8IeEKRZcYUgbybIG
gF6sB+MxMHxKk8a4nLnTyCxWYbSoKGGblmQ1o1J83jrH16O6MwOpvDsbCd5Pq+uwnJ9FinZlFa7R
6G/pNv16zJymRnO99ekSXT7KvW1Utq/D9DhLdLCTShIpqvmEBJIl9anszUBdPldkv6Qt/xiidzxt
U5w07GRj+/o0PriEzv30fN6Ssl7t8OA85Vo8OToZ4RkZpykG+4mSbXtwOdnccII7tySwvp7UneKr
SmOuWghKetoTvwGKNOiufjjTbN5FRwRjZpo9MzDH/MtCTH4+xOC475yENbJTVD28wzQQ6uiHXI+W
IzorPZ1gRkVE8g+4qho72Vlqj1B1NVxSFaE7HM/JvJacCwSKlT5BprJSsgGj1+4x5/EXJaqtA+Ml
LvEWklsKP/PkNkIOkREf8mPHJ5T9WKh/HAKMV9VqSnrCQj9sEP0h+huSvpRUnyziXb0z88ER8lqh
0InI9iC88nWIj9B5n8n6emmAN934b+SUnf1tbWQ9oFeRFIW897ImowA+8Av181KO+OCbjGmN1mH8
vp87/9Rh89YdEDonLpHIGLiLQO35IrtfAL7gsTx8kpKSBXDZcjVAcpOn0PYgSNXOY1w8MiurRwHh
rd+tGOKqEwf2V+9lTXn7YVyugIH7fM90ZFV83LzTAObbC29qvomhCy8Hirz00Tchr06lI5PbcN67
1UIBFuFQppSHJBrIxvANoRrJ8hybJ2FgSrCpS1i8anFhDm9R0G+j7Ji20aXssAF/162v7BG8iv7X
qrmWXxemPTE3NKy1sX1c3iLofqodVIeZ4fRSSbpmUKDqK+CYca1Ju285GNBKCzytSkurcVK2a0vT
UohPr51v2yQbzXdzYv8wxR/llu0nwqSnyNATsDkz2EqrsXANTU2hpZpVKIuDxs6Nmju0BqCfFDxE
/KWDu4bdVn7MdcdLN/mSUhfT79+bE2wZ+M1XJvt48vCgSUKb3pdk7OiN8abHl/vd1ywyl4HwNoKA
TmMI7Wb5mhR1iyQN8ZDJy/ZwYcxC46zYK4PaLCKZ7sRDbthzOQDIWRwEFB6h0axUxqk4k1kON2Yv
f7mIWUfhtLlplZvNZNMpWzlfE72ls3EOG9EVWIBs5EhIwZ0K8gHRoDvuEaLcz7zMbIRgZW1pfsAs
93wCarbn3ZVT2yAsENjnIqIVocRdkT7G8sLswBR7y4ERPdhSHdHol/KQx/BGrvy5RBRDwQRdiC8y
DNAFWGooRW2sGiq4OAspE7JaPbLyA61lpOu/KUZgWg7Ca9wXlTWk60EdwqRCIUp2V1M18QDJCHg6
RRlRo7rNAN7birXEVcl7P2Wj07osbcXJJaQjcOiIf67lV34xB5KEYcxxUqklwPQHVs7Q4/befa8+
mZy6Q2TPIHSxjdUVbxWdAJhGMvfApmwDXHIoptq4qEjRnxEMjI8IYF1ywIqYMg1i18QJkt1hFE5A
kXG0kVeAsy4WvqWI/oaxz7MM056rlK5Lb3L4pfeGVJUskJbOQN2X4EcnrlJvy02C6AzYLkbP/B0b
/D6mRANWENNkcD7HGD3yGyI3nOZ0u0RpOTrvK0z23e2VCIS0/Y8U9YHBVgHjikpRdg8obKMKyfoY
VR0/lw4X+lbXUFYSy5xeYlaScoofAcg2bPMCcVaPHhEb8dfoZ0RCaF+oH+KWSnoDjFsCRjR31SYQ
mUWrBuKm3JhFPsKMCZCyIejX+4DU+c1yf5pz31rTW7ToNkhurzSveTNGzUmQ8tAsspnYTXARryhF
IlUHi5XjakthRQ58z1bTVvZ8FZ+HRW6jVTMKX4iSLL00zI4GHvzZBLkmoeSJF92V+PpKRuDvrhKu
gCPUfWKS6yh8rr4rNqBG9asMOHRaildH6e6FabT5nJJWKv/6qWADdIMgaUQJOLq5sBfofdMnxZsZ
/hATHEj/4fM63EVvXLfWcsSKxzYyfbkkdEhG1jeXiz0BDzaCwMb+qnCV3IaJG7pRB58UNubBYotA
ZCsuqy8qYNp1TtPE+U/MNHmDxGzQcSL4p3hUYpEwWabT67ZZEN7koX/JoqQ8oEmGHLvXjYbn3RJV
hiFgRoyKI7780WfkchiZXhbO3PAyYB+0Wrp1lUkMfUE5jXkbAdiu9dpuFhCXK/HnKjMvp+BUTVSa
azD6ppXfwBOpd/+oiwVtymZB8vFQjOYphpD+qJsKRbnBxiSqgKkTLB5QlT5XDhx0jlujyLjTdvza
KhS2o/w8Fw3o7ZWnwWxs8fdEbtFQduoF7j26+kzP70RYvZrJ5W37l/4Kh+1h9rpE016M7WREjj+v
wOxoiJHnymbZqqCcREqe/ax/l5kZBMyGVS4GHXNnb4F263aTjlO0SsTfXjgWkTZoECMzC+woJPog
/Rz4/1IQcudkMvXqEfnvD/RctcCFng7q1tbLQaZqhFtmM2LnV5UB68+zTXR4bpTkNiyUX0Qua5RV
BnjWMtVRBOJ8Ft1SVSS5hS+jvyfWXTJMihj22rIt4bAqJsySEgaaOyzt4DGV41ySX2edLd/9G00u
EX0k7fLcik5dn3v6KCk/T5cIoJTaop60WJGN52kC02ogPx4ppa4MOqP7kBqFtaobcupp5gf4e0W9
Kmf+Yi3tnyEqEySe2Tk0/3EBtRsuZG5fUk/MvhYLuMuB55rXwbXXzNBWMO2OkJzD0sqDzXCZFNkt
bkzNKNKSpJIwNlqak3NkqWHp8Yb4FlIgAiV8HIVgYkZJt/uDZpP0mkwwRYgPuVbX2jdgXvyvZ7Uu
R7gkQU5WYSMcSBul/4+i10OKX/CTBzTbBDg34qOWsOhLOA+ZjWoSMx3qDIrFsaY60/F9wVq+v5m+
TGKoSf6SPmQhiIIJYVZHnCXp0Ya86pCwZWGlMics35ypjW6kSTuLuEKtYiTcTJW3xTjnmTbl/zPm
zVN4qCNiHkN8zeFa9tVMWV/jiGmRA7vNlmvaHwbb/G1/DCUOMI6QAqCjzkcbh52laHu23R7exMZQ
dDLqs2N2hrcJ8frGRWvO1XELFtT7cF/2uYfQH9iuMafryn6Ix0UMfF5xo07824yMp2DVtug8g+KZ
c5MiCWrcxkPItdUutef1APMPa+zyRnjkspdWXKs3+ns5ulQCxjsyOM2dJpRkmr8BN5bjZEQPhhJs
4S8BbKPcNh04hTHc3f8UQhlbqbeaQGnU+aS7XarGbx1gN4c+JNccASaLL5i37zlrdRvXcBL+IDyi
1T4MGzXmmSyC/DjqG5t7Gk9BXpUrB22ofGItNmg1SXC4KgCHS7ZkaI4z1p8aSdkbQwZAo+GlKe4A
z6Oezpcpqqaa1T9U767P4BVAGmz0XIC/xk7j2nUgWCH0/fdjaPAV+R0REGuegO8E/eLm9MJ0lVHI
ye4D7olOkFFZtGie+1UqU4VlEIGhYaoknqlFCGCDH0NU5OtBOULogXOs1B/HP4broRDODz78FhEf
myuwKGrbfsazhW21INKQ7m/xxd3sJDr9PfHaggPmpWOT9d1QTdARsHRUCB8iExF7j3Z5eQTz7+Kh
fTAespfA+X3Ke7bFMsruxxoI73yfLd+3EIBZXW9dIqekpCYbk63YqsHHbQylzW+SklFe72zjcINe
ynyZBfeZxTIDqAOGOHOqJJwBN26BQ9b0mSxIuncvCcZXFRW6cKHOHQIA38WwtwzyFJmk03s34yjP
zbf04JQ6ecS31F+VHSKNMT58pj2N/xlnBDf6NkvqGgL1dfKI/6l+Y5GIatGCVWGtl2J+eRIwdKH3
8D1iZKGS+dqeg/aNVUFf/k6+PMQQo1h2Kt3xS1Ow0dsfl3wK1yIk+GK83XWJpbCB6pejsGH/jPzn
dnDoF/MJUdNfG7rPyn26U449U1DAB56W/kIpVgvcrR3ZRtDca+d5ylYg6FEEPJccHyiTqloU7p4D
yDTJea8l73hZWicsS+u0Y6F21xgq7QT44xMa5Fy90JF/HKAhk3ng19rqe8Xr8yknUMx+ZBcwn9VQ
Lby7iykiZ88XtyOufPqyYQr7VMLqAoFz96KqZbv+EFJ3yhStTWyN76M7Yia7cQh9mDutLjLVov26
he8F6tJCmqRjdLcy5QC42Ozq5Op/P/rGhIYavwOWMt3nS+EhALLgQ0f2rSNw3dMPTtu+jUi4qtUU
UhvNV0XH72nNx6HmBsEX0MlYi2buRLJ4PXf2oxXMqifER/bwVHWBCjdPbkT21LzxkDrhI2PY90wD
C1XijN/7g6fTTviH1bN7gsIXEsOSpvvdmHAYFN6AUnScwCUSXflQ9oziH7PZ3VBnQDL/NowgrEET
nBMePoEgW1+I0Iq4ywIDAq/Sxw4KYwSM1FpQEWAximZQWsdlwwWMI42KxRXj2YF1JwV4kcFBwcZI
R+vOTbv2dfppaiheQiIlHDkx9PX3HdxhLuVYMaYohFCLAkvDOZWHaLaG0udHJ0B7SXtxt6DSKvaE
KTxrjK001JPsYYcWt9EPzIImsd4TMFyoFY+cBhuY62Uhs4G+iWHMhwYNKzvgycArHUXZ1UxChkkp
1z+vCaXUWH0IkJILA8GKx8kCVbvvOJM+H68byVfRNbFIGbrFDbVeAno4bYzPi1EzSzAn+f0WAVZs
OJJ+755xIt3dMWvKXuc0hIJvHUAFAgVwzX9yyFAUiPwfFk2gSPWOkL8qLQrQQkWGeQ1itQy5xdMM
48Zvr/s+w4i71eO7hU6/nVxSSj6a/W5S6oafvbiWreVQhlWbmyrKie61R3SUDPg4kjMa8yoFzVNJ
cQr9E+7iwEP4v4AIokUxIzxE27LG3pBChjvnU+D6ydeFLG8Ex3lNliS3FuJ5EWFzPctABh1Cn/ro
9lL2PnkCiWL3zJydwYWFWX6UVnhIvp11Q96yS2NkW8WPL1ku4050W8CBifsp+UL5Bt1PdbufHGPp
Ib54Jh/TP+M+JOMITzIGjnDVxxkyadP/VzECUSPQ/V+0CkPxCdGqueVq+bUyX8yFBTCIAv5Xhj2q
Px3MZzE9ae8usNiQKffKAoQJdXWK/r7ydKCAplhlVTgui0Cn0YskTxYs0Te3YOZAbDbrD0S+zhHA
UhHR9CIVyb2yJIOBnZnlrNKPHskpEvpD+9hzbj7Q0aESHdKbQYtkqnGLn0lbS98say91wmN/0LmS
1iFpBmThN8mq63XpugtmZ+kcIHxasXCBlpcjN7Nju7wExeS6qeiVcXaWnoyFBpYp8uEFJkVsifKB
ttQ3ASwSqEd14etqCGId0Hf7S12ZPcQ08uZTmCAbpXdO2M0e79NuOWk40VSXFc/ARYGmuMz4tBVC
OAdxSDC50+XSGqzmqXVf5mLBNot4ZuBlCt2Kk4romydqQ9/7bOTMyLoeLiC+XNpeHrxiWfiIC8ab
duO+UvnwbYFUiQbhokfJOMGb9MPswbZDQuqfx2jUUhXN9RcH6mQg49ZcGt6xPrBxlA5KKxzFMjNI
5/2MVZ5TDRYB1F0fvghtfnijFO5zjwyhZ08cbzMIggzZQgsHieRoyEczUpA7gUhFxy5V3gvKCawo
uMeGNvxiq8mTDkZsXxk9Xs9W4+eOQz5t90vjs4v47ZaVqBgJ3WsNY8REsr5cYQRlQkah6ZgBA+Zv
uh9lrcjb9Pd3AVVrt8DQL9gLNWpQbdd76doxWpltH3BfLUNsR+7wwcwJXJUDDS1pktdJ8rw447yZ
CNGf8JyH4XHm+rIS+77Orl9P6rTPWLhgHE6z0q2tJUJ91RsxgAfqdZsVwALnB1wHXPTnGRwLJ1ch
006cI6NwYSHQTvT2wdFsA5WNjQmrV5lj2NIPy7s5UdgyLGR8VWqQejrNV+P5n1JKFFZHYHWBGvHD
t7gBSJtfmB75CpjA4VTnmEOsoxfkH6mCaDHDYUtB0x/aGilw4hxScR/fPUgw4J8DHqRvdes+KRc1
QE5joI6Wj7h9nk7iR7p+rz3kKvKhtnhYKLCHTcJ5vvXgBmtPwSu6x5oXpT00hn9weJdQqIWXHCm9
3JglRY87pBnTvKwuOyeSMPQT4MyLB4NWgQL0PxXKnAfrtCa0xqH8HfXQm0tqU2a490wEA8a61YDM
8Sgk9ya7jV1Xzvc/3AgxAqnGn2GOw3v04yZxle2b3DaTtOYR0SO8Ayg7lGeQ9ReW+F5PthPK7/DY
LCZa5ymvjxkq7rl3yALIYyMzgV/Y04kxXgmkK1lhxDSTIbCbPIKa6RZGlUyI9a8NLEw+48QUTOfK
g9kLx8hQ/JdkDs53vB3Vq5R0vkM3+AO5PAJFdGmQZ595Zd7yYPhBd3iFWCu49JisG3+294NyhMq4
JPun6M6sCpQhO9+9DBu0tTn0KE1dYTuESlH3arZZIfJyr0oxMFaYpjiDItHVmCjm4kEHrCpcne7A
pL9vFwQL1HERslT9ms72cNB2JSUPlbA7FbloB9L2B+TZureQdcJcFGjb6aDi4lcDIve9hWpKGWv0
yKN/dLrkLaKQq40iW8wzDz9CQP3XJB7Vp8eHqXJIR3BLiq5uG0QnGKzXQ06+EtEYx3XeaPzgflXh
NzwzH0aXyRA+IeOUz3OVojHoMgky+m7CKLl9sF3NOEUJ9+vqpZB9igpCs6C9SZlpXpQUpo6i244E
tJ2x9Ks1LTWYNbIEb08l6zOBMV2vLIisHvC8vZsZBloSxBo6gFXfbXWVldAolfVhcWCWok58uSPL
7WAUhfH4k0sb7CWMy/BxPULhXHFCbgkEEzddC3tW03u0+2Z2IuWkgM1/dyOkus6u8o9DaF/CUmfe
5JTVHQN5KCdlJYmd3hR/QZrj4bqdudHoGfzMdiQXT7FZDYVWoQV5tnJ1dMa+vpI8ppgLiSmfPbtC
inWvhQzi0x+SY1bdfkw9g7RXqk5HOU0pRIS/Khm4QxTZsSp9NEfHafPcebgJjBBm7yw4yjLrCRkx
prvTIIvEc6vu8MmzJULIMw9/3PO9+nC/Janj/iEFqpHSyqIWs7RGVZ7AJXQjEHUB7hpgqSbGmWt4
1auGRGd3BK+O30ykhasLPWiQtnxw0uptKeei5VKJ3043hwnAuslOq1UnKNVtcG1v03HaCImajFiH
8rgpWkVb9qgB6DRh86NMyWtShjXbLpKwvEIqBdmxDTJpdnyJFayN9ADEensnmyXy7T54xJm6a7vt
JRcvp1dnZulr/Tgft8l/a4m23jHmCAUUzjGODSo2mLLS9+OLVODHBj6ak8htG+sJapEfXBpkYMAA
kJOBNmWwDSQFalD0mR6hOAKcGIC1xzNHlCdk+Zbgju+CTAi2LtkjPmPsJv2KXCcogtl9uECboLvi
rnRDYiWJ3TmruaqHIg9yycORgJiKcCAdOjWebFLWaRuTriKSsF8CZKgOPOBD2Blt3n1I1A1qYlPf
/m0Xqh+bORE+Auvx5EAIoesgiNKmyffhMDMZyJkSxWGYiM7DG4pFE5PHbnUN2gtgQeVa1LpvC95M
+WO9dbJh3i7v/JNEsb++ffESuj9wgqZybpjtSvgoM71k/MGkrFDdKDh5oXfWwUyx8S+8R9FI9o8Z
D6GIruitwG63P3NnywPdbZ+t9Nkbn4cihWmYaoWZaAnFxjIP9DdmrZSF+rOK7y5PwZzcoAnPQ6kT
O2Jq0JEVCRSG9FcMVrh9cOSJ1g8Dlvts1pZJy5YOIEzJt28tXWs2mRpS4ggAUnEcYIa9B4tS/28R
0fVrs9Ji6F+wVo1hdt+xZmeWNozUdbImTLILUY8l4vNXaXLBzMr5+mGYtN6De0alsy4bibVeq7BO
fbOhfDTsK9neAZw/O3OqfAgkZsyrPb8bWaTQeVTYavnqALyWhhazl+py/4aVqnsreaPowLI/Zy4b
IFMihzejXHPZLT4fzHS5FpAiBOj4JzRuF3i6wsm2qXA5UWlCpH8jKucl+qXjYw9rwb9XkHjeCmbT
7clCVl2Qpd98KGVdTe5qaxVPBISFel5mgm9/fMKiJV3r78pnDJ2VbNkVltL9eWDihiCJ0MNeZyuf
0KZCH9eE86I1uNnWNbKI/S6Al0pMlLcQ70dzW2ycYH2j03N8dkahAj+1ldvjlu91pvLbc4/J3eA4
/bv5N0LgBGvVJiVHZ3pNFIqtTJScbtGklJlFwehz5Ij1iDbKDaeb9oPfYMND+x8XFVAQb2lk6dX3
P5GHjv+V+cxFexIYxOLpMQLp6V5Mr6pgzHdny4L/ErC5+WGyEUJ/S6dMDQGX/cIEMzBAGdn0AQhx
S4EaLDicBbaXMkHbs4Un/MdqnzoT5IlzzSfUnpXgJEPK9JCTgneQg+kF1d08bVlHMWSFge06iqRd
248kfzGFb8OhM1LHgU84d/q3QO4JCnVXZIjP+2wutiEiXsIrZ79mxW9AhelsXLc95wD0Crzr6E1r
TQSMJ9fzpjYVG6LCRloPDG4DyyOgN3DrNQPh8bUiOY8mjZcsRO2Ffd3DIFXFBNpXXSxjUdkCUfhC
rUHyUkuzXG2KrQu+ppTyqttDNT8zK0iXee5gi7RmlIYqSSrvrhYsZwdRyKvDr9u6S934JRVxU2VA
8S8eF6vi/cK3awJZH8+kvG7hPvLFngcSAXgE6sMVUKOJgjWAhb32UxuoxEdRSBFlbnIXTyitV8m1
KCxvmEzhS+EaQx/rZM9GSe1v89mm9EPUtHGHGCFCl5CcnGCV3/W8M3NuBUvaENNLzSiLtMnZEbpN
XFDmX4o7C25rasftDvrN6MXfDrJOwFDmIvDTKYlpWSvHzZa72DNkKGXdUPuAOpjhrS6yVDDIR8Ca
k7o6dxOKGf1yIMUmY1HdmvKUJscddRTrkhw31Fnw5zZ6mad3BUdwHjaIDO298D76RHMXt4JY/Wsh
VUGPfDMPORQ6ihHSESmbIEfDXoUJjeaWuf0y3IjVGfsto5+lviy6d84M+3KWygVVsr2b2fdidecp
+rKdhjobDPiSbvZJOdIWjO5L0P2HNoWHDApU34gTl9BHFytpjnI5gyny/pLJJMJU40zpF5ABQ1Tl
20wQf5U+OinNJnAuFhhOwG93OlsxZx5KFmFJHV7aDRf78EVyFeA0SToDqdkwmYo86ZAuwQ4dRXx6
w/64GdkY2TD04pfFAWqKvgOF5GmOlUtumwf+2QEGt8MSVw2j6ajcg1cWeGVPknCwTgKH6+hQ0IV5
++n666EulF1ac5sgcDSe2yaDaoUTMxyFoS7i6a0yHkDs0K8rfc3hXYWnjNBVIX+vK8Z/BasiaG+E
kKBYLbDAeMMlCEnCf/6oVMZNzGl7LerGINYSFIR6H2uGip80JnAuU+NrU6/RZkouQ3D+Wtnoe8iD
7S3EyW9u5OqB5AfBwt8YBx+48zMg3Ul1BajdXIk+6KTz6dvEEvEzPxFQ7sBhRIF6S38CAnrpHCls
7rudE0zrjak5Cgslr3ghPF9ZCADzD3gnGyXP9XzlmXNpXvrhgFkvm09MJ0dIGgK2x/1ANAVhVslW
8aoNERfkFGzaaH3Ydnh6w9vvuVEukhXVvWqTQDpZr8Cg4J15NagHZpARDRz3oQzCKpX08QgMVxaI
2Pk7yWcSqtQp5JiMUVC+IMzjaHAu2S25YwJxLlnBR+nk58Z0W3gs97RlfG43yWJaZr/8JGXi5NIw
J0lHsz+bsS4r7dyYUc9UbYzyiQsvOOaUzHwtwUo5npKp5Smc19l6c+sXa8E+vA2qa5UNYYGVv1Yt
LqDxPXrXfQtm0KIGlG4idxmv2Iq+xoQj/J4ukUUStEO3qxxUPsTwFRN1y+cwk+54tG4ZitKFa8Az
P3EVRLFyFJ9A7eb8emqCsy51Tn/9srOAhH1ibDFcI2UQM6iQcc+fAihrPhwm5Vx1El6F6WAhlJa/
M2rJM9r7XbuXiUkKKSPAC70Ecy33K1gDDY1yLZSwV3gsyjece4QAkX8pqvovFUrlHbm4U8tM5CEu
xmvc1VqjQvqYze44E3vleEvJJvyxWySXUbFxpcfXQTTyCGdPw1XBDXcW36w81ZLZLwT1+FzCPGYA
A2k5rovvSqQ4uOGa9pMmQg2jPpUARxuycjj/LxXE2HbARaMv6nNzHIJsSVObi8PmVX+g0u14f1eX
hH1UrTrDmxv8+xn//yi5ZzemOdbbUiBA+5RXTUaZpfk4oyt+6Sef8xEX+SpcVFvIT++HccFp0KID
BFkBiXUE29Yl/WRHEWRpYCncSGhAeo7hGQDSGstUDYzTYtcH7AjB8i7JoDRBjILhvHGKwkczckmP
di6ajbcZUyqAygvKYWvLRepmPXHTrGuvnH+HGC1tNXxJ+RwZxFTp4WD0uckBSqhCzZTfvoQVr0Jg
T7whiGLLsNstrZtM3YPQ0McGs4Se/bkC1OsGPIyy52x+7a0eYgDIVpIOHY/t998LO8GQct4W7VJq
fZoQvDA/NdRJKvNnJJDtPwTkTcZNpD7rc4jRYb7WMlhzGJZJmn8YF4swsPXnIfdClRDL0nFHaz8B
izWHPVvjR0NO1cT9th3bxcRTmd20lhutRmX05gOGyWJ5OoURP87S3H2PmzkK6A11kR+KYaUHYMYD
eyYjJ62yApszmhcuLjO05BMdbjX0GlW4SRK+dBUb9qE9/a+2v6YPB0oALA9mqKhSCQRd9ml5c4zq
XiRQUGV//4UA+/Jy+WolejdgypD4Um60uaEg7wjMGWYlMY+Tw/0CThJXhyOWqxdLcnXpVGvh5AQD
8HU4A5BCFg8UDE6KtyK7hpPxEhWH+ioUNIaHH9Lfg+8oncaXJuLySPvDR1shssfCZAN6fSPO/owx
aj34w/UmFj8O6W6trwC86/Xh7U9dUdMS1mYChQwDrzcuhRaRXFF71QYT7eRY2mCJuPiNlTIPATr/
d7frM9q2CpmeMKhupggF1chpdUa1+4RUnjSS8wP4umaMvFPYis/Rna2T0E73IeyDG1RuUsP2KHJk
QnFOa4E8uvuPGvtl5rvT2XbYeeSfhDgVe9yTddLexDtN+ojSYOez2UM2UFHYB/tsgDW4okUWfm3X
0jHGnrpEGAZDFVG7Rj2lK9TLVrjaeorwNyrsZLH021CnstyEo6ZpX8rtOlz6blj1joE2TSiRlxTK
a8a76v1xfqZKAblIPRWQ7qt0mvBPsXP53l1xpBNRWeFe9ALFNQ3zluuRKrR27sexQqKJHkzfiqFk
wXEgEDLQEUxDEmmxAp8cbPNohSK0T5zO+L/U7YuTkkRLnEyCOZjkoAbFwWPNRKO+Tx/XKQw2W9LV
NLp6wjmXCdC9RaHsoUMrihib1QGmXZ9obsQPfiSO0cKo9pcnjU33Ll1x17B+OlqVwtCi5Mg7dDSK
DIuVeJI28ewehws/Pb8rD+hdn5EJBi5yLESup5WtdbRBJmQ2+L4ugu6XpszpMEX+HShHhKisG2lK
ZgbsN0enCTq3erVwvx6031l/q7p03wXilShiVDZ01YmvVieO+0N4IRb3QTuLmVZ0mg5f1josHZEz
QtIK00VPS8RdPiBZL/dHEzWy1QLeSCVMdDKmLhW4wYWeUy4kzyUea3Yo2lTSgbYtd2/2KggKfkBm
MauREg34gE/YySo1nlbPnOWG86oBB0EGr54yEtmLoXLgiz8VPJXJRjiltNlYo+i6KgN/0BpdChEf
IdlGK+kLtAOQxZ6xxKxMf8b4SR406u1FrzdcTI6PdtiqptXbZayivVfKpsXfwffvV0lu0Zw1Bo3d
tmW8RjCEVSgDRwiKDwTJH0Ihjp02C7jQlT4nQG2hNCb6gmvj8t/b234Pi3T2Llin5Sh+nB0E/gZi
4/IaCF6GBA+o4R2Gq89orkup1JRamP6a0Q8BVUjw2wi7JtoYvZdP9+v+Kymmcx3aycvXxSq7P00v
VOM5bCKcONvWiGyeZ5g8sfQtxfalXDYB/dvM2Of9TNtbqE2JUUy8t2VMMZySCsl74kxrrHoSazm5
TA6izsmV3nIeVNcE0GsCmWpDS9p8CCgYYMkZ9Gjpu30R/E/c2fxh+a7+2B1270sB8JVWRRPVBhh7
W0e83zi8HLDThVvMKRuztetfEnyYuHZHMqO6ARzQVTsoCioBoCQTa0mE7v+UafgNDLgzS23NXsJ/
GX8LLsXAaSlZpHc6JyRwB6w6vSpXXGBiMyx4x0pGKROssysE21hX1sMphp+kdzvBCJqd1PTVWnPn
BNp3Ypk6E7mEXuRaE3Ipoo0DAzIIL9eu+t/tRxkJGt2T/hTsFS6mOIau6Z1TRgCCtwjb9Gz+mpvl
ZfZjJ0Um3HFCXqtLgpOjbOO/Du7X+FNdWY7BOi7g/7OHfdMEAVGTqJRQc3HSH8OSH2gopkss1bQ7
AkWO67gTDZhwzifIPdbFjYUGu+dbRK66QlVWH7RY20EUylZpuph6a3SU7V2+Ouo0fhaLD1vwYOZH
X7dyA9r6+b/8S6TwwRyEYFuT9UA1gxdxhML2CdrGGiHufWmmiynupVprhQiFF5LCfqrmB+AN67kZ
uUXW6qEBjGLK0ssee6AeyaOcxbEScCxWiWdDv6xQcyOkKsyvgs3oPSb3sxW27hS62GT68GURUqOq
JuhO+owjKJrrO9NQ/KQ9hfw+OdqZJNWlxxh92M6G1wXkJ/BWPYZkE8Cs9tCGXUqp725EoGgQLX4E
ZOAikPCm6RGMJ4vIgzuofY7tq9cl23FkOjwAk1ioatJf0piCvYSUXEGvMQKn/umIkRu5EWPGDEQP
1JBRB3tuK7LKsELT6pZtjOladJwZjbavQou6HlI0vUKAGEKTvgQdkeWXcClyTsZyXrwPdx5hG20d
yHEbx/nOpIyOFyzOij68HhW+0xP+QmA9Sn+rgcQ7YsPutYqAq8Q2mZR6ZaKF6DTNa8VBRp3ibnpB
xoSFyH1+ifnTbQeKXCatEBAqBUy/KQ9xjqGA319BkZaNKyYFZgBETMTmq2ZapqiRGBi85oG/Uh6s
4+gx63oe991Jn74vS7NXGnqHHNpAd1Y2+7CsLxd/n4rl31P7LVwOOTDGI+WvgQjYf0AwvdxtQuk6
bPRrzCwVM0y3x8pd/lG7TwxRTS6qW7hnFPsdlW7Iia1nUxMhzaOgwRtRsK3P/yb4AwX7fMYyffyu
fcMCmdgFr9T7cSG0qXbgnCndpTU5XwUkAQD6C4otYVbugjN4aV13QK4eJPys/CINnV8LEtOu689N
3VCA8fN4zGGxPLvIJ+FPg7NHbtv+iU4MOB7ABgF5w5PfkQB6V+Icr7UaK6tZPieB/USh6AadT63J
0wtJFXG9XCjKdVZxgRfQ2JJO8H7rHnzR4+uqLXnGbszMqdgcz/1C6R5iF2OwckAjw3gGfhFdiah1
MqgixKdV4F76W5WziQY6jnUSLR+m0Lbiui3iZLoV4LJNz4sKGDq60ds1HaynxSpA34m3Nqdjnq0a
LHuxAo6AjyOz9cPRZqQvK0PhLXXSnpoZxYUhFVaTm4efPlQC0dZyoORLyDpoTRkJGw+q8AtTjoCk
Y6aHwWkJLQJAg5Og46PY0uZseIIuEBXIGFD8Yl0OAl7U2ymwt+BBfNSZ7cqLpnxaIH3bEF31Qy2z
GjRj3cmvczIM7xz59Gq6WUITeKIQ6yvx4+xKijgw6B8vDs8FNntky1eI3BWgxtq4rIYe8sj3LIk6
vMrVnnpR9R/CFz2TO9S5Ji3e/rlySS42tzaNBxQP/xTJ2DxVqgYqmBzl293N3JPyzk57maFFWPeU
TjzdnRCShgZ7s7+6Qnn1qkAbb7q9ED8lA+jaAAmXtWVF/4LV2b9q3CMEXepH6eY2CgQCz1puMN/z
w1C7DXM4i/TpnHpL14oo1sGs5J25EugsuN8XGIBKhFqjs4iltYNMiJxTAK2lQBwrPMTtwmzCkm2Y
hstV7c+EHfc7YPGeUYJElm8o6tp5gV6y5FppPpgRtyaBJw566MKldVILmdC1TAumFoY+BWVxA+08
HLpeRABkDCW+HFuaAnXhKcWNGIKYnw3pdOjkEP+qzHay9b0hU4StWSbdTERdXIz0HvqIjXo5aBEs
gJcz/Ot3iFdY2AKK2PHmWqh3IgZXa+DZSQfr6FQqnZJT/4meKR1zfIeAMvVC8aov6X/iYyX0YH8+
DvZ9ge03L/RVvHAeCT7cClqwkHpJyXZ/uWWLYeYAaSGuavZ8YZ0uQ+WDZBvUFGmb7PVyxyTXP5Xg
bdaOvEnKTmKMAZmROZUTI2+KfGAkD9SVuHubdinjKUxB5qnZWx6fnAqebGh8WA5pIvYNjrMqyo/e
hFOr6ebAXMBUAazH0+jAb1qe588xNz8RE8QaW9MqlzmwCqjoyr1fHDysIkvqAUh6+SLykIZ4OiKH
iZnQw2ac2HItl+yC3lyfiS03u03bDsQajIosJExvQUefohrLXrWqEP36/AHp7vIOu3CwWPorTtCC
aDWI4bysavHOFD6sxb2e6F2vuYXfnX9cKzimFcbR3JEddmgWa1jglPsP5sT/bTG8LPa/I7AljhUM
ncYeVKX3xzWj1rbAFD7e0svzrUiOQ+tQ8a74l3IvDAAhp9qRP8quw/pfKjEBdUjvLxyg7fSdAIGP
hiPxV2shs0I+dHOFDsjgZSk7+gRu54s8VgJz5/z/Ui4pxX78ZLyEPRQruz9SJbj/V4Ldc+ZY/ohK
wnxlLrpU9+BOXYWGsUEJS0nUZXykv2YSivJLErfjbaeJX8sNYr0iOc6hMQfig87P9U9+Dj0BZAfO
OOFXeYoUqwt09HGFL6fbwAosbXklzwzkZiYbS8lMcaqRxzwFau5giry3stdPAqxCUy+MYObsRiQP
UbzHg94Sw4I9k5kEQqhvG0JZ4BVpEku55B2OuHG840a9CXpgnHGmjgW/hNsedr+9AYFeFlx2yTv0
8VR7rJGYbFzkhm/KAM3WxSNWqJA4N/PIkGMEoD5B0W5JyJ95BWyqIH3UtmOkM2SG9FjzxIfqHqhA
OkXJdGK7VNwkx3yRy5Wk4zXgS3W+TZeEOe3lrIbo9k0DGvmdzUkSRmEY2lKR10cAAy5FDnElfkex
5+RWniEkLhQd4F6rZm0TK1hfxXAkyZsCsI9bTcJmBZY97GHl3RJJMDowMvn8LFFXzlJbIk2zLfRr
6vMiyKopXDtQvb5RzoxzJP6RcVqDTk+kqG6+tCIgfk0rdB9tgAvzjJKDr1zjrNI1RLJ5whmupKFN
olycEjqw2hyFmeWb8CQyIE13D00d+1BCdq4GMgs8I5uyD3lYtdb0XFGtIyXZqRkj96eLMGLMzfyP
/53311Q3phDe2PD7c8mZV+nHte40UkAswDMFfWWHrrQ4ffSMD2ro6/6XtfrfkaN7HXNrg8cIoXcp
ydJvLouwZFo2uTBd82d0q9KVeKShkAsNNKl3w//pBhxuwGHJoyT1kNx2BNB+Tq3Dk9X+7rqfoA2P
+Idrai8QuR2XY4Zi1cZHueO3l262vFVP/Aeh+zjGO01zYjtDNuVsDBhLOM33OTW/e3VSr2jSa0eT
K5xbl568OjDASXgORV4MAosthFE6vKOgoUt+4hp/BxqC/wc97KTTlaDOD+vTSmUy48Q5EXDnrT4U
4/fl9Tn+zMsm7aOXZ1hjeW9fe3ugYph+RwvZbP/sqU4SUwubSnJs/mLvnZkv/DaWUUFrQBq4M3dO
NOM3tjEnV2/EHun+zv1wrYRSBb5YFBMB1Bk3kS6nXR7EFwVQQY9LQvtxshT7cSbJ/k+WCDMpzLNn
2H1iobNH20uSQ7rX03JzbH93EdQWm3vR4RI20tpxTMbCdOaDElkYk5xyX17NnTVDx9+kaEc2K6wc
a8Te+JY5ig8FkGX2BB9EC6eOHBCrm/PKIxUeY/uTYz7j6qHlyzzbF7FI1SYn//wtI3pVlPyGmKyW
eCywTF47La/4Bon0FyB+d+W4gYlNiotI0PCGL3RDBfSjTOkGmDmv07HC2b/qoNfh34l5JsDCauXK
oywH4kvIDLKCykBlGnxCYe/TvOmVUeXVntmPOvgO78nImRbrB6GyZbLQC/Kzyix2l1pmZcc3kO1U
Xjq6mC73AuIODD2UpVB4wZFWstz085vF+0BK1WZ+mAC8DqB9B4nmzFSuvAUizS553N2BqolPSGjr
SBq/WLC+GP7F467inDOrm2hUsXj9ruGW7hY7nXeuMoY6Nl4Xop2z1MfcVhpAEHR/mlDuL9mYDCEt
JyGpV3k0gmNz7gkKTC5H+c9ddEC3T5YR4/Esc/satglMvK7BCMLpus3LxYrp90w6dioW2hhURbmJ
1YouBQIWggN+0j8rZBX/6vx7K4+9qF3NoEUakI6o0oZsAJQJsr1jCWeeSuLZUSOQMreQbd7uWZ09
YCLWtaUsTlJe0GK2xi04SaEZb/i/G6/00+hfe7+gv7mg/lVXRkxyxyZH3mW6jWs/VKbOLjeCIsI1
a+2VYqGANeo4WjWGqDUOfOhbu1gGSiAqepKvR91OaCnT5wlZ+onWDj3T2Tjy/7USI+/fuS0ifJSU
B1ncSFudjn70pgPdh4JYm+jUVYyuC8zf22k5eZaTpnFyLTHwZKgQiDvu3+JDf2a8qFLw4JiS2j7G
orWWJQ7mMkDnV9ySdbxZ2oQprUr/qL5cYSToQ89J0lvToo4laR4pZzaDaxsghnYkxqXfKNMfB1Yp
Zg8qwFzFVofnoRztP0gYBlbw96ykqklIh73pJNaT1lkS2tjB/ZIlD4K4Ssm1YXcvTJGNHtES2/GK
NWPe/zpM+eEWqWasXumYTr0Dkxvuk8UG1vV0SnGdbjG6vA0s1hqmTfFBlf60RNasfgiUa7x4EleY
4mogeRlxG7AO3kGb4z/XsffCs2ul63hxBlIUCLfuVhqaKfo1aJVgMi4XX7rh8LvFDP8WLbxKox8c
fJf4TVh+aWHwjSRL1FsdBqTbXJk1JEZc4JmMhkvvDHUBD3tpZITYIg6aLtcCykWiFvI+OclwgAwy
ul8Vv77CmAm7S2OTE9xKBxUTY1NqjdaUfj10JpjD/azI00RdBDWckw91Cmi3xyPJQXQT62nNhGsl
wuBStYEWy6zIc+j91mWidzINzhB5dn3uGOU0z6Z/CgA2mPYAMnKl4CEpwQTSd5VdgwqZxxfr2Dtj
XevuQwNDzYKRSW8qoqaEvW5aVN9ip05tUt1fpB7nh25shEReiqmK5AjNiiwZ0TvdQHjWxJTYeSFk
ob5O3p/TgeHSgPFKFaRP0kV/s4Px69Gx2cR7v6lfxapzzxzGYtOHau8SHfSFRGjsgoYqedovEhv2
8dG3+9cGxuIlvybT8I/PsJkQq1zqJOjbD3ffCm7mHgZtT7fcco41e+S/ZNrnK8YjndTsUwONrhmx
AVXuhAuHYRa48tgo/e19rkkWWkjO0mxClbEp6QL+fXKuAYZqE63w8eCTQrBzIPx0mVhs4R34j5O4
jSCELPr/zQGm5dvki76rsAvAYSlE322Bl4y43sqXLHuGf2W8JVOngHGPfcbOhS2EJxRANUN7gBSP
WZMRZlc0SAOgTZr39piEy389OAtVFOeGKjOamvWpSe47GpaO5HyhjvK3c8Jx+DJE9/dp90dZWuHE
7Ahn/Gbfd/kR0sG3KGQZ4RzsLw+Za7xYNg3JcjXg0HohjsAkCtQ9lqPjxkrUL+sCgWDZbS5PrI/p
uKT6FwW/4AAW+1nFPneZv804TFENg0SY32M4jHH7Klt0nS3F4vOm6ZDuLWKAHjXkq/7rlmYh9PAr
xZRUjxnOdz9U4AANiDaBpIE+OC45oU6GSTW0nf53X4BO36rHHsGhHfE2ZHSFzp2YKNkOGLby3LBY
pFjTG/ZM22C2Pn7iryMcELdj4KTwpO9ld9zPZYiph55+JJQkC8u64hxCrN4HTj6957EnDKfgF06A
VyCFESHOQskE/j8HOTeqX2rGCD9BFGi0eF9j7/qe5l3Js69PiVV4dw4dudN5dTAb1LQgtAA4Ezon
TfJDTU3NZ2M15lDDV7f1PdWCQnFhHZC1c8UArIVv4iKjOQW8LeSl5SNZ2KLPzRIf+qEi+S8MjRym
Xsej8bYiBS/R0QdmAEGP4zK7QC0vEOedN/diJkJbkL2Fuq2UUUychEP+DF+QOJ2x7RxwooEGUcXM
6R1+zb+XK/BNoGrWPIKBdm0e4M4Algha4TXyv3MLHZYAdjhD4RTkW2QPjJ3Y3dJ9+bobhBqub2Yo
qhstsZsS5aXPH7o1TGpcIWGLBrutB9Dt7gtyYOOYp7gTkJw72RXbpySRsrhwN7hZTLos2BPpnFP6
H6uFb6ps8z9EzJh5DdkcFyLuDVaLyQ5fJkRnJiv9/07zLV/6Ez08X32YOamnyONVS+yxX50dT4wE
pJ1343EezASm8MW2EI/rSajCN1248NZc3MM2Ztsha6yp3+2b5snwe2r/vrw71T9c7OoJlVrMlfCF
vKg3wNRZkJO7D0g2vN0f2zJeOUPhaEcz18IcuRY3GwTDuHQ4DK6iuLLRejbCE44WODGjklmMqYKw
I8HkOWKgdAidSWXwYKpZtmnG5unxPyCzdpg0WawSP4zzAGaHb42jSI39FFnOI9Y08cE22bGK/gzl
bcgnzw4liityzmk5wPwOCsZxrJQbatffsPmBfrwaoDJbn/tLYr/KldL2Tef0BaY06+07C/aVu/SU
XP4HuObLtMbnVi8DEm7MgkoHBm9D2z7DuMPltylAlLkf6bMiWKbFBFnxGjeVbfjhA3fKcIFa4LMg
FyaL01hGPuv/H2zcdZORzdNiV1wRfgkxd22hnh+pr11I/HujR0daRGCcMaI8WQ06fwLKzANtgwis
6+5DTakyx1RwJpvBY4ZV9xIK2zeDD9xTdYod7f85aiOddX/EZbiqcitL7Lb/Cp3+SFyO99iQbC38
bbq1jDJbabRxZLPehw0XoAwktbASOGK+dNQSTu942sxnJ8jM/vcAje4709jSwU8wMxCT0gyFo+Rn
qzpwWaOvIGIjaH91AarBH4jXKIarr5jWQq4/p24Zo9VstnxlY2RzV/7IcNSsvKIPcG1mMoTZqQh0
sRo+WnYRKFjMpHWUBiuz1WotPX0jYkQuSX+SEMCDqxR62PUJ+dIhzHyluTLS80MWc9voNbb+HfHK
DVj5H1pIkFwWGDrIrlTWMD+FRY9y4zjD8+FqBg9NO/iymthLINQ4JJEVCuPb+Ml9E92epaEhVJVq
/iztpaXto6OlAm/pPwb8SPbFY4RPWOXlS6xmgZ6bJH+x/L6ZBl0inrmMnksYR3DdIf6/Fn3bpMcI
1REziWrUhpFfWrKLP1zNYzXAnuSNmJCUEhiTSxW70Y2i6Izp9vCjXhA2lr3zE3lRYs1ss9be3nTG
kz0PLtRCezJjYZ58GVw+sffxSMrbo3JwSG8jLkr15JsuUIkvj+iwrsOKfyAesyFflCbnEphIvJfz
ghwQgdWDfoAzWjTzT84EviJwClvc4HGjebhYWNCiOh2i+5sohiW5pe3p17hZCU2ubGh90nEaP2TX
Cmw1lzhEqxywhqCngLQXGfbZ3m6BXHVW3/okkIjfKpAT2SrngLIeuTmsryw5swQ/xQAflixCFF1L
ERg0nPscQIfvcIJy0Flkrk/OavdTQeyhezFR/a0c8wMHjc/MMEvCG507BHWDVqoN5nVFz5+QizHb
itw/mhDC89ujYajxafhx44TydKOwRQpfjdwPf6/3bqYMqZlWdhkiYn/JmQpP7GVaE+07XSxjkrY3
UdoMqy92vI4EipzGr5iikjacOG7ygkcqUfoFNMbYPovPDJZvmPk9IFQFZVCSEcY8Yz4SK+E1AUXR
Q0wSrT2W20OVDxUrWrBYs7/83rZhfaMCKEZILOWf8tuwnrKFxW+sTBxXrqDfaXnkFN/3tITax9S/
6kYl1ogxnEddAL0aMvqVaCoEG9m17L/kxvBlFtlkv4jpG1pye0qgSKSOVoztePPhJmpwAMsuXCBm
yuS+htMpwB3p3+A+aYm63+THWKPWnfZ5STtLOqvUbG9IaAH7wud4ogvEUeIvzAWuj1FddO8vQrV5
Sv5P/aUPIBcdyOrg+dPBmTA0OWWdHXh9LSkQzA/6OWfKNkXdKVJ+7iKWAw4179HWUoU11USqp4N0
x7RvD1iM+QYXl1gTbj+kJmd/UlU5NJuDQUSXKShKukdYaEoDIGX6R94F454yTeUlp/w/Lczstuid
OlpzL+xGPD17P5KCm5n04miOnynGIs35W3uLL7JAF3tmRaRxMTgKbhkCdZuEDJtr9v3q7vW9ZCYH
RVve5Nwpn8H0bA1fzY+/oike9aLnDsbfwwZELxwJQ0ZFzyRl4KemEI5UZtP/euE0K/ie534nXv91
vS6RtN4s0APvdS6EkFwo9t9O+5LUTYW6S4Ii82IGFejBnw5+65DSI0LmI+jO77x7ONA0jFKNvBdo
eYcd8ceXgbZhEpZgWQn1oJx6RZ39JsXTshI01rcIhhWZGb6Cs3KEl+RVjtEejdGJhtHa69i7wEgT
yk/7/4L61ScmfCYePBL2Hcu/0bJOHFnfiMq1G/zTRYZmeupDt6qw5cclcZizrM2kNHiA9whKPddI
zaMzB/7S1ecoKDyF4sP16fKkNdli9/DAZtW84/o0T9WijSt9eofPtUTyQoAGn1FZ7KmBLgfzxOv+
bUdn77dGlW0iqQoAr/7MMTRdkBMVq63t39KzLP9KRqDt2/Shk1UXlzhHKHzf/HkIyga1Ul8q2olm
iYtf/KnnzhZmsKFht0AkPelBP405wcafYBZwfloa9TGnXaDC6EdOlQc/IPzvjQgjpm88BKe6JxoV
BLYRYg7cAw9FtGhTx0Uzz7sx8AHYTssASAeNPhQW2SGEkGqZSTHv3HsCaAJyRf/SS+QyYVOoF4Bx
SGN1g+LpjstgjRUId9tmrY1yKnMWVHSxLB3cxMjWqI9rXR4uz5Jv2/yHzuK0A9R8PlORDKrwmqYU
abtxz+HWJPjnfFup0IitnvMuMxfV7JeoNcgsSqDQQtOr3TEZX/WJQvu9W80oV2Cs9URtXmnXrkQu
cN0gm2vGoJT4EVDVWCAvtah6kFM98ri66WFgxgARPdOd4b3x/gJqTXN01IECUbAMkDtrEmupj7pX
eyad7X5q4VhzuWSAXstiAC1xaeIAaYoaYi77QAOJHYEN0TWuYQUEXMAw9wr3imZtjH2qsU15HxQg
fr25jOzG260jibDxCQ7Bi1uOkLGbzWP4tWbRnc87PWoQBwGBOwj2ZmQ2l3uFEbCkEZ3N7zFDnydo
FT0LRaFlWkIoj5/P0Ysz3Fdsd25jFm46vXMv0wWpPv2LQVj4FGGqvKMM52O86J/jvHkBQ0N6qz+i
mhDO3nfGi78GsLWkavrs4s1asmEGL3/jDaDMD39VcxK2nHE3bS/fw+2fk846wxjgisArZlczVfDf
JI1VnCdVfkl6q49L1HJnticL31eg2iYbh43oVqVVPbRcIL4Q+WOmZaKHX5pz3jdom2tCjFe+OwKS
vBDp5aTc+y7Py3aDGKE2+i4TAStMV0Vo7cM999BI5aucIVO+PL2DmkIQlCm5g9mJjLTp7INOJzwD
gMPHuPchlhcAarlPpcCKOtOd9LiKAc2ASzMaxWvNS8gcgDA97+w1126bA0oMdYaJ+BB1PbjZLbiq
CAJhMCXm6oQwQZAMoU+KKf2+LpPfAjE3VpY1RZbePUMXAgZqgkCiH2ZWFDiPGu0ah0Y4u3g7TH2r
MfqXBmzcLbMWFLDwXdHELnlkR9rPCT2Pm3unSA6akjRlGkZLtxBm+jL/VFhGlSMRrQ/B8U4+fdA+
09DDhRJT6AnvaKMrtNCyI7DalZvVms8ZI0wcnXReiwl5r667AU6hELDjlHBj9kdS5thOlEAeUTAJ
N3Jb4UxaOb0b/sBThGADT4JjT7InOLTsWGb5JKXliVwl/kTrYC5myVh3S9j1foOwx9YFy2IUFKst
r2yI2TB+kA7xWvuqqVLWKK2AXuY7X28vS4/hnfDwVWD46ESP27rG7dYb7ugDGA94Wt3LOt35q24I
MwRciBtD/MpKz5HGBkbnL2IFNgPFrYpqjFmD19oBhGuat1B41PIaRtuxSRvBj8kCRBR06/FbX/Yc
J0cWScuMZGb6Ifwjc6zcP9F3ozT32WLHPJacFnoAjUBW/RWPfdBD8UMVNf7jEJDJ/KNwntQWMmiY
mrSJBMFE8oW9fnDhiJWqh9WISuZscbl8Szs0xDRJZYowaOm19ZtzujDC1tMj6aR/2sPAmnrNiMDN
CHQCVbbiHz1wGicpQ41VRfEbrwXeKOGZDz5k8Rbrm8FJVXz+/lvgR9aLsNA35RS5B1Vs7RwpPJHP
TL2yzny5V9BYDITmf4gXAMOr4+roSmR+VeNbVRT9moG7i6MeaWG7XJ0pVUnwtH322tMOamBITvid
3jeE1DWs+MG/NvDCJwZN9TWa0WP/Y4DwEd/m5e2stjL+MvXy66TbGmdT5htj4Gu58rr5JX4sitl4
3O+2L1/1Ypc/STKfOeqLX2XNApGreKqm41Ok2KZq5yAG0cwkZmVSI1zSCwnjX5tzoCu4UYkTg/Nk
o+Zdf4NrmDqYIgyRhBGpxINWG6oxhBF5YTN/JTqzOumIGm6b/4ahAvFbxsolK8FFkY7bdYocjMAO
4Vphu6gwLuPW57PE6IHpJeI8PHujCjNVqbkkfzLol4jU2PGDA4o1bJPfOO/7vmeb6rD4+POo1H9i
Eg8TLMB8HnbUIru10H88f23++693NjhPZwC9OEu3IwSPvFTMJp0O7Y7371YHhogg1bivIXd8h/0Z
ksiUiMhOoltS44Fsa9zEGoyf1M2DiMTYh6bYGirQWb/Fdy5uImgqxvXAO9B3XwZteuQ+TnolIOYi
sh4JDASCy8B8gUHmPmULnInvU10tr0wXB8xGkq9dMgwCk/PoHp7zvPOJScfVJ4V6vKvPNyCdF2MX
JMcybp4l4VqgBcgoMii5q8kR0cvOii0HdnyIHPOCaR2FsKLeCZfyjbaB33cwOBE4Z3ytdx3FjqJH
e6sUvZFiadyLGV8z7xuU+djVfa26A1yZgiEcsNtD/ffXppRT8qdUoax6ro964n6um+nk6Rnj6L52
b+7Qr+qGzBhXZJdl613nuaTHjmtDtGL+Ft5QjUFP4JMWSY6CN589kV1KhwewiS5IhvyAjqxGRwaT
UzklqptYUJ15kblKMdIlRCttDTeiezFIKnjiH9Em3fDI0zYrcpM4Q5iiR1jJnrA5sBjzdiNmPbio
pYOIxQS0DsCo7jmflA0bk4YkcivKgtfCu17st68E5u7u22o07NRWj30jI+dY5tsjCgLN+vtZZ6bW
9FLbXpKii7EmNOH5DqhoNRZKUdIKPWB2K8U2rQ7zk44zctoedYz0iKg28ukI7zoZc1hJzBNP/InM
hiAp5v/SZ09J6+8a4qYHkL6B4aGFYyTcbuZplAfM9XhJ0/4wkNM7JRBI6sNJrjcFJT0ac4cx9xzG
TdY1uYeNZpC5mLDPU3vLj2wozLj1iyRFwX5lx3GZKXv70/FFFzHy8rRjOSQUgkcnBVUHAdkFDMl6
10omfdO7RVN2nwH73JMe4ChY39RXmQVPCTNPJmDHO6ErAjtNcx/kpe6qE9p7gEdPF9qPJaX5c03P
+3wqEGOfriksrsXQKB67NBAzdirO9lsHCBRHO1oeD5e1CT/i4YU6cBGsZIJaj0uBevnlPlHGkLK6
mAsU6u0awJZ2qH/bdspRMJ4r3bPnrw2HVlC7xy/TmB4FRABjvSjtKmoxft/a+s58JTHAT4RR42xe
EvxFYG7RmVQ73sC6RYCT3AGeAkeQZjBzYSueS0k7c9qISp7BgSC3XX7Wt+L/dS5Xium5g8r1Dmbu
B9YemmjQPYoNJ17sUQuwsqndsu4ebTUKJOIA8hi+i0dSya2g8CqNW5Ju4g63RSoiGevys1DKT8Jg
s1bwtVl5SF4YBjgqFrme3nUxYCC5ZxkKtlX4QsLjf0B/TjiZy2UofUAdRZTxmF7tpStIvdFB2ixp
nibk0sOVJd/Nl4ShiCxngMRs3B8jWRtWRQqzRj0ppbRitBpZ5MeARbKRDVzzrr07Ak4QaLI+U5z1
eJ++dntpBvxY7bZ+QDe3Q69L/Wb2PA7fgisBVY5tlMRbcOEQmwhr66RnpHjcWdyI7ZgcyVWFeaFe
9h8ea9CxpR3omTCJA4gCgw7xTCwCJitc1m53SmODhXNnNCO/x2DgRNlVxAcWJRKUc+HjqF/KVjsE
keJQ7+1G8KLCTcJwFKdOnuviWcS1evzSPNRHZuSQH1Kn8J3+mydXrWWHDaseNHwZEgvzP/bXm0nP
TcONNXoYgdMrI2mLiX7lKo+nT+nibeh7GOZxOdQNfCBdTrjr9Nzhccjg+ZEVEvG4XjlzHnz/mBmB
GGF6GKPssU6aWUFcQaFvENqDei3qWk+IkQfC8Peqt2C+/YaDcjMGHJj8mBwbo9kxDqDkYdyVvD1e
sASWEGh4/03AKN2/OHAfyGTiiwEwJ1myGe4ixnfs6x92EtvzaNkIQvOrkdmgjtzS/NDhhxEltPTb
xDF6GriJYGchc/xhc3K4S7pD7NRiKT27Z6KfX+dw+A7HTXx53osfefPtVArcOqGLNjUmDwner4jc
Tqc8nx94gprSsBPBWaavVxus7pcPIuD7BPK49vdq5KoeD4ajKXJMxb8bGcIrVLgg7BNt6suF5zkS
1CynkNZkhxo7xHoBrn3MrHyjZ7j/uCFlN8zF9/QSVxchaxK61bTwElo+AF7EGXRwMGqrLOESS5no
d0/IHLDFDwZR0bu/8o7+hpVCatdBmGc55e1DvWFioD/43yNOT2rhMf+NS2AaDLMjC/bWQc98OYs/
GUfTigTrX864+tTcyB010uTYSe5uSpem68zR8yHG5wqX+p0TmiTy/G9GSHWe3Z7wcokRY0Oldh3t
CjCWYiUD5i0QlCW9ef0rRl0kuXAdzOULRrmw1YSwU4xni045bg7I5S5BL3WV9Mkl3Q0LGNsXoVkp
Wsi9VarTBs41xP39v20xnRv/AM6H5hku38+LqqsKdNJ8/JlJWPti5+FQ9Fz7KYt0VvPtgkntD5yd
NVH2IwkV4m/4Y4aFNlOSbheSLk72UtTOX0FeDyExVaX2D5U0sbg8+rqaMSIzxGcY7RUK+Vm+mnii
imtv0m+/pzi9zdEu91JDOuRZGj4QapjFmtwsPgHsomZ6W4i/m1v7CXqcpNxDn5vTDDBrjDXsDeRi
siWF/rxqiseIYQtdOly7yhlFjdS4birbFONwklF1rZrKamnzNBLynMMMlw+benW6YcxncZhElb+w
0BdZ3TxAIC/L08gwervmujNtJgESlxqYfciywnkAlF2oEGKcFs0DRrd0Aov+3pr//wi0q4OWFN0C
EUbllKnFV6ou84TvOLd5rrsUJI7TkBRokT/YMmib8DC8e/v7bbVUmb2XGNrbrqyrb2x3drZopSjO
iyun+yvYVoCTCL+niysmEiBJ2FVdzAKussE0RnX5SwGnK3OtgPBR7tNrxdNi0osindhvO1DyMllp
Bq8IXfGckyvTYm7UBhe0DdCTL1Ldp+es6CR/Ac0I/GuG/40zS7DAG7z4N5IkBbwcUjpiEbwVduiZ
j5drUjYZBxe5TcNzdM+toEkjW8bo71A5wMtdJvUHuPr+yl7lNO39PhpJt8OkrbfFJziRRDzdv9QQ
mYePcwkrV0Y6I2lG6W3M0IqmngZOUJOIlBPLPxKtlGy3Pr9eA5LgHg2MD+tAxZS5B0MdNxX+C+Ba
WJwXzMYuPhpCi+sCngZCBw0gAM5Ddcd5zZFQndqtU3NJnbZ2V6CXV71jA0YTNLqbIcDdOqkj4yrA
sUhtZbIR71bVp5z+2/zAWBP3+DscNPoVCcww4qtORYkoyvuF44KUfKcZp1N0NJ9dlToWlbbULlZN
mdHaG2w3tzy58rWGXuBn9IYQ2rjYoPaWVSlbLTEKj2mJAuYLMC2jgBN5fTA6d/xFXbxGJjGkN4bY
/ndf3Nbynzvc+Mn6EsnAyiBrfHccrkbPdPhXhIC8N3SgjJ0QLwVPNBmUw7DmUEf7n9eeBSG0kYYt
v0DeWEpX5Qr7ZJwUIUAghzhr/PC+I+D+HVCIGnxvT0SP84KbXSY9RG02r3PpCIfRqQARxSC33OyD
Wk/UNrSZveO+tdmWWecR9VrZ1+/McqfJz+0gv6XKOiWi96eOWUP6MA3wxX/VNOv1ZHT3H2huvvUd
x731SpHzR+gEWHl+Q5sPUhBGUW8O8dxHxZ1k5WbHinc6vrF3KAtnNeZO18TVtGI7Kk7rYK1C71xX
VUU/VBb4te0NsKtcy/qk9M/MHj/jHeareWDmcRvxhBfsZSDFua068FvCZBdoIl8QJrdiO3d/biUb
UrQa1nuJK+tMT+DPR+owUJpxdEkQqzOEZzVUqqQH7/v7NVtGY62AgrIIGtGwKm6vJ4nXwJun65tc
BKcaWCNuM3SI4gEwmcei9Io7/5r3oHy0dSBqPToKm2RzUq2wIklzWXm03KvwfLnTgnez9bFP1x+/
VORGSFQPFVwmAaWSEocfFnL4wYv0rm2lcBlk4kNVlrSBChXrMQLLii76wjuBRveb8/S4b7zOjuqH
GypDU1et0BOflwebzc2vJnjVXGa1K/sa0mMws/10YrY/6JuUWgPovAjPOodMUKH9XwU91IsUvmig
Or0mPHrR4mJzAMjl8Lb/CzOh7hmIndEqDhMyyD+ZKqTK9PUrom0XD9LSH7ZzBawcpctRNvA2xF60
OjSs7tjk08Q17jZ8Zmb8/keJpqTW/pr8ihIAmoblKdK1QUofaSC/jO3NVo/RWjGGQnuvsghpEJ4h
wuspuwKWhQQLTEc5ySFnuKXPoXFgENKD8oLrO+UfC+DaBCEw1/0W5lUIuR0Q4qPN2f0KEbev8urj
ueKvYOtQhB1R7Ebh9c4A9L1puiqPNmoaFHgvdM79lF4ZmpuSmadUdJqTkCjU/MJ53qXCrMPddiD4
FCqguxbzbevQGfwKnCCpQ8InsmzcRNsMgmEDjpX5SUymrn0rTEGJbwdQtRkigjfaUI6un7qquCfU
Sahfk1+z5jvnPYDcTGcuqD7H4eScdCWHQRZDSOK08uwi8yW6eXkg6BDTZ86rLnaRu+91/AqSdwtV
aTvJtBU3U5NNaIZdVEFzWLdrhXytzbK77thCFQgQK1vQ/aV9HqRxvs9PHrns63MQSBIP2vuOuE8/
4ET6JXYwvtEXsaDzqsGTMLRaCtZMvAj4gVVVfawtOz7WLeY8v5QuUeZ2kzYxUAieMZbV8qn/Ffpu
ox0vDVHar+M/D8Vm3XOPxIUhs/+IX3dmhk6MmxQ9PmNbprzsARQTVqbAcK+rB42ywfsohO+fmQH/
ip3mpG0PxV85wVHMN09R9WIicRiUgqGL8647kMX1RImYS01nhW6Gh3tr6xAIPTWp8NRyAgOESE8L
O0RTQL4IfOWqMANvR+E/QCbJ9++wujJ6phsS9omkVvFePhIdzU4Ylze5rRFqyAPhFh+2HWuupZQG
qM6g5+YtKSVEXNl9k7LLKz5UY/1ceBkMDkpNZZxoPdUPSGxppHEyzlnW/uuykXhhcTys8gxFxcSe
Zwz/9yLfKWHlfX2G+rVp+7av9+QCG/XYcE2ZphlvXUedVz+GSbq7YKX2LDZj8j7CgjvDaWwL+TeW
f7IIxLITSdvwY4MA8WwtnpzfxSeZ8T9Ut3EmANuk9XTTauY3BTshU9lEqLVC1ICY4fkhfWLW0iBq
DI2mpfER7xaTq5hkkOsKw5UfXjIgy08hefxsqMYDwmHDFHshMjWXfatirDQO/cnAFNrE3md7rB4J
zB9wQ680rPSdCHtL0JFLOVQmjyqHwht0U8I+kII6bRZtb8SWCVgbZ5svhWELTOA78N+QcsRx377y
KXTCG0UAyY+CG5XtGiK7Hn4VH0n+rfIZPhTMoi2AxHU3EU6SG0Wgo8aDdJXVEU7JqIJwFfs1IeVK
hQAY7OyVKhDQOWPTh+43Yf4xIxiz3Snc9+euaTKfQWh/RVUbN3vUcXy4/rsPGawaNeT3ADOBPOgA
cdA3VIRumcDq9Sm0r4aacBZbVfqsZML9DyfHWSpTW7Gp6s46+LmRZOh3toh4o3HXFeu53GtagBre
FI+3ILXE0me8hZuW9Bqh0qPRcggBYmaXEP5ubAJrH/btwYLqQ/m6Zg4DxY/twKy9IkzAMdyx/ewV
TeiBRbYNli5WRNo6Bn+Jj8cb4HYTZhyDDaZPD0Zs45PtwAQr9aAmcsDOeMwCZ2xAknhT+2DIFmgg
v9swHG5MdoA4zm6T4sfA0Hm7sdWUfX7CAn/DHfqZV8hlbNfKMF2dd/mJGudviogG1EGlcJW4eqAb
w3/bQ+W61S1iUAUsHgRt/L9b3ukyERuwr1Y8o7CAtyufEL01dEFPCD8+zlEISUpqObpxBJzwtG5b
16uhvd8aTnwv8xAYRfXIB29lMRIM9w9q6xSnDETFVRliugep/l2/+XnLe+W1/Co3oNqw1hXroqJQ
HjnjCZ6Sfeldq3EIS/6Vnl7InnlnJ/8+hpRlanv99h61RfU9zTmFNHLX8gaP/RHcOKG/c0dS1Z8B
D6ThQItw75jLlZUsJYtv1NFm/13Bo3qy5iSmn5stcbrpC/BDw6Mar0W7BRZCKnkoPji2Eo65jKBK
ljeLBcP83XxDbLxOGOvOGQ/HygNNYOS3DHO2eqIhwOSi7kNsnKlSmA3VaU16e3FDJQxXh0zLdkDd
RXYM+16zDdLps77MwpzH86EelaAKbIwPicMwHIPJT1yHahu08Ne5L4bEhlICpCvwL1PTc6hpt48I
iLGM/7PAhjp8LgQnH1s9COFGbmJfzpqqGcQumR8vypCfwSZa6dvlm/Eo0MtqnvZxoIg0RtRdhqjR
9Wgv5doaoEz7oAPhA/FdjIcdTLSBOb095JgVCAxjlxj3DLtCaJaYP3VExYTWeFBrpZKnoNa+Nzpj
3JpkaeHFonp4JO8o/pzTML3CJDS+7Q3vVaPM3pGOmRpWyZUmXNwVzMDIdPdbnzcoVt60k9JSmCSc
r/++iH6FTXCxRSBgoWTbf3c1iPvs9xFwqaB+FpIagf9JAVa+qcJD3FKWyXiqMyZbLZwmbLNTnI+l
n0aPV4sngk6EsRMEjpLTO6uj9gwg7cd2rq0D/aE++f07BDgXxIS4QtKWG4XelSKonBr2xYbTV0aO
3Qh4iCLCYZm33rdHhLd/DUyx4H6MCFoBQsGKUFqibQoCQ90PtDGTAnVvJdm4gZ+vEF7jSYEO4aQJ
uMKcS3BgLIvLG9aWz4hxjNGMmVSA2i6jcTiJgMQju2xJejeMb0hmffTIMnqvDagDXGULSkJfWbTR
CYK22WawQmrS42+5P8a2Hi5SnjPw8hEjjTVfGIXG+zp9c/CkItwAQyv3M3MhwY9KHMfzNQDOT31b
fAzzqKVadAdwFZ+wR7MLNgvY+7jNnsmJ+VFgEvSOaUH8bEnnRPXmH+9HXwqZc+diEZRBlFZv5teF
Hu2uzQVCbyPZC6hYx5po50/amq9fZ+z9aAOy8UMWV9HvAJTKloOSi0gOgw9BnixloUZIYlotET9g
Mh3JwVEWKZU9xPm79N0mHLNYs9itOzar2VePqkz3z1/b0NLwEV0IxbkU1wUA8Przt0d+/2fZ8WPg
+tj3RjNYPq2LhC355VgeE8F1dzpRRgBnpHiK3CwmVLp+CSLbMBLdHl50ZVZs4llhBzjs7kPcJB+Q
yCw++CnvDud4DxyL5zp3vyYWxMXiFGjgns5NY8hNkKG2LXuFkZsYMRuE4WbSfb3NnPvoVeaTrxJ8
OXcVgVJQNd7T/OD6AecekjAAWkYrNSQ5Ww3GqJcH6YJo8AUHRv8CD+LLKv3JSI0xy3145zC5hRAx
AARTR7JsUCHTvvslOdSxH/YPc3k4yjXrZGQjPUnSGavzJEzNVME/lgsRa5ki7VDYUG5i3eOwxL7J
kFUGtGuTj85/bYSCjBNNpb31mtj+C6ZRx+hqUCaJCoz3nfGJG6X0y68OfP5D7XBbifo54plHMWpm
YdTbg8IRopCBWp90NOsBm0PpGbzMJ3Sx/29+bJcQoIkGryaPiaBPCHm9DpGcT5wJUw62voO0RGIU
dXK0ZaaX4TIyU1d/klcLzYe7ka96mwe3E/uv0h1zEEEwKAxnJd3LZ+zTtpJijk7PfoAoOHnJoufq
tYoVDMmm+FhP8lOAPU75r0OLwyZx8EO3XkX+4GT9A8DBjd4alE1N6sxM7jk7oByvdNUatk+OUKu2
E0I7FpAIXsJ1lzI9eUYVV5rAo5Ocvi44AKA7SPzcUhbH6YwoosO1bsP0wWynh21xO3hrzsMLa/4Z
rT0AtJ7fLAg8keU/OTzWRQT62FoI1rvy7PsaqJVHmouen9CYB96yOPROrGsmiPT/Uh1/90urmloH
IDy8Ju+BBZy9aWfgSY9kNT35iSuiQlVkLbD+JkdGBtrWiolvOYEek0BGflz+/jld+++g2NvWV/QU
lsZ7KXhkLUKQPGXpDFpR51C6HfJ17LcSrqm4IBY9LZVjQPnCheCgvkYjV1h0oIYZ496DYtztNhyR
vN60kSw6jozQu7gksU2JPmzzuVpOJDGDPAsjqH5bUQ4fbBlYhT2aVXv3CpklcGjKDLX1IDOpC3VM
2fWm4PgHkmaSBekTf9I12oWbAoGSiyOe8tTXLCyO9CUqTD2Y6hSFWyzSjChviPhQIMyMGiqwM9oV
sazl4u0r3EmM6h7RUTdA9F4iiryW+zWe5ztRKRls/dbLJilwKJm8f5EX9rHLRoFCEnsD6WzNlbWB
m6jcpQX3iDmuReQ0Y2+08cxhDo7CW8OvFoowWcB+jvhv+74GPmIflvfK/V6DDCzLMhg1dwf/sv4+
hu5iAsCFJr8ohDaHI75l7gtQqB+uxk3owh1AZ+iB1zHToM4vLDGkUCb3CRunApVeYmE7fu6JemQQ
tyLAi/rcp40c1uV9gsUtlmY1mmb/u8jATl5sOIuSsStoPi4yikyvu0DTLnFNAGUZ1vmCIhzC5Riy
9RHN23UA1Rfs2DcdTJKJ3FXBSpmEwFho199QdWwDGXxMNOs4GBs+e/kNTzszSGLAB2Q6uLy3XGPy
uWSrrLDc3NYln9KLtkUa/smqoQ/8cRjTnIDuF6bjRT6MMS82U6belJ1JIETwRXm8WiWhqv0VMocQ
vv8ga1nnw+siyKxWvR3/VyE75K/y7DIWrwlCXpbr478zPUt5p6Gx9kC863/2X+qPU2Bckswm67hU
ZUGCiSWe/YoHUi03PURK2ZddShSQFiemOnX1gZrJAAFQtpdHV3Apor0es1gFO5G6sTorTyXGcbF3
kqAtTIfGHxIl+w62CbilSb/Q+5pG/+kAwg7GRjilqn7mWPoG0nutfG8LhIJkxKgG7s8HBnMlWSp4
yTQ3s/YOF82mZZSTiKw9NrYx8k+b8wqXyEmaz1EIc54ISHhReAX+JjMRNqHzDSNtl+VhaRkLxI/G
KZVMPen7MOuJVzoXfjULfBSvhOJx/cZubQQEkmE8Ju9NisswTsCTwY0fBwneRgvLfZe5fOFBxnCp
InYUa+zp0QSAvunsCGomhlgK293lxGKt+kJLO33Vq4brgfG83RQgbSg5aDFo2Nt120wKBc+r0zXh
i/PqdpaXvEFjdfhn1Vs1e1aqmFLxppLIMEoQQtrklZE26liY/uyaAhTXjeVOzY/tRIeSrtdiEZI4
lMHXx2uVoaGDKQ0CwNBT++XrxkvDNZN1hi/hcStrRdIQQXgWnCt7n91DDqmQrG3anXwJ5mDpU/lV
uFzyJvmGxOk16zYjpvR1cxtXW83Jsl/xnMxW2R9U9WgwI6qNYt7KHvAQSBV1xu0hQpmAny7xySab
kkYRMgZBT8/RfhHgwv1fHO/IQNYxY1fU7nle/unC5BEFRXIuz1oeuXs6xiWLKrQX4nbDyhJBSl0g
Tudte6IguoXGcQ33AZGIlIqnMuKA6AnkPEloUWqcZjTfpD7f4ZQnEZnydkgpwUsdiZ40fuAWvarX
y8ESWOs2uW5cZNhqY13yvl/N5xYTE7fZipsQlyP1SlEYFbitSDM4Red27zZKOVNyPiuaAfH+xyli
W+seUVcKhmcqPakL5ZPo386tEWE0LF1uLstVTk0Ku/UWUz5fA5SKOpkSJ95l9M5LkaIMOK+hPko2
T5T0W0QW2RkSdrwkaqPmoitYIsjrO4vOWDbslMqZL6i6hvHzME4qlr9tqJ4c13vJFONQssvLueCJ
JzxKDIr68Il+yww8IlLk+3wCHFiQlTGpbfMGj/M3Bja6W5ydQAYb9W+Lz+YeFBGRcmY2E8xjShe5
IIByLPHMk6T493TFbMzrE8uBBhvCoAGvrHrYAQJNDlIIGQGVsA5xZWpxHGmy7kGho6tTScVIN2ie
jSLqHHPA4lNrzY9NP51mYWnvkDlgbLzyJYdoj91JdLIhyxsu6p7GPT65g+P+MKzWKYkZT86gV5K0
m0Uc8wl9TbDl1hb14w82mwmcRqADlmgUFmaNtQXVGUn9ND4ElikCCp2qKkP3ulS9MohtWu4bfBfr
QRXjGSTZMiJ8MqWly1paCTXX/zZ0tW4kHKZ6tO/Q9mUDyWSO2wpxMkqYthDwnLswwt4OSbO973Fr
/hwsru5sQv5t+bQnQq+JejEAsb1hMU9oXOrEQphreigNZS9yH6TRZRBufjCeTMfLcWwT9ZDzyuNv
463vhiVyyehvPuu6LTdFzPacdejrvJo/MM5DZvTnne6YNWa/Z4E1g2heHwIez95WEFK4mpsQd9ff
ihtdgXvN0X+QgM7uqDWxdHSH9HinLmTbsLM7mlcHsUtTmW+HyNUqs5F14pobXBcLi189FwIjv4lE
HXDU+/71vk7MTvD5PEYlgLGHW/hJ4kSBVcq35c6oeWmQPtKTpSXJLhDvkyHmbN6KksBEybhd6KZ9
9sEOVs0JngVPSsF6CjWDprOACliYDpQf7hIQ5dXYMbBVOFVvjF/RPPHFo14M2NQ1138hAlSJud4v
CfsqZrR8FuoA4y2xmgknTKeg7w3LovoKANuYBqZBpxYC4q4Q+fEaZn05ORByVY/h9jJM22VOjX+y
2GcnTW3rBF/iHPzKuioWwXFCeF/6tI/sMTzJZcZPhbwbJnlaylK92o9VGkx9wsd5lv7EZdy+zhU9
OF84JqSwv8m3GD/esdVqfhFsPbnRzp/QONwr9z7vr4ax8TYqUccyb7SqnKDEnMIm/lXeToca7dRG
+qEbfT6Rex5m4hxe5rhNd2qtu6b33/0BBHiNs+XKGqVhUH091eNfybNI2gB9wbamp+9OnjiFHRHl
0XqAg4ci2AJ80penN13CMP/2OgmBuUtQSXDRsjDAA7mACjDl+tYGdLWopVmojPED0AKluL41plgh
PRiJDk+3SumRjL8bjYeXNZJrrOrMIn/Ru/wQ+zQepMrZ3zrxfXj7JiLGDqHNBuCU6KwAcRl0XSLi
r1FqRclsVfJK0QQmNtcSIBhHFTCujnIdT/ptSyU2KEUMx1LpIycHFO2TO85qf7MT046x5sy3ILIz
QKAoBT7ZrsPHJLVtnPNBOFE4JRtpMKXXFzQvp2ABu+2N0xeoK1gB2Jlo1TrVpCTqhAW1FSAKtg4e
h5bM3Wo7ENxvwa4egmCsLe1Nul+FUQ3zVqveQkDpCoUblm+PV5nyeeITyjNBFHMBohbeptQvOEiF
5CEl9FJ7sN86SqQPriwmogW8r4xMX3/YXij4AL4Yt+H1cOU5Vco1zM0EN3qhaAcPgT1guIblqQBb
m90eeIBxs1el7jymTAasQNbh0AiXZyzE0SKwIy06t5ZPfvBOCV88C9oBTXgEhS9d9sVbhxciC7ES
Zq9nCkgtKuLKs+jWxrDFAuioHluwfxKS/bfpY4Ud62S7uzOunfg6bG4sisMqCukcFEzoGFwKF/sU
ndf2L3mCPRAUwjefn7kDMj9fBWMZUqv0ut/prTmmDafq1rcrr9ioHsNRUTam0uivXF8N501u9SiL
h49cruNmUuB8nIqrEC5YhqVDY+CUC4LlirD8CvIgzIIBRfQszrmEk6WElPyJjRvQnTuwTv4SPVbq
BQ/3MJ5s5YqrVU1ZYGQ1AM3tOMLkQjDqZ7kIoCZfJa+AoxK4AY165mhLspVS2mok2+6YKwza8MP2
fjYy5aFpMzeLcx3ajIPZZVKRXyZ88hmPRZQnH/XsBKvvrPAZnnOtAXkip95kIXm4tE9h8clPhVSj
uUPrWmQintDmT63hkyHVlAJluMPiyS8yPWQwqLwQRkLLwIrBSMLXzD5jSEXtbhMBUDuihunp7NpX
al1MGJoBm+2U9lJ8ILo4wb/uWkXnvaXqmNp1oi8/T6PsU4uY4FfVvDrxQRpqreBedHa5P6YzsvNR
dWqFSjLRt61uXEQAUHr62YOtWHgEbPk3uU73/lYFlkkbBt4FtWlmWPy8efLdg5Ha6fGd86Ue1K6w
fGTzkV/6jPLaANHYvrDg6u/9osswFjDOAvgtM4Yl9fAUOHcGylM2K6slMehP26oL2Ve4OUd6WEwx
MzVxRDWZKd2yt8o5lPAPr7NKQgyfiGBsQXcAMlw2mULHtjGV38SHdOJNObIQKZgwe8DxBDMZX3Kl
DXHEidhngVRVB+P7tMcuAx65/jSLc7zt4c5jVHQOfnn3swChOvqKcAYFD0Ssd+XbM4qd3Yb2U0gX
z2YOUGIk9WheMRXWFiQ9YZFBMAnXZK6WywP3b+6RnvOAABs5CsLxmbnzbSGHOu5lKWC9pZn1yTZE
YcL+ksy+GUwUHUy37WOSXf9uGZnL3N4skNbdFwgtqCx7HDOhCnEGFjy6Rr2Axz947jX78ilIdHLj
Z15jUwbds5QWHqRyQfJGwU6V2NrDsjDBerzpi5psSwOO87d6fZQCByH10zlZUE7Z3sBRovoOJv34
u7/j7HztI5J3yqMl/XUBQo2DoNcwGPX5FpJ0edIR8RPLoBKGNMA4+Hg0b1Ge9EarNHG1FEy33yiH
rDrMTqkB9t3CwgpR/pnZHTezXeVork0JpxTYJIA8CXbgpHU76WcWXO4+tfp1q9nVJULH3WzFEzta
0RPsa+vZ2QaeFVQneU3IbvNpe+y9qIqqcK2K1pg1T6VXmoikLMWQQylJ7RI3+mx5+XgmSBQEnABf
UVpHmuaydqoqXErlNSGd1Ly2ed2qSnwKEwKNhZBwU+pymACOOuX6XRyEwfg9PmJF2pPnF2m5/V8M
HNOzECHQIFq4F+d+jv6xNEMI3C8LYU/4o0oJY0/1THoIRKYW11xlO8Qrd9HAgJ4GWkL6PqwlBkpJ
OIKx75uSc0lvsrrIIPjrZDAsSRN5TL3WP0iHkVlERViJw3rHNswBiEBrL6gq6k8ZdeXy3XYREc+Y
OE45BzPdDO9AMNydlSC6oPc+N20IcIEcJpFEcSQ9E60aO/RC0wp7lvUpvHoyiqAaIX9Ar3wBf0rb
eGnRnb4neMzIxNJ9vmPlL+FazC4p1WR++OVaEVN3DzgROBgDUQmxxvVXhnh0cQZ7+x3qB4dG//uW
QsOOmm+ohgrTf1PDGR9aVwsViHHTVx2sUnje+DV/NapnrneadIsccKEfCWJM8jtHAUanSwLXSWD+
kmkylqfamHvOOlLisuMqr7wu/r0AxkNvc/yABNLpESVkGhnNu1nVvAdMb3c5m00hzUe4usTLh5Sv
qWbJwQN1lYcsEV6DjtbEfQTwL/gAnpVc2X2cNviymRRcGRwipHBGJAwcEDaWIWqiSSHiVmBs3hZc
BhCdrRYOR1GLN95LQLnu/CUP9+usUvcIrl9uUvx4uqAUbqmfnnohc4Q0iJyvUd7673/Oann2XqbG
WtdtzY72n5UgFel4dj2KuTeF/edtlK4DUzxUFbHTaJQW+tjlqbrw0DLJkOfK6W+kLqfzL02s09LM
7IBRzlE7uXcLhBhWYbEfQiSa5UW2H+1f+S3pJlcztkTpF6W7BMPqwEcXvBRXHcnohaCWv9Xn8tqf
723J5kPTUDqmYXh6mTpOczFlG9tdyTpbHfPvMOn0Awy9ZnW3ycf3gVl/8R1QfBwIqxpjBv93dBlw
bSLdKCP2Hf2Bstv0p8Bv6zGmyosSJbM6AxMkQCuFAD3iFHu9JdwvnJVLShYEEqQ4UXEVB/jr+TNT
NkBpHZyxPiIO9My7DswouWWaQDqFzhS65wy1Y8g9L5PPuRNxXICxCbIcinD2OoU44cLfWh/8Asm3
ilFMsh6hXAWumK47JzCPU8K98q1Ot44Mt4jhzHq2nZhKUwnX/zI+oMxBQ8cBh00zWA65lxj1WNrB
oU4n5PdL8cD61jfwMnuh9+Sg+018gr5HVRLdye20vfZK6qvmojeG7yvqTNqARsGmVrO4GusOrmG4
fiqVwYxyFwY7oUnVDgLS5TvuX6CzMUVlknfIARrBi5sWuXDp7GHC56aTPuaSgyw8trj/h+H69Bp5
cXGSsp74NUVrpIbYtXr2nnfZyX/BtTisoDCAmWFVMUl7JtZEiRLdMZqbVQlFn/APyuaPviq8+URS
dsOH4AuQoWcRFqJNS2A+oJ5o4t4VTWDV0MdJJT+YlnFPZsGicB24dxX0LAtbfhL1W2qQNohgpq1p
UF8qEdTG1WP2LhLZO1nFvDMW7biO+R+uFA6ZnQZO3dO+2+MiLn8MR1AIBuI860uiB2EIBXf9uQXb
lymMxGRJSCepFoZm6fymR7ryCZnN2IpfXSd61SdCYTtfiyGjpF8JLzNKVa0CrrJ9NzSiuuLZn+6H
nhxmiGwzn43mal8Z46tr0O1dqNxCnIVln/KyCcx3SzjpFMOQ0s+Os8LyoHWJpct0KK+/nznwP51a
/JzmQLXsnuXxLPptHCZwNRGTb96v0o2uGL+VF649PBsL1Bu4BZf/SPZtaaTGNQjk3ritCK07UBYf
hRRvV/ozBHN5jvyUkUxPQswKUYwKQk+zV8jmEkHRIEXJoNQUzsJtVoaqYDllrAzuAp6LzmThAD6z
me3GpbtpfEpMvjxMFVKE1ympkJx9zEei523L0Hz5gAxIDo6XwqK0UlST+yW/6IOGq3sMKImoRAlH
hJhV4ZaEQEJc/uNXHv8Y8wW7nMGri2QNB+tA2touN4obaPsAxyg34vfx+Wh5POjF9jBQlTY1vZtP
Ib4P8aY4nf9qW7Ef51XtS35p2GsAvbX7SvvwESByGbIK8bZ6ie5JHlksmyHoarJ7Z0JGOsW3dt8I
uRvupAwR2WSTaFBz7QuH5RI+LqJPfTiTaWy/desJU7gNN157y9Gu6leSRNBSkmElDexrtFQkyTgD
o9+7EetNJks94NQbaBHHJTB4HN1LIq6gagQngVIWUrLwBGf0/YDI4P4wohOcP1rtThFguudmS0wQ
XIO3fTCL0DnmRkHEegTW3z/syq6ZU/OZki3sgFKnwjvDJJ/iNELKjC4ANLkrGieW1pb0sN1uGKBJ
bNsdgTgzva68Rf6hgiBuX22CowNH2u+IL+3kie3venzYNWoWkkX7nZuhhAtApUKh4BcK2BSyezax
cCG9dQiWix3A/OdYD9RIie7lEHxRuarQeefWHHD3IY6CzCvga3Hr6DyxZp1rqdVoHZVcb7vejmFE
9dnj9JPgdrOzDGuZOuJLzR6Jh8dpv4eqX5jtNMOE334F1i7FxxHte61Jf5o1AHNqMbrHK4owzcKF
a2N2HpOBqh+wja2XSH1ayWgmbDAYgXA4SzBnXb5eWaiyI4waDltXWW+U9dQ0sYSyCfYtDLVwextZ
IbQJHFKFfR+AGC63ZzAhI8Aa73uxuga/wYP9RA+ZElevSVprT671rY66G1YIKMOHySSKXjNabsfR
SLNllazwD3sVP8YjgyMn5EUTCpWmnmgLJqSLf5EDu2xnt71LbsaR0VNzh3MWxCj/9QYvTO04y0LD
lPGTaxKKWKkYW8VkTZR3WAJgWEWpg+DIcEsngakOtWiqLc61E+BcxdtB2FU5RK/ifph/2tJ60r3I
afPc1jrcg4gvxn2mXkJb1eyTVLgmM1vV1/KRrvkUSrdlVOPPI/jQhefsqeNg5mcThHu20BbC0W0e
PC8DrkhT6d6Q8fbMRtW08bE+8Qcc2tGmW5R4xwiNugTEAgxeuWQyDMLD9eX2+111XeUb7W3r+aTr
lezFJGNUHofUqgR6LR5SWv3dIngmhsYVwzyHD9eqpdBPpMI3OIcPh4TrbCzZ+eFfZ7ZC0Dw6HdYO
oCPcpP62s0FB2dfdTzziazLYRfWtC85QXNMjoa3Z+au86KnvIyZJeP+T1P8heoSP6jczBXHCk+TL
EUGj0WzAwPoOxXTIyA24fwr6SpxofP3jybyeh9inYCblOFQ/1ZFU7rPuZAM/gp04PSrwJDsl24Vi
B4/u8k1kgKEzOBo06w40RYxdPTZ1qqPLfrISrfzKwy0cExH6jeKjbN9OZt5innkVAfji4cm3cGd8
b0Pq7JEulbQe4+X+Nk7Ax4jUOYXcHc07dHptBj10IPmP4AlEdRwbrAu5ROcYj5ctZAXXLIzUIhhm
capW6+ATkjeioKHMjPymVIXhvFNrGsKZrM6LVkgsQ/Y/TDpeFM93ClwPCb7w4NHRZ5PrhfCz6/27
MDFrYd0o3HAZx/VgE6Y4X3U9YUrfimcnH3np3fS3/cOLe/IG1qGb1NyvgW4vpmBTCWU0vQeEQcUI
1nXB0BuifnB11JvlIiEsplqZXEnSx5gvXl17GFYS9B92mM+3nYVUwwOzPzqfjA5iDrJ0z8CwogV5
UifFQ8hS/4UET41HAw2S2B9uL/YuCe+LQOQfeGn5pPRsZkyYUC3pjGhOXkW1BreNW0w179AlEx5b
Ioh3xMrSVQRrVfYDrgz7nqcwEOPKJZiKLcfOHajQ64k+JLlnVqVYXjUd2b0UrZm4KdyDmR9UBnX7
N2wtwNKPbqLuH6eMhCmBfTvRPyUsVArTRNldjF3HeVxK0jgcZWCxsErkzHklz/Xwf+JFFeACMf9P
Prc0ASV4SRPfFsqWl7cHnVTYh0/ldnxEwrSTUS7OJLnWGZ58lwBYeD641nyA9VTIpNhQ8BdorK8y
73h+PQRJ8KsdLI0fpBsXE0haQm4FyGP9DtRig9wSaWw+NS21rqzUpHpRjVLZ4OmyVfeWEEwH1sKA
TH+7Ezd4jM9PWV/3dTM06050FICTvV3Lk6vqSUA3399j4WlvNp1k5zMrk47ta4vFgQXp+UiivMZi
NLW1jgh1PakcjwnVHtG5s4eG6EwVG/AGvpJzpoNZ3ZgHeoQ/x3+0PHWHTmvL0aBYaPCuDu8E4vTR
qrVOQwwsjn292QnydY2lx4eNH6jUnufzwf/6jVhjgBon1Jqy/CBM3f3hg6RrECY1JZLb4qOx3iMn
QJyDVEGNG3wYIx3V3t46xLZE0DPMG+N94oPhSSD+yJ4aAVpPZX6u0Q5uqNt24D4kg3haFTM5LQ5C
3f5qx4EfpNedmcf9wyVUJrtV6f8Ab1GpNuIAJ2VCGURgrbC2LS1nXPCg2cJt3vPWh7togsabXOeD
gllM64gzRnmNhteMO5xzjzCI2IUedzzm7vCJyYXMFo7XI8igbjQOFhiUNCN5RAJ4hc/2TGOhqEGf
qht/n+8wjW00bZbCzpzgF/NDIbVv2gFOtlhNN3fG/suE/BGfqT4If5Tf78n8+Xh8z0/HF3NxPNjs
3HeoyosWPj4LrHSScyXWhOv8aRLQRLBDOPWbx224GxXZkyVrnLh3zrOTjOeVY3rjDlgMMZ2QJx3G
wSwpePYL5iFhhi6UHgj82WY9H3+6nWBGsHvtD96bbdXQbNHOI0UYJ0YV1oOow9KeVcT84w+nPEz3
oIKetS1ckb0aeazT7685GwG0B9TA4pwc+Hhn3/01HAiWNFj/ardIc3neZ6P8I0ZJuc+3GYOdPb2g
WR2mqEsQKkJbCFrXr90UbrKLMXBKFjKiENNWECknuH/Kl+I4hb2spb7a/dugKFeDzxXvzKPRTfwC
BjtbHccs1yFJ4BbvDj2lud9+U1+rcnWGS2VNf3/puJa3wkUWz1Hd0e90BXK+ndHgWglCHRD/Rgnq
7DjC+EKO4qH+b6B+0NYBVEBJStaKQvTeityXNm46cupq9CaCM9/kq/pairF7wnjJCUKyNQFiLWy5
j0eOgJ1i9QIr2TrpcfEayUG4IbJR5o+TTjdGzmi2hrmT1yNJSScJ7bJqxRWzy2eEF1t3wSifn8NF
dd6HPvDBWWp6kpL86zotONzUyQYTuxhKKtNQDcGukFSZICdLoDOw4e01XCmUjZTrnYcEbERWk5yH
V2EqNQT3TVPrMpH/f/sDzsa3kF7yTQH0tr8R5MgZUZ2b8Yy8UqCeAvPLG7Qg7fPXinJ5/KWvFbUM
fDIVDf5ad3rnl0FRMFzkNQSVy6i4kNBzS3nfGzlrM8Zm19DXPmba85aBJmqK4fB+09KMSNmT4lbm
yJznsrOU3dAMaWkyrB8Bfqonlfh06ccCNkXFEclhiqVr9efgeXYjMWZDvav2QJuGYpSg7BBGPH++
mzJ/BXDYF9+onM/AbeyP1C1C+ljoUZNhepoKj2Yc0xf9YrCvgqkhiyLAq/qbsAfLQh5BljpeQNVe
AyFEHXd8LTjvUMQLJy+/kczeCcvKed1zXQndTTGWpYV1BP5p07SgWolKyu5VEYO+hp2qfGt3ZyS0
Co/i0BYviUoRSNkugEyHq8yxiFKMxWqZ/zs8aD1ZVRpWUyPK0eqf7nwXJkhxYwTl7ywIgyz+xK7X
VGSLA/tNVAG3AUyLW9gHu2cvXKd/UxXqm8aKNgg5WjM7iOxg3C/QyYcPUI/qtwxHBHFTtROZ4VJq
RsQ8sEd3C9HdQBJEemhL0MCXOhuP2ZnrjvQOKobeiypD9Nuau7InUa38/mKc1/TFh5MbptFjRLKn
T4jAfa0XA17gfmsSatUAK1LCNelcXHktQ8UcQYLywWn6umtuIS78Vavp6pMfv5bvkCU6hX42WhZd
ZfvEKAW5+w79YjNeyw6Hv8O+2FUfaTo0s8ADqyf2jWzjY18XkqWyiY1gqNSTUoHoIGZ4/aKb97wJ
kQMN77YgRnCie95TVIrxEvgSlR2qUxsDLIn8SfLR0IojxK+OnW/SLkfroXdtVnnTGpXVrymWDrkA
Y5xXaa7CSlh6Bmq8MeYjVrewpOfU/R4FC3KNHMphqJhUQgmoJSZFNVW1Ja+2HasxmE7H7iqB3f5t
hLc1ST3OgeLF73akDkr3v7Tjs9gieAOtAO8GlalPghGocgY7M8HpocBksVhQ9w+xf7lTfO3Qlgu3
LTrFhrw0UKfHtWCRbmwbmPRSTj56i4dMUXNo/0dMy3yly2q2AmcyCqU0cmgiBYMJ7dAg0jNjTRF5
oyrrcjpNyUchPsrj1ElKBFXZgNAVcVeYVx+cRLIhUfAiOxUEc7pN4oNLFA3qVF2muayvmNy7Tx6j
igXn3q+qCXMWKRoBUU9joJ3AfbSH875usEj4xr4BewrDVRFTDp+krXR68UHyG+iXVytYynLsnA4z
ywywAyzkJZTjt4qAyf9yT17X/7uFbpYqI2Op3AjomfAdoFeJZXnEjlsnOjq1R5uL/wAIM9Z/CBsh
4V8fkD+c06sHvkSBD0NJKvwCGe1CD8iZcglny1JhIDcoP7W5yg3NEYCggqXG/Fb3JKpJVClZfwsj
PLjXSXVLXNe7rVfkqftCj/ApMO3UY1TrG5b9L2cRr4FqBE+YpKiQ4cHFLgGgyD1yin7FTZV2gYvS
nUssTkkzYOOcu00YHIjd+dRTSN8KxycofNsG/d6+Wa8BCN4+/7k9WJDQQDqUbfBAGSn9fgVQH/g7
PTspbOg05332lWhuTGsnIhMRNDyS3P3oMyVyU3c/Ig2GFGHJuPVUXeXMm4i0LMuoSliUzAWhsDwE
Fxtu6iFHJ610u/Zdk8E3FkVP2H2Y+nuaVyX/yUdXPRAenb3eDVJcubzP1B3QcQFmCmhQ27Qk9XUQ
8z5lGwwauXEpaBFdBgSkzCbbiQThsv8BMCeFcMei/Kz3X38ZyXLFcr3U7S+YzlN1X7d+Gbw+gid3
jqMlteJC2jLF+QKVRVoMtksddvZjV6d/DsxLdehfjGpmxUIowruZNE5kASZ8sjj6DnbsgZe9/Trd
Y7juQwW1VsfPwrv0/BCsfQOqMwe70WfS+JukuaKd95zbi3awyctMltjJH9Xe0PDB+vk3Z4xTGaiU
Zf5ux2rEDRQharz1V/IfP70jzBBGUFVcnwAuejyMSXglNcq9lXgUK7ayeIS+ey234lf3/j0YBKxY
Dvi+/MFJ0IuBnGva+tPw74U3jOb2UJlrqVky7VwZQiqD6JPBZQosqNnhpgLZpf/tk7HWo2F4ekw3
vCd13CU+YpXPEFzSv/MOLF29QOXYqv6emfUn/73BMRwXmNmkA31DnAbez2v2sbu9/BgE2YukA+vw
HB3cg+yn1uxP/QRQo2Eyfo//vE14HGmymmP6PqmCpawp9XEAHaCX8P4WQYZ9TibcoZndzvUYZzsd
BSNrTqWfmwbjwwMDc+hwcjskoVE7cibglNhxJ0zPq0qf88HCnMs2LBJMXJ1WJMK75MyejJ6Zsta0
OTRLFDno7oqTA0oBGf2jk0aljlOicrQ7jkJRL3JLerF1esvWWUIHbuENG8gxZz6ApQtb8dHP+YtG
Qp0qcjvHxHmOz+ppitwA4AocUDC+W6n/j1/w6lV6BCXXtuSxOGN3WfwaYIBDRduMeBCkwTEInsqF
Qc37QpukQvcfc7XugpiOozswInehr6DJOVvw81K2VEgFx/lXeqOA+j4T/588jLX+y7iim8Uj4uPg
a8ZpoLbaLQSRu3N9gSQRWG5zKRwr1VZt28guPuLU332MHMqdm4UhGyitWZGiWcbWZAq0p7CHzK21
QXLMxmMHXCuPracXW4Sl6EmyoBGY9Jgkk34V58t93Zfjc6DO3BaStj8Djtc+uoGdEZogrma7AR2z
aAbWsEnMjTQFp7G4YVh9sQTaza0zMsPP3OrIYTuvg0vaMULKCQ4WdqapwydDqeUT4NY01aiwcwTF
D5cFwh9xaGUES6oa1OtA4v7igLbrXo5aEVJMCoE+rsrSM6m0vDtEL/xqb8/pSgevASoxCV4I4i9u
bI61chIyfHkDrnNb4zlZJCKxlpxrEVYZyAgFXwBTgzgKjV7T4RsGoynbFvC+QCFN1qQp7i6yzCNj
71yrcdJO8xcWM283nibVFC28h+cAsXYbgCoeQ/Sgxs9Pg6RpP84keJnMeXTqwbbo46JsgCUUJbs5
yLcrH4liWl6u8WjDJerHyJaspgbnu2/eWv8AVonLLIaMjQwzzy0hfp7iCg0qJGUdtScCvB/mZF96
etPVMWG3DNcn/TvJ2297MVRJFvt9Z8Kz6S8GECypzvvKxt/HXXComfccIYQdHmVzgXGjHiqoNfp2
jtloPzwIT+Z+VxafNZsfhAjJ+ophxcleeVZBjUZKUZgZSPZx8Qp+zKO5uuqk7B6/L/lN/SNduPcU
sfvp8kk0VaEoiroodDc45nHoZu8sQEa3edCqfBZmIUQNXKF49Np5ox49rr832PZMiOyzGjCjjucu
OLfQ+AfRoYS/L/zlFX3WpC2EFf1WqqLVXrjxj0BhbLKVyq/0JagbLh8Zgq1yI/zUQ5fxJiecQdli
+HoWOA2IMsdbeJGDQOfUqlIGY1ZU2TVhHpIC6Am2yB1YMUE2AH8jpnr+IOMEcvudiwhaL8NZbj3R
t7AcW7fiMiRHQgNoDZHF7Qd3hwJWHH7B4Tn+Zfzq7WIrP3xqfJD1rPcBiAl73hlsWDUqY1hcRX+i
NT1JCAXC0I/cUAHKHIq+09GjK3l1kWHKPeuUWmatRx4H6U87PVzwAK8L3wn2E8oJYmj3rG34UwBA
9IEYRJ0XYQM6kwTYwEu/oZlU/FiLpj/CJaIlwpGbQYdcf2fsHszmQn4/1aTrgEy9yBr0orZPgvsq
ziLdRe5jinvgH/QDtJjgVNiU23DeOJ5Nt2J8UjaTxHANLUv2k4sk1XLVQUy3O4PsDniIwk+oFFre
qoqF/zT3JqRZbUKTwEOrJsX2E3cpqriCKqfB+FsZ5NVeaMx85IroCyW5PLqyn7QQGTyB4bSeZjdo
FmTCXpxkEUQQCeWcgkCJCh8qrYZ6ksxxkI9Z7QinM1914l9QXXrEShc194i8hMZiOHvzbCrG0qpv
ZEkCwJnzkQbctJGaZpZMTm8SmzbnEZYrVzwiu70+CG2MD8pvuK/sSeR1++rz+j5pyOcWv4zbOZRK
nadhNOxOkiH1s5yTplBI+cET4yHNC/HsdFu65KwJ8LoQnqvcOAY/bBX6ep8J8AGXUT1JmomVHvKr
V/VZwqZBe37v5Fc7lAaOg01vlEHzUClyFWQtD1KiIBNvyjz4m6ji0TzD4xx505Sj1sfnOpKkgMQD
vtprZscRdl4Bq4EuF66mpf7N2nWMNfgzA5PSa1xx528x4FDkpb2L8QgZqXrfiOrjFPVNdXUWUkzv
LL39jpg6MVYj1fl3KKCNYGzeoX1APj0/daZEV2WRaxBahFL1jAzdQZGO91ILxLbBIdAIk8/FHU2d
Ockq09fVkzLPSZAKm5ouI4i40Nb6O2UZQbfX3B6ydlJb7h0EKeCIxaUZ9sYWON+4H99DV/vvh2mk
EBuw9jek+UBF7q8tEFpOokvaS+pmV39RRcD0OK1+xFlhbDEw37nrE+kLK2qDmuOJEyXBnEPOw/mV
TFHs7xeOliRxNI5lHPEaoAe9YyCosoggcKEDDpK3nQI8LtbwuyU7SjW0e6PcYa5P9u+uYOK9fiA+
stnLmpdbdCCn0gRWWxYfLc5bi17wpJ+nU3zCRE4rtvkjr9BEXzCPoHmIoqnlafH828Yfq2o5SIJi
zVFGuEkgKTFBR2Pt123Jsze7ZwwwM7CFBKGJM9ZhXt0KBECVmwF81jYoFZ5k3yxTXGJ+u+h5Oqc8
rXJQMAM7wY7f7UIZjyTtcutctkDIR26Ahj75JjQbVAO/Rbd6FYZI2eTX//lOWL67AxLBzhC+l7CY
g7KWefA9nTbwYRKp2i2cfYBPXLh++g08Oy780YQS13sbQfnQNWZteUlljNoBjJrlrtCvIHoV88RR
gNHcMWENlHob8YwbUqHylPGv1bQ06NdAhA7gPtV3pD/YKO1w/z4xHlndoAdDpH3eBLE5JVqgqkKv
O2wFFjC8mXcA53YMAIMzqy8vi2CE+9aWq61iN8olQ67WqxJUVmjj+bUlc/oEhu7pbwG5aDUfzKG0
QOwvL1Mk8Pwof7B+gZ06ZqOR79eyzvU7i/m8y/jHOUn7DL8b1j8IKT+WCCueDy6QeN9XLBXYRAzK
o3wtPCbyotReVvxx8D1TLcjEFWu0BYWnHd3Ii+A9KqDYLnIPgp+5VMbktoeQZgweiBrqic39WQIN
8/QQpbOb0N0BaVpFr9Dzw+6BPaJPyz5fYhiM2otgk2JApkusgi57n5Z4ZWcpA/BEs6hOaU5v0yWz
NW0RyFENH4Uv54fdvZhVa6IhoDk83oTb5Fu0yygjYZDAHKGQyeQKdvKFMlzlpTwiPl5S22O8hMVq
syyENzNyWxWzdq++nJK/qctpk9TXWMerahYHulB1+yWvXEmP7nsUfXtaCCNqoYfx6ZyKZJdlK8Lz
NDSr6wN/X6PSM2f01pWHEBOoHKzlddgmfxSevgSdcZCeXkuISS75V71rq5o5Ok6W0iEpzXyUCMU1
FOvAMXRS+O0o2VFgAIaPIzlBCTG1LAy3jJiDJAGZEVAGBS1M8grSjYLlxzl5irUxmwJtdwspKUKG
0KujiTzPHD3karkQQxsTL4eziNH9Pda+pLYLrp+XJnwmjLczdWg2qwGrWEeJfMZD4nl8nnEJSsXi
shhLPVAh6WSBPJUJWMs/7cwc6RBUrYRV6PIBoriLOI17a1qKmg0XCE8w6+iBIlSztg20vIaHL2I3
pS3H0/NBRD1AIAkDsU+xm0yyasJW6Jn5BRAN+FJQtvilkDAe6mVBcJ/Be/7/ofsG2EZHaVtLWBuP
1IQ1ancZLlaXPgxwgAx628IsRhERe7k7FZ/gvyXb5HL59x4LckrMKU3Z33/Kv3nnBsXDO5h4ADy0
YMJTssVNju+Ztg9a//V07+qErx6uXXNQCseYXOgi26oUyBmge8dc0O1KllRqyM6MtYgbe/KaFkdI
BpldAWHqsHJ3Zq6Ow1ypeNRQVVre1vU/66i+WsRDEkVrX+UhZ7Hup25ubMDyNRXXW2QeT1wKmcgT
QsI/QdgY4LaWpRbDLc/wRrs/22PrThw5soBw/zmfz1UvPaTcMgHvI0O+/MWkIB/hEueI7NxtS8ta
4/ECvf7N9hfyRB2LEYX2yth1o3mWs+l0xNT1IiOjZKySWR9DWeoajAz3TKioUJo/Wh23Fr2gq4Hd
TeF+7P6JaszK4SC588dE2PdJEQ+Lrrwmaox3ja3XYjkjlI48C04yDdGUENiA9y3qC1GBfn5AWAQT
+gdY4PGrAs2KBX/a++h75gLzd/dqBIDJ/GqfSAaZFLbtvx3gAwiIe/PZmSAWNLB4mPtX8/yHbjWW
O55RQmPc0nlEeu2fsE5iDj8FiqvMpQxp5z9sBV7L/JWgPdlNHyXa+A9SuS5x2itqliUoBuNWxXml
iPbpFBUY+cpi8htHnpN9QWaby8CgcGnJAFk5t35H1qAm5xQTqTPOb1F/PhlXW6rMMrvYpdz+mtJW
tveK3Mw4H76lgBy6NpHHAWntHr56PAYl3I7oscWymzDYR/MF02ZQXkYpckBcCImGz+kTQrYGCFa3
Bnt7xax1jNbSLYYqCJGLcV6F4sX/bn6E9RJXBoQGdFa3J1o5Yo7ZmsAmIuPP/mglLS9qbcLz3NEd
xTBYxY0AnypMRinUFBXK8NZBs6Cl45heOqzdDDjYBkT/qomLtchdAO9NQSSkvJ7W6EQ0CVrcRyCY
XzYvIf7gl7Dvpq9cWTCLypiyB//1vO9DWp0F7HVqmUxuOgUY5lrONVcLj1V+P/xR7T1sPTqzkz0y
+aw+kGBEDgoe9kIu3DvMp8mt7WsFCQPBd6YuE2gPKAVCevltF3KdwJ1MtviHzTF4Qf5D/1lsO7GQ
FMmx8By9f9FOKdGJjcxzeK1WvJwIcZ0a07jXzLpoSyH1N7kmEWx4Z6GTDfvTwE7Unju/aosdXdab
hHqZtBxIsyC4uM6GAj1pCJtO1Yg560OoRYu9ahR85MHaOqD8I9GmiU4P5a5ZeImTG7XUagHQ0N6N
n4Sqr5JTLRo84yTLN8kvK9aNaQPJ6AI6F2t56Ilni8KAm6F498JH1sUJOaPRr2tXHu8ct7A3PRkm
/xOYUf93xtwykigtkMvHeinREMYaPr1B29rXDi06me5NHa7gjMLkjjgOcNlGxiGU0o+TFkJHTk/M
PRt54ZX0FtE1aO0XP2m7wVYMKBluB0ZD/hQVxJtpYR6XSPyIayfaU1jVwc+Siw8DGOsoh04rNqpm
SSSNJWPVRJ5JUlfYMpbhdoIvckQNYEYhadMZhTebkHk4ZEsfTezAiW2aZRNek/IApfYwyO8BfAtj
xWFQY5Uw439rQoyg3jJ49EeOiWqUpbecK2SubhMTuFylkuzWgVch1EtKKDRJOIdfWZdTlP5CLy+K
em6Xi8zCxtrfDLBeW52zHiMi6/B3t6q9xiWdXe376Z6IPVSiEsG+gFm9wGZVWJaTD0g24ilDgFzK
MUCdjrizK8tbY6CbDNC+XVyH3pSM6hZ6LDlal5EaqlvlygIqK1uydGubR3lnSos3p4Cv3Dit73g5
s4Oziap3Lv8FSsRlAmG53sDn5bgOCuTqSBGK3bFfrZFD0ueV/HjuvJMM6NG2ysn83l0PYKwGyoZk
kU4C9uBtbhVbiNGMgy/RWAEpt1mqkT6Z1OeWsm08rDA8SpV+wZOC1DC6b0sICu7A/wVbdBcOsVHB
EZmmr5nLduFrp+1rUEf6WHITWztB0TwlTtBLbteFP9AJlcfmUezJslVTqkmOvXb9rDzoRRHuJ5Ie
URu7ZH4LIsLvNEdEg4lSfnQqm5hWojrXJIM4IrV8nzHtBJYwz0O4T2vz4LYVjq8vx9mr4+BM7gpJ
yYFQwWzYiMM4A70o3O3yt4cfzK40b9Uf9WAvHDtr3RnItIGXlEV3w08suqXXfJrR98RxPMQfewgd
RZT/Ijq9E2urYDpiFbLuKoVIqSXlMlffD5mxyMYKI/0duW02MSRLEiGG4BrDcEvLBUQddOJdbg8M
pjzQJRB93485eBaK4PUjOf78RW8zsPvX5aJAjcIHypNquDQZ9gYSW0gRXXUzLd6uVTWXKuVxc79B
8GnktcvgQK8tTNFhXn/Mg/xtE8hpXjeS1zwtQYthGe1bzIvNiMQ2Ltdt1p65i8R/Rt5BypGBM7ne
xf2IHWFmQb6JFHea3mJ5oPv1rSyXZ4Juuue66DFkafLvG8nBia+ww0fK74gp5KufWQ+3vpYrwsln
+Mpsq3MSISxgPeMptWPymhnyJLDW1XYohepQjqTeDbAs5LgDn+cZoH0Ee0xBsrQOUJ0fh1ujZbR2
MiAjEg9So11hG0iWZa5ciqZn22kHrGOmy8/nIqxLPEFjjsXlWHVeAzeQ60BFOIKOmpz0LaQw8YoD
akDcNR9j8Gtzda/0dnDsAYmF18TOSmw40Yr37mj8fUErlZjIqmuGKEezy5Qv6DhRGsB90JpoJWgp
mHn59O0QsLrB6yuMUKv5W98RPpjxRqKINUJNMGD4QQcv6HrqLS++Qos+eHP/mr0W8zeKbSKiWCgh
PYN1WgCKeGh8FByyUOUthxU5UY70DrLeac82FGDe2cD+XX21Tlc77Tf4RaznHm0cVWiYVy3TPOIj
aCydbk0f24scNoDDlXgFsphMs0aH2LNfkRcrZIotYMJtdQbDmpPzMPO60Bk5y5HVYSNtAf7soK+U
dSeg1VF8DjgQhHxzaMm2I0GK9VaGW0zOybtkYdukbevjCpi450faJzjZKjJluw+BY06dPiOFrx6p
eAxAuR15FTi9JWuBUQgRERE/qs/n+3Tf/iZKZA5HHBW8H+wytMj3+S6VZ5w8YqMwhLTiTjCRLqFX
KS43NUriuODtwOxKmhA0ERRehbXYswuS7ZSs2SihUg6CFZOCd8WCQVqMLhiVGvl/whAgh/GMyPPL
6Iq0I+JLCkuY/PWq2ScigGqdZnJixe9EIzt9TRibrKbIYfaEiMsmuoO3wyUCVExyk71k3Cpg41s8
Re+MEHB7bLeTk+nl362V+uP7Vca7sKj2QHQHL3XER4Vykb3tcmMZtBI0CdxxddNDMXocfyy++hv2
Ay8adjhqohlwlP0yH8SLMS4wEqeHrhfq9eThih/PohyO17F9DDOO6NwFq73OaAUgN/j3u9HwBABX
chGd21Fg9WhyVpXkz8yZCqpPCiDpHGy4SvKkkl23+RoEdLVFdic4L84uHefR851Rdj10drNp7t4l
Rs8s26Zqh9ZsXzk8fWhkQ/9RIYZ71PYyjAS5pm1mSfD8QVNRnziQkTv6noYWoAfVXheGW58L8U+d
gjYc4fMDN6l39RDIBAzVQCKg/xvXWYv4DvFuDb+GhaCw1ZA1GZI5CivHaiDi4vIUBDvbEgfplaVH
TpyUtBXNjPuUKaWWogidi27hXSxCs+pWvt3CI7qZFdiqKxlq+EyNx8jUuS+WLznec7tv4J9vuHJU
M03h9LV1SJrWiP9AvOQpUzTcVvqTd4GCZfOeeNryX7sXaNtmDSKExrx76zkWDd1+x5RGomlDNyfe
rwiww6sNz742ze2gZAJmsQkY7+Hxg0scDiunrzf9k4351eWDBjUkqp6U5FvFjacjO/LeiDCgnKMh
s7l7GEcDtmwhDwvlBcvvf73dC/UYxBdvzVkid0FWkohlBzCvyXmaQ3oV9SYdIzwx0Wt5sZe1vpLq
MuiYOQ0a12kY1k9tcsC9vYJWP4leA3/6ndr67ubp/em7kcZ3LOjqHMp1tFAE3+gAnwnieFjfcK48
rvpVrceCEBJ5jGtMfhaUBzTgAHjlpyNqmgaxigocHWgHDc1fHsmosGMStpbEmGuF2eSig3KIGtgy
Bg082MNcK4y2dNsWsFhdswd0cfyI6FOl7OrIUqFSvocluNF8dsErU+ZFVoD2tx4bp+tP14s2hSwX
8hBZI1iGzgYU8z9HBTOXiM1OLAMilhYt0H6omy159Ubfy1c1kNYYewPx56zGRn8afHM4U2XauVRs
4e6KZlXiT+xlNZ1P/K3aVqDGdxPMj7XYzyIlImc1iNXTxbTv3vKN9G27foJ6e8xXvUsM3QZ5/79G
ldLXpjBG8Q2bw7bwGN6tksWg4NvpIqGcnrRnENPlTOb826EikATsEP0ZUV3so6tC8N2VwAuUjV1n
0cMHgOumDzYlVXGbhtgCMFgvYf+Ysl2B413fBVUuji24Rmt4u6SXz/OK3zmYrGe/NxMk8zTuddBy
NPQBw5JmQKTEEYWSqxEclxyUHjh3w7Wf/ISuouS706RdO7zLZikey/XtkmpujvhuZiYAW4RAQJ32
/qGuRV7Fhtk/fa52q+GV9cvtih903ZtNrxr4DV1lfQGyjSVuVOZSSNkti8Ey7UWPbNDC5vbEEULj
7kRHqSbGTByX+GC9epGH/jz9jnGgZr4Sd5t5fumInzPPmYgSPKjGOlwbY+n+CIrHBDD4EbRQ5wIm
8RW3nOTqEmv2gUWIeo9Hh5NTBaFpYf6XUwuFQXieeFPGnZL0QG/UG8V/ev87Zw8gA1Uig/aoTN2a
eW3L86YuVKcUTuesVGfTMAM14cgsPQrSEP05hGRH5whDIesVnjke5ie8uqKVXBnDV2awgS1NGK/B
P5fpOkw02h9GyT9U39uDzjn0ux2o0tbQvTCm8cDdV8n5tDge1CaoHXCM8CEGXg7ZBKAqDFPER+zz
cWQ6a53/XmGIwHGYom3V9LFi2B0002f4SycYXRXPzWF5VIS649UBvESMRQ0gFSdEb83VEGF6frMN
k+8MJrhxq8k7ZGOyEL5bv7XtZKMaKGPNOJrttymiTedLvBRnhqEP6QXIcU5NLMuaKvePy9dI//Ui
RLzjyC51J53E9KmRYLy4GEkkjOxE2/iaQVhh7qRtZvyF5d+Nz5n9j0jmRLxvhhkv8aFAcGkfiUfL
k4x99nMJKpfvyrMv9yfjzc+J8yTEAqBGu4VPU2cNwrkMbzC4+r3UU/h1wVm6MH/TMCep5IxSYP0s
3rqTIigwJhWg+VYh+Jkz01QNh7gbuIyE8LIzMRPt18hxSsCuZvSg984/4FomCflxOJDUeKNzm9az
FGDa9mG8d952cYsF+6V6nPzSBng32574kEcCZmyDBix6f6mw8eXUy1RFqhIuKQTr5vfgNQCezDUM
Opcg6VFRqhxiCVRE98BlcqHgbuZh3JzFnFTHGxENythyDHWX+Z2Va/t8IfBOTad6MzUT99oKD5LY
+SSPHe3gw+LTSjufDuhrd7tQiD/TegAhbLrQWAsLE9uCMSF+fxNljG5j+NtVJ//lT9JGcuCpOoAz
kvm/tedF9J0yWJCJn1N/E7o4tDUD3duWAlYSTPTYW5zmglWvJBwDCJyBIE7OyY83KPrIUtoS7yuB
WOBMORv7bA6H44t3aV2dCzG2HYKY2q+QKvFdtGZ3SWgmw4qvJW4z2+54RIZPh8h/DGnLKbyJbeh8
wANuOG29SYMSZFGpPObD4OZvRedOZmw7q7McRun7vu6Aw2aFUPudWfFTqCvQtc4YGsx5HCP5rmNj
uJN2LAjir8d77CaBpqGUgSf12rEPGls9yEINoCdMJtuUNkx7/FU7SAzVD17cfc9QqiSkmxBMiT7U
Kh4byTn3LXUBHDiittU0PzqwpMP9T9uYjkMSNkO2qV+jhdwixatR9XMGnTaWlz5nZjs2v2BUFxy1
GU0HC2DEJ8bU5+3Nh7tzeFZlbbBSeSWpleINXoPiumxauQ/PUDCElOtaRDoXVmVsw/604k3veSSm
HGXirRJj0QBbpSP2Fp3Vq4qAYHgn54F3mOutkJ+n1x26rpGkiOEqa5bVSk4rdeHCFGjp90ViL0ZX
h/yVlMPGOXLSe/h3gy9asPYUI7kDluur5aya+E3G/7xrBkgm0QSIS26GXLToaqixcXJ3DZX7nlit
6fqH9+jnTaUzaQBq8A46C4HkRO8NT0TzLjdI729o0zojgpkrQWv/ZmsgG7J6W2+stqlFX7/zS2Mn
x4RwrEszITKyIxQIhMBXXhslObqsWTTxqirsLKyIR0+rxSKZJ2AqhvppjxHEE0vQpjsG4JDqdh9O
QdJ9QST3FbNag+zoIIzzHAG3bAhAjPlJvVb+lDLJRpa4EPE/iBSXkTeQuN4KXM8WVXJsNm+HbOcT
/27+K1QbGZvyhiog25CJPHRz7ni09dKgCAitDzRIndFWUdRA6M1FMgCGIDbEzjnAWyskC0BLQSAZ
rqOOMt9301KOnaeh7RbPJBt3+LzHSZ/FtVnLbomJMCm4IG8xjyCJpGFQJFfnB8T9Ef/5tMI/om2T
kCjLgk+xx7ioHk3jIWY1Hr/TDsDs6a9LeO0YGtOx7N7c/IJtx6q13SUmnhLa6rnEJt7fSJ25vQiB
gXbnCRoHnaRrgnevRYanT1g/Gdx2iSXQ7QsWcMEQLRm1ojrykKI8g0ZMOUA2Rsz7gzmyCn2uo8+J
ck3duOo4nDwlb5WNXQHPjOoOn/8mW8yZrOHmhGzwn2r0lLCvaQuiJEmvV1BVTiORwa6Sq43eSg6o
mR74+35xDwBwzyJNBfWa1I1zeTX1H9D1D7LMItJnjQ95VRkJbiMrpQCYPr4ZNiOZtmpyv9tLr0Pt
I9tA7USbVzRXTLdmV7GFlWpSj4hYhMkU1oFZ4ouHOKmDLL1d4mgiwgtUdq0gpBuLnay8LWlNnkSi
JUtr8+hX1GjvMCnHGwTFYyK9u3DeSIYmlKa7gzmPlbAdGUG2L9gg0xxp5oLK+BnPTciRGnswIS6t
dQCnoY4Mi/X5dWNK2nd2bpFobFajGgtALpg9HO5OWE3rbPIJIxcvWQws2N/6JKWskLl3BUNbleaQ
ykWYPMVbEbJzIQksJcHx0EqwisSp3419Z+C6eDM6HqrHyp5/WWjqGRhT+QroPvFEPqx4dHqD1WjA
RFl3L6fNaQkF3V3Y8E8rj8jufNSdyYm0UVUpUbxFjXvT8/IZnFcf03X0NMlRXXtxw0Gt8n/ETwt6
0flRhofe4wu9LXYoU3DHII0KLf9ErmntNN9e2TyxnpLWSuv4GK/6yS931Q8Wt7qe2cyn5DfwKZgg
wpVioInshUUpL+X9T1rUdtR6SdXtbw1P7gU+s+hID6GtFl7TKhX9P4eKc8ZWFi4n9EF+AnNaiTZA
WcTcwAGTmvec46Loe5UHFaZo/67CzM3ahuoOu6B0CNaUpZKCPhzRGu8/MENXpFuejPyNbbXbfcYI
3AqfnnBPScquBXclPM+8LEuODwSc+xZydhuFN6UIIb1vCGUZm3eABb8kS3Rg2eU/U5Ho4aGWUZ9U
bHjxqxMno3zUOz/p9plwKInbn1qGdPRbZCsyZ1oufUfJQK2c0lO1GzHuNDm6tsoyVdUaLhtJX26+
EDODN4CoQlmCWdXJmj/o8mWmiAdpaxS0EAhCECb5v7pLtxnDlg9fH8MO7I7BmlYC77pJZmv+tgWh
VZkdtX5sghhw+of7eHxNlBhZP0ml0b4/KLH89KptsTh4WkXnm6jd+8p3d3YD0ct/nuMfs0ajA+fH
HgADY+QtcEfYimCzfDKnNgZqDKormKqXSBZeR7/RueF9Nc9iB7scG034UcsSIsCfubUSS+oMG73C
/oav+9DerzkZ6YZprQrqwoy4uK7xaYxSp4KRVXyuSpsRuobPXCmWYYmKFhV/348Ygu3mG9KYen5P
NI+gXID7+MI/hGpc1U7sjjGd5PtWahCvFCmAAw976hkblj7FjVrV2gEWfkYvlxxhSZvQtyWtO4KW
dPFdykQeMAcJF8+vDX5WOyX/xUSUG473AQklHMsKvZXlsjSIZmcD3EhM5B/R6/J3ChJlva0sXFfn
0VEe0ITnfyXIPKO1cNoFaz7RQdLLz7ligCR8CdZTtR7rpjvUjT9WLguXvGp1LClsYPnnOe8F7jaR
5Hr3x2JbQR9zDsGpfzl+7YhKNw6otRy8ZiqFFqth4vohCyR6mX3B/3/hn4+LfXhnXR2/PvcZdaSm
gJ7QH/c78JyoqxiMLWBP8jPsBX0Ki4neo086XvhWdWurWkGN0VZFQivs/J/ElOmvKUpgcnCt/FKD
K5pgV4uz/68sLAomby01ZJOddUFCtwFSu4zSuO54tPwBcBxZ3uZX9v6Vaa4hNsXZCFv+GZyGoXdv
wJI7TXeQX8ZF8vb84ibULYjHsPU6q3bP0WKOnqthbC4GSuK4jA2oYSgE61ifeAFxuvPcuDh8bksa
Tjumca0uBcO2hQ8Jj7HObbW9RRX5bePB26n79oIimHVmtPVeOAI+NbzYsFIflb8+ci7vulAE5DW9
LaITLZl/+RJsp2dBltXbYJ6SumzeJVMvfj/aFMf3abABS8L9OQwxha/6oqH/8/kKDS2NKpGd5YUD
kjzigNEOp96lTKsW5NWI1XG+bquWdEHbbwi8nMocn+q1Kilrw8Qaa+4CuCEmtGlClO3fABMvY1v+
TU7HwsYCYbRmxDM7l1WtZXNyJKnb+iS5w4NN6G2wsJt84xA2jlsjUTndN6WqDw9CN5SVB/M3JSGC
vggHFSRfnz9y7JqC93l2TfRM6gPvxIm9iHfVREcd4GaZpAKe+3orwJLs5xuZH3pfTns2sS9hSiai
uHjoVZiyokmjV7jouIyf+3XOf0iZEcs1LrQHBrSwYojwcfDKpU6jWq6g1l3itUU2HIjrKJBVm4q6
rWSVU5LYXux/zpLcn1Mt1LJLeTBjeUTQZ8bLubowv+t0OwFApBmaXzF13fzwpUNwDu/RHM00KfvW
BdlOmGxs1YVKecBPKZkoJ6ZXAdDRirqFAZy3noZjDBNzzsMB7Peoahs8RgX7/2fwugCAicMKc07c
KTgd6rW3xFPcldo+obFymkDb7EMU5zHxSpEXZUyfbdEgrntzbFr3WyKIXfqGVtPV9hTWmghOa2bB
TYC4PmQToDaFn768O/Ykunw3UoYH4O4k1HNG2QpypLFxjPeATuv0HjxadQVWhvaKQeKzb3QO5E54
FJpVuE/IoqwRZdmU3jiVevXhrlcu1sHEqpD8AnBSoT4y29qP6v2eBGX9iBWvsc+bJcCmNIwc4V6t
0o+lEKs+YeWcOm89lBre6tcDnA4ouF+ekxD4NtXlo0+Po+L69/iI3aONVIMPva10m/MhwuYz5XTj
JsLCuGQhgYnhjUREtfrIXVFAU2taTxIfRfGlhNpwQjgfuG5UOFFqkXmsvi9nm+0I7EUIsy/u+vmQ
VUKMcdws8qWWvwl0ZYlJFMcSyqLNPHoFGvB9egFQuSH82zH54EvdhjOL7CK90FUyq6W/H6TG2pgr
HI5uLz94nT8AMiu2CxSpc5ZTBKlIkNYyfY2g9FkkwjvsPWlsYXkjHDPMzo7zbFJYWAAYO5tGaAse
IG23UP6j1WFI9OR1Lq7YX/flNWcPG5wLIDX7gUQnU+cJ6jCaOhzx/8NpcL6ZxGeEjDt/upP92yEZ
/p7rIAcCx0mbUyIBzmrTTmMraZm1mfVGNzFV64DxNBW+rmgkVeDJNSMteG/EMdRyDL1gDI8QWLGx
2KXKrS4Qx9pgjv3ySf1J1QJsd+YJsbdZ2gAr4Q2qNbGLVR0eJP1/qFCKip6u1Mpu4/WruEyDYbpB
utEhvzht/ZOdB4q4jcpzCHXJb4Kp7ZOu0Qr1/vDmiVZgmRCekGBYV+7m2pIAUqjShQY9WiDDVJu0
Hpfe6eEIHGH16fGEkCBhgypj4/HV3DS/y0cllSszJDaAKf5wjx+B6VvZYh9Z/6f5L7z2KNYAzaHD
V+tEFy1F+Dg+NExOy1CUXtxMp1KBSjm0seFtbZjSFLdcizmCFnWkEaB9Rdsf9orkslWbG/vEY1Eb
BEi0TC/NPHXWHOxoGhyVCJXtwdChmL4XKbgeQwICNHV9pyPoPLEuXZEe9wTVo7SLaiNmQFnp/22B
mWR4/eY1Ftw0l50Cn4DNJ9IU8dSuIUItk/AyyiWE/tV42Wejs0ONW82gEmkheP10UAKdmEH/BNvz
xPKKCYSacKCJHwZnN411eUGDwfPNtxW9IHhpBZq4QqgN8KgOnzNMtdhFQMItjvFWRYrFm6j33I6r
F4J7keZA1OxD+568KpWOSsikAj2fFEs2x0QMrRgg20wzrXNeNJHZHEZr1UVcDFNYXF0szH7srxQ2
wZah//YnNx6dz08nS5JQjVF4Yd3H1VJLZk2lYU7uJuqhgHhiihvCATcTwavIsuqIamWDFiQzGWFC
KV2FwV5ePKwbpKykN8Lly1LeYpiiRJiQQ1EpKl/3x/KnEg5O60GAIM3cTxvVvpB4t74WzRR1trje
m993Ze8irOfFFKI6Xym16KFTllBq6lBTDpuN80tAMyj3K6SFCkCC9RDP+jBuxKyUQnxtVAWYvoE5
oH4eRUlH1YgOYHsv/hjBRMI10AilYFh4ZlNT7gvBedUit1UZSJaaCXHY/CJgvMrhqW6XWr8FF77t
1CXyl09Qaei4lraMefjmQEozm6dLKp6A61aoQNY5M585z60p4l3Wwtpl5kN2N9G8Qos1SOiLrrL3
HBcwKVkhheQNIVFp8B6s/duN+fG1zUohU+ya5s2DsVXFgbhs3cgxzCcAP5XOh9LfIvTmqge0spH3
xuiusgHIi4yxXP6V46sHddwwOJ3dIw2F7MaRhTczqg6lH4X5MLBrhTn8lkAXW8vZKW6hA2FapoUW
nRzdZI20vafWNm1wm5n0QfIAPF6zPJhqLu8eOISRU7uB+esoNDeWRj4bO65/R2CtfQfGs5q9FJKj
EhfZMnpuGdIKzkxTs3fFx6s6pTNo5j6l1fB1sP+touV6CJvfvceetyJEFfnpZn5ig64eALdQjMMX
SEkt6P6PqW3wolOtoECKo7f742XHlVZSoHdN5XKDqHiT4QlOdOeGhW6eedrISaQUsmeiBqYNZZnq
IBsYSYAKyI55vf3d3XhdJqAmmuBL/OjmHTgXKUSyn8rwQACs4hp8yRXwuroS1tg0fQ6lRf1CNOou
nPeT4Nc1RQglDRTrnTb9aCu94iu6VtYPCLzaTrkaOtTDwBTNE9omAFZ017ubhejcGQ+P9qI7p42L
5QIEc2vEs4jQn2ynhPQPPMG4ELtnYUKBBNUZ2cZWgZvoSJn14b/IySzmL652pUy4RNYkXnI06pME
Ru6Rp16BLZTeBYjkFUzn112ajVbVBjdskvjfUQ8X+7Bh+J9C3QQHU9U/R1NM9cIVzUbzbrW+DA+R
izfbFWxyrOmcKbotbioqq4qAHxBH8pzkHgLIW8xWs5/8OYJUrwVRW+I2DdXUKY4L/A66//wEZmVh
TU0jOWte5TNzMfuHvPMbAsOPtJBEuHZJqHDnYpNBsb3SmQDlGnBKeSoXB5x61x5jcvbZB2X/jCzN
Bp3juIJWU4oNA7o8doB5DPd3RRWilpT0Pw2LOVj8jA3AT0M2XMbxrTiKZKGolomdoSxXV3XrNBj4
MFiUaXD0+/tQ1sSIbcxkW98Qyjble0DsFQQQ+5D5MKGo2qWyvZvdJm7DCKRj5cyh6cJHt5Z614PQ
tFSvyglTrYyX2HmfQTcVjnjxAHh4IuLenEifdvN6/0AgvCU5xYhmsHVTzdCz6oKvo+G+k4VvvUex
hsJlcu/+gIuZmqvtfIT2qyCH3hC8wiUP4vticVfehgOMtdb4aqOK1M0FKRMl/Fc30FsWyaYOtKHU
lGdOh2To4dKfkBzrqW1tNe/WOiyBzui9vhaU/v6qEFOb31a4ZpvHAM/Nh9mdd5wMQ6CeQ4uD09+p
pHGfiaLRxM/qApoS0pK6D5bYCPXGdphMOFQsdduf2H8JbWyGUkKzp/Xjqfy6hqpUwO4qbNc7STX/
bM5KhGR4mVb9Mh8Wf1MKyfZJlZFGWzGpGzpfLnMT+FN2bPNGGCw3nXWx3lIrU4BQ5Cb6/aRVPSRn
f/1mlBF9YasIsHmUTizbA7h07Nv7z1ddS7X4ipmcNeVkvUEuMOPmGmNqSldGQH6gVpCRedEFUz2T
tzFGznc80pqCvaicxsk2DOqmRNfslwJhxK5+7dsKh65c/i1fTJta78+guwFr7rf6hN6dvDZdvU2q
8XOMyQTGYqh+OqXbSCGFHD7lwmT3TgZaOoPQENkw6kqEE8Fpx4uC5Pk+vRQoJubLj8I2oXqs3RMZ
3k61NQ7uvgavgk5eWQEH+2DumC2iPhv+fwm22m6v1iS6V7Fg31tIR1zMbHI+MFLWzZ6BmhUxXX+M
5tYbsm9Qwo4Vp8T27PbaFriau6fC1BA4IY9vDSC/0/wtF/eG9pJM2oy991yR2T0OvrINRX5PQAYH
ofejZx7E4dzcXDXhP9QD/SdVkkovfdQ7xYDPD1W12bUEKlFVytQC/2ck2zw5M40psqaJCgj2W8Ui
yNi1toF5cMqIWzQfCjeHFiy8HeHP6t4Vn9PWa07iP+l5+WlxbYCsEIZ3vsTWa5cENu8h30NzP7tt
L5Tv9Csektr0/0rBiiSF8UFqYL6xbha6rKcpDvsW0/HovygjgE2bnIqSf96Z8h1DTOQ2xF61xqoW
881XjVlHd1znzjIbO1jwIxx51Ifq3gY/XT9dWHNAtQ1GS/zuzyI3ZStyF/veTEWBJWSQqqZVB8Z2
gMqDjw06xmcCTAzxAJHuITveZbfog18fCIncBRz2OZUwL2OlNMDOSxIUN4AS7hRmeizjmW81Izdr
IHFvEbT+Nbd+7iOYvjT6nz/FvD1a7eZ4lX13ZXnkFAtqCwIjNp4L5qqrL2kFnWNMAwe7bklyeLfG
TwfjeKjwNbvpS0bCl7YV7yn/+BnAn/pUHiEI1bkdraR7Z+WCXn0lMPaefYkPK54uLNCOOh1S37JT
XEEh5j+7IiONpmL1iYegx+Q15PbWhzYh/q+2zMXGeGTOwnt5Uz9VXIYMfnFsF2upuUA7SjchTqXn
V11ChiJfyZoJrsibfEetQQHq1lJdZgVWk3+MQR//TZHSjOH59g2/VW1U0ijA+nDNmFbOgaUFBdVQ
/R6SYByt/Qn4d6tg4T06DdeuDtq2ZH/h0frzZhKngSZBubSCEZzW3PP0sXldpSn7kP2VWGxFwE2j
g1C08apKv5q/R7geLu6cBq2IeKyj6aD+PbCpRlmGmoksXYk38bf8xlI9xCA7UKyDQNDsFE2roww4
SoTUCYTQrD35EV/RHQkOmlsUqyVWgMRhfXvGW3i/2xwJuFAojB/4e8R4SSpw9mi0lRUrf+VmUwpI
EYTxe4ysSp1N8dyXtcTTZnpw2vobP7dJ/5WkCJkWM+wqrMJJoV+uSFahWqHT9AjKagwOrgro+fLm
nFTC2iUGrcVV+UPgCBHRWYhG7zH1KhqCR0X1VSWWbPJghdFxVUMzXPJvBvRV9gDWj5EwntSLfBhM
gUFszKdP8HOjNmsXRaOuqRdz0DxosUVL9UDT5QXTTy5YWtfR69Rv08LIHVKteLA8PBoOBwCfpEB/
xp0k6f1kVWGSDVaRis3RY8ESnYO4hOmSYXqs70lrsJWmuvmKzwa9kk8eH+D9hpQ5GF80PUgRJm9A
MLRV7/m2yDVw1GRpuxpZ73g1nLMsGBijEATPsgiNoN2kNPKgJHgzAr0UuIIvgH6fTLyJ/cVqKQLe
rekdl/s4kZF7SpYSBfzEVP6jaJAfu5cRILM5cdGfdLKfcGaXYb054prrjITRjnHQY3c0MIVZqf03
mGsqL7+nHf498hoN6pYwoFSn2GF6y3WjDgOtrQNNRv43gNqkPTVU1RdP9bbYWgm2ZOkb2hzQxJHB
a4Vo7kcjJeVrMvj9msFxEPZWLUgH14e1l1J2EAszE3e8SjsphVeP9dpsMtYIYrk7ogwgn+96Wsm6
+cdUXGt5SK9VsyqCew9rhfm9X1zJQlHmzn7uEr9aYzjcbDD78hV7tA/kugpHz8mcOqNaJMtxQS4p
rJzYSguef+nAtunpJg0JiNYrHSzEJKzccJHY7YDmtIqNvbsVGd0tslgnVl1wunthhThjCH3CIO8R
gQL3o6vBKROWVrlv+urcOnlGr/5ZHgDLKqNIq7hGgbE+wmtqGp44Uebr4ijTs1HWnmGy22G20glZ
j7N5/qLwMWJGA1dLyJd+rnF1bKgJJhHp+jv7Z0la5/Gn3i5ITNQ/P4YsFzgJiwLC1lJeRkDjgTSy
a7zGQ6a+zfEbJFUBhqcwILYprXvnO/jmRosNXKCUdz63Y+83Iw/OaMWOLxGDVUFWju0A3s1eEUsl
pzZBc9i7SnVg8qUEMPtJbwHIaDBrSFffrNbtRk3CsuM83q5LiN54opYn3MAS+idNv/IXJJEW9DVQ
fhtjhgmmZoGuPoNiTq4u4c63pPHMQ/vpR6n5xFTMt4SQ5IXmM/fgHniXUJhbbFqtZV8BuHnRsGVk
JN3sphsX+z0r4/qzYoGQbvXYLTrlIs98tuNr20eVE9+QtBSCMiEoWeecWvWNkVLnjDK14KX26NsG
g6qSw7JCY0nVl7kPFE0uphKCTG3Mj9T5vPFZvAssa2tYiIk+cRveGZnHflCQ7Lo9x5zF+ub6OBxL
M8fcKrWa6k28v9Jgl/wqVONKnPzB0OBWrI0gZkyLLz++gfa10OBqL1941jUFiVNRiYn5tK1KVXml
WblVz39mwJ5l2UvV1IZs8BsjmKXt616N1X0rgcwuS99pvqqIRRRKZOyMW2+Rt8piCN77wr5+yP0k
wOb03DGuPkfgkw1cKYkIFQSz9rZxRErjuom2Iz0zeMHCy/Ta6NEeUeEyEaIIg9+ZwiPWzeKAGw4x
uep+vdGE3HwXaIl6umoCExW6vG8o8I1sXm2flOctttT9ehdZiyEHJQjnuTVqAUwmzG1+mjMMUuq7
aH5h/v6RJyMCEqIDFNZwcClCZr0CrJX46JealwAzHNIPIDmts04tjSZyGFiXW7ttTSCeR4Qbp+Uk
hYS1fGJ1yayGRsFx6X1kwt372ZWVWaauncrwBE1lyKKeVQKkIO+6LbDTKKcA/V9pZM7CLVUX3MvV
//1nmOEPRJamQzMY4JjbGmHVYxO5bF7mHapN/YndBN0s9b+/2E7vRAH4JVpGTPdVN3C+CQxE9fjt
OStaoaT1/N4r42Vmhcl1jMc9XV46McRig+CgPSeLw0mCe1d2i4Ps3zk4VHNaBJtR7mDGtsGI9kvN
PzNVwVp/e/jQDwrPPiZLbJILuD9CQ+HBHMxCqyOzi+BR9hGbK8yqYr2CeSi7PgmfikT7osnLyrRD
sLBj3F+2fGp6/AnNzeyRupL0IkKXiqbWnRl+4Y+VB4I7b5slSZb5PwPphNf+5W5XLnFC0cFtcn1Z
k5W3kQ044Lz0q2zdoxplJY6AFoYHMaTMzOYD7soWzuQh6lZbOYfi3Uw+uPiUo7YTKSkywF9nD5Vr
QnOlhmn8YQ72pJPLeLOYrA5sCmz424Xv3+kAAsviy7+OkJtMj8SvmKcCOfrocWHNBqeZ2tc0dN2f
U13/NqfvEOOHvxLlPJnGQJjwrVjC0Kcf51EjfMrtoge6oDdQcujEhNxRH74kZ4S/l75fEoc5T+Tk
U1aKq4ONLO97/mNn9Nz5RdgvulGxTNiAGdFjyXn23rlxZZyvIgqnffvOBFc5OisQ1ZkyioE0UXGQ
5YR2kjmkzzK2VF7val4t/QtbZ0JugFOO4LPyxlpQkIVuEG3L+U5b/ezUEysNF3z7GZBBqbtn26+/
U123IpQpdaOPpMlRSFWTFlIG9XztwPPCQ9QrJT+Tpsa+VBuIiv5XFSyDm9bkHcuA519YcWITALhE
izfwGaeuUFJL1tPhDjanzhETEcYSxpsN3gjPLTRivUqi/41K9GbOoBQSAIEFbUmU0SpEJGVg/CUh
z4mRMW95p4PSjB2ZGt92QOcBFjMQ26HTIBYmN7P8Jkf/d9WltOZ9ql/wcmwr+oB+Pth3ihDmAwjd
Ty8re4U3rGA3m/X0RLg3QGZaMgxdTwuCB0fyTBAR3w4UNDPk7HSAjBGGKSmVDcWi8MukcBzdH3QG
FOCCLCG6ilSPbIFlVS11EDWAsrfoPb5jYzfCc47Ibas9j8/zcfF+VIkqVVUjLQbClMsyr0BjP1TI
3kEzNiU9OXqHo7QFyrWmlXJAa80xI1iumVg22vlLsA40UG3LapnoLVHIAJmnqe2QdjXS0UvtvdP1
aLGPKr49+XLpQxHZXSbwjG4LVwALMhMfLaNdV6manAuBBJB8SHMmX7nvVAd2y3xyrKVS5C7xKYt/
JG/llbgAEozsogGdSjjCYPoMqSt6hiIcW0btK6j9NGVhetQLHPTUzJNR/ahjrjTz11iBaNdKSnpH
49h6wYnh/lfQmGy6F6Gk8IsPG0CjwfPpeeO05qqUZ+mMA5U1aBOJy9U6Y75f3TAsbgCk9ZljLZMD
cEFGPY3WQTFjSCSNlNTCGJjlEiQTt6V2N7F1ZbIL5G0i58Bij7n2eoRTVnq5sAUPBTpe85iRUujE
d8X2suigxYzVbvdEldAssFdjnKb/5LMH60D0WRlKYcv3J/gwyeLYgtIbLh5/c1hzx2QbLDJT+mee
ZKPzMBSaz5GiN6iCismWLqtq8IHWdDYd9dsaCBup2ECuWuE+u6qqvp10Uo09noqTDGT2HsUB7koz
SCkzesLxHnl6WMJA+b1YzlMKRZAhNVwBzDAJZbuKPbFNWCnwxp3aYvbm0SJt55DlGz8SFcZjFDUm
VRPI8rmdacKW3n6bi/Y2j5Pvn+HhsCJTZk1EVd+JUqHyv3ZIZsA1ZseNdpC9lqXhBqnfM21JcwJa
fV1gnJ04cCHXeTTSCVv7ArwhA5Q+uGx61WZr+j9h7/v2FsbfVD2jB3a1dBZBb7N4gxCEKcJWs6bK
QQV/cigQG4bXrihEaQPq1vlQPGPuFODuTK8H4FgesfQMQ0DTWnuPU+A6+dLDQUwp+UDvlMlQ9H+e
Pt0u5Dvvp00I52TaWfhViCkAqkI9jM8pl5clzI2lwiLZrgOCNPMb2y+nZbKg0xuN+KO75Hq70/lV
X6X5GJxWE/C5gEuP8qX3FKV/uCzzMdqgRpKz46p0xoc0AnAVFOeVA2WFWh7NQdIY9nDfw9iiVy6o
Z+Br8HOwD64xMCzjzef8+mvhMrJoV+t1LZ3/gYOwDrt0APECbFqk+MDwXu/XIsOLqfa9AQiAWvjz
cUWSUcsSaZFPiofy1phJYYx+5ayzYns+OfE3SO8dO5CwXfmDRw401Q49SNg3ao59nIEIEjyTLhfZ
+H1jJQK07uC5bm+vHIVFqotRNG2vVqlmbdfk6raIZWpikcaFGK29LeDfxpBicunem62WStZCnV5R
G7fTIucOPviL4Q2DtHYL4tK056FuN5sPvkinBh1f4g2+L1gDe6kdVhS2aLZUNbKPGs2uNFsWlXan
9EbxFJKQnx5Ry+3q6RwYw2iBi+anIe/ZEoqBJ+oCiC4+W2leLfAw34ksbyKLmXv+NfIdZOtUhrAR
fB6pyzvbQaUQ+3Sa7WZm+f46V38TP2eweecY1MjKIrBUHnQFHGNUkC4p/DmLv9E9Up2jfdy7hzVc
S+kHPMlyDsSPS5MK0jkk2vmUyfUGjGwzVkvQjaOcyhlvSCnqo3HmHb6zpo6iVVpVGnsyMsuPygbH
hL55okdcgrishb2bh84xiKFCxFEyUB2DPyv5BEI891hoC27fuGiCZFnHJgXW3eBqq452s6FBRLxJ
RyOaTClkOJIBvF9JOwtCKgUa0imLn0HIwnnMG6YqKa8n+QJP1f7u2OI+sducOqE1NiMzdUnE6EuW
lUNYIJ3Xl9DeQinAH+qF6wc5J9M0ZU3DBuG3Nlp/ASgpjVDuFc4NyC2UfmrgqszZLHACgjVLaxkf
HmosGUoSHI3BqehMj5d2tpmBT/vWb/MUBS3DAjPIk+uu4CncvRxTZBzg+z/7Zt41bhST0ybvoT8H
ToW7k19XBbers4X6n8FPGtMU3reA131370neVx8wnZ93PubCGiD0X9MGAQFQGzO0xipTq+vb3WYb
Fk3S0D5VG7+oURsh6Loda+mPiZrxcG9XMpGAN52Jdxh4iw4fZU3pt9xHpjSmidSi06rySXMaVDY5
vjTL0nz6c1ZN9NLQnSFvjmFrGgAgmjCOX9V4VXn94RoSGH82aAFAHpZS7GL5DN7ybaNIkM8hdTfY
/sdXMp4Zv3nWdtHNLJ5BCixpuH0hgn/i101pHCN5L71VbTXUB3vKhRMTrFVTr4T8yuwwtDCgcCDj
YDajWWtDSI3BYcIQUWK+28ucJ4h4XsMyG8xi/9Eup+g0IGTH1ML7dKwFrAszS2KgI1oJp82blJHx
ljA2jtTwKbQViO6mrnMJjLofL2GY4S8zmSLAaaoCqjn+2HPe5YpMyfaegmUdB0Z5mgqK+dkNviBN
TyNtOeuLsX+a0JmvbXhwQZ4T2TIr7RKEJRu7NlgKTWuT15A6SzzNMWaM0e2mcdDce7Nj0lGlvsfA
grzRtC7uS0NS/6xu9L/QDeg0ebn1Gwkvl2qSAt7fbKfgG3Zsqp0+6odIFYcqY0+OOaKY16ABnjdN
arIpdT/lPoqyOzUNmxEkAjFNCyVtcqPzdTJQ5RSLhUAilHRZP21JZubdBnvfWbSSCURyir7MgBzi
acu/8UP2r2PSu4Y8Ga0Sq+8FTG2YDj9vPbsmT+vqNCAEDnabDlV6EGGe1g1Ysa0zGseopQf9tEb/
yT5EYIVdghUvH1d6PhLExtzNjj4aSBb0I0O7Dxf/EXkpqSoWY7ncxtxW8UKKuVMpfoBp4LY59VFK
LqUuQ6oxpQ1zzb+PBa2RdYcObjnKSOpIg/JOOMyFQO0QFm1YIAXw/NoVf5VaPDfZA9ohVhbjiFCZ
+G0LHGz3MrwMvhJthg60TichXUjhNZOi5cjH+WnN9pBvbhyN+EJe6cGrg1xZiilcxTDuAO9FQOiD
qqj108Bhe7A/wJSQJJr/TZUElKJyhqkcK2GUtAuDtGGGjEoNOghpLJ+lRZ1xkSDAvswlfNk8fWc7
VKCHfGF+GbvpUT8bgsbqiNz6nSy8E2a5fhR1o2DkXRdHT0HiwdKcM30Tw84EzckIZH1XZnXb6g3J
jhVLNzHy+/xqrP7ojyLL/YDyRb9XayTacCXNgJcFZd2lYMdVNY/aAma3x0YsseFx7bgI9bJmXrHq
sFTOzYc7zFEXhoCRmDHazZu4Z5B0oE2vpeDTv5dBcVgwDEqHpLn9D4EF4KPdoPOgPo8n2ktFf4qC
WKQa+F//r1zWssOtfvDgtzQFFKgKFaoK45iB6hOp3TJS9XF6ZEm6kGXKki4atqDanvxPWQM0MnbW
iukWrnY7EQFmxoFhRzRN9LjHUtAC46zaHcUS18Qz//tzYRzi7fwvu0hwdSVcZtm8On402J6FnC2B
Z63ZCmy1QXVjBuPTs34FESp8dT1q6DOjg6Rw0qhA0mKI9L+CXcJ4vHXcAdQ0j+WT7MmUAJkLx6Nz
C2r5txoyonb4s6lM8hyASMZ/feadgzHg0wIUJSZk5Su0a9PRP8pPOEQjJbse767pMjky8XUw7Rju
iXNVmLqmaVlURYML5UaitDi1vxMPXpkQPcqiJeTGovtYAaHjEqCh3uLuJ47rLkmx7QtcdQFN/mJZ
HB4WMU8IxiQ1lypPjknz1UAe8gJusLX23gwDaTCZpmhlfCdMVijp5D2WmbNnb7+xxcIIh3BMrk+E
HXxbxHuNEKQYtzSDKMW+wwUW9+D33AfVwZMv9Lw4diDfNSmTWa/loclrDzvdxoatCbL5qiqQpddK
vmaeaQbeA/8hcm8mBDSawpU8Fos5fI6f2PsX/q7rBZxrvhVXCSoZHN3P6qRutLt5wgqjo7Gs/Rxs
JC9XNEP4S1ozCFPF9IGm1SO7nuRyTS7fEdEIbQXVA5F4ib+J2DWNHqy6XeGGxpAUT//XU/iyZPRv
TaZxbM6lLcwYvrZ+R5nfY/opEcbJVZqvcpSKtv3e9RrOS/EjlsX3evE1MP31Y6gdETiLekU41+zu
lLEKDyruASTh4LVqMYtz7QpM6UB1knEn5KiXvJV0ezsuNHAZEaC6vo9n2pQP3A50QsviiuayoqN/
8tD55Q75cSZaTzBDGPsOSx68w/spTtPixQPMUT8+PE1lTT8FYbFXYSSaPrTbl+rgLyWu2Q2D8wLW
WAKRVI3pvtYnbTLRzHrRvgkDWH6SGsz/Zp6rSARIcTPqc6IT0fsgvIP3s95kx4CqWtS+YD0j1Y9O
WeP9CArH/0POfZNMVvf2NKm0sN+uNMVQdEkSmhq9MDthfuJ4ATZTc4A329e5GbvcvXMi4B7gBuOh
4eY7dGvAay+6uNiozrGPZUxHv402ScQX698R7FzY18WQDKX3hhs5eLuxQeKX3oBb3mgt00XJyxaK
rz/px56sWsq7RBYvUI3IU3Uv9yKnXShEKHuFIs/1HG8bCE2ev6It7DLS/xoxIsLva2YzLHGndoRL
Cvk1B/ODbFI6FoI0O2WaBB4N25w2b7/1BIriLM1bs6q//sNfKMaCqOLI/gtmWGBpCwqvKPk2Czhy
dy8TA7eJk6qyWSiPwXEMK7MhXODvXrPpDBMwFFMui5a7/YRTZVY23tzpDpgS8hlF3vqNeCDQirl/
TyM8ayMuAK2MMvRKEG4EWr4YtSgopq0pheQQx8PpE1iijsW7bvZ/0AhJt5avylTcL3RvPVmm9pwy
573dweVAanayv1K2TqHoiiKPAlGKMMt8TgSb0dwuss27xrO7/oT3x95bOWSV9HdeLO4QmkwriaBp
lbPs2pE9SmpPQgxB6it106Jch0mcEG6W3vXmic6XTiQd8GXtsWIXayTVgcpOHzZuVmwz0jvbhzk/
c2GcVoyRc8PtsSLcv8OxYdUKoEw9yqrT7fMHq7QF2OO1WNJ20Q8TT172h/h+ZCfQKJFAfRSbpI3E
FC2oNSth8wY4s6OB/mwu/Tiv9A2fruP/iMdfEyRzF6/AdH/1CkTAbuLhkRj1q+cdL5ymb+1JfI+N
1LDRWq581beM616IwWmqK39ZwouQZcWFKb2HRvk8RI7hsc5iNrCqpHt20FxC35/qs2E0zX1PXgca
AJfaIbcwsZfYEEVNaId7NSDhj8Tk1BPUo5NPqM/wzsotqgMApi6UwP9EiM0kQS1510YT8HzHRoSV
fELQALlmcOafHsScHk/C5aZQZ/OauVmU83CoNJGsX2AqEky7I9dv+5AekbnP0DEns/uKLkUkNOi2
rQOayWQlJhsr1ghmJUqgDy3qnYabcBTD/0GFVuP+EkZTKs6NMAHpIez+UG5NCI2nW/YcArDIsyYA
dgZF9dxpInEccWPL6UQohICBo3QIaMuxLxm2A4OkkmbzD7twxcGJqXSmpp7jz1wP7r+nOk6g2AIw
3IJNuoT907zflPn4zs80x4pQEN9gz7cirjwPqW348kJQ6PRFmBjcPh9mtx4Rj7MJq8sBwQUOCa+1
BPnBhbDSNjwUcup//oxnv01BW2qet3UP6AHAjFjiL9zBeF5QOrjYKuvcAWcXfwh5IX3BIMt/sbEf
HA4eu2uzkJJKC8ZraoySMdGwz9CR0vTRXeHeMWsnfpdrwMw9JmxWjxYN7vogVK21nMmnJrO9zKJw
YgN8QbpsRgYF59DcwUGE+jusdHmepZWZsj2cBPVO6Uoy52TrCsvl/18lvvqBCbi4SrZzom9qVqF6
JiH1v5C2wiIrxS/hCbmdfb6YG3NiU3gKxGk7IV+uMbrC34vwpLZqqEvQfcQx81WR5qv6+kvSRNCQ
LYbHglOZeyeCI04WJWfguOUyziicl0Iq16cTV9B9zH/yuueGGosY+MLDkz80mQ2q2knGW162X/Re
fQivO28N2ul6kN/g6pKSoXhnOYilu6O3bm2+oclOri6S8o+0aVELi9wgrwabGCrLll2a8f/AGCvv
t0zBqnuVUbM96jeiMjHxDUnBimXSZsKondQB4aTyILOWtQ+/aEXJOOSOVmqzZYcEphEp+EYWVAL6
ob5R6N63BffxCnObDVpO8xTjnc2jtUKDEhcnZbjwI+SVlfKVFPxAFRuVRDal2JN+JuPVpATAFbHw
73t8daeN6ozRWKfep0qAAkaxr65O87xxUdhxe9GeMojLfp+sk6825SUWMZqabgMHZ/m1QUxjzB9s
eOINuGSYY1/bYIbRnHGLcH/UwHiPfxH7L/szPC+XcRXdaTI0VmPKPB1ucZo88GjiXPAXzEt61Cpv
koC7VhE9B5nH8ln2r4TKtq/hAbHeb9u0PmQOXZtvBdW17eTlA0aGShPVr0t7TA1ArM2gk8pAuwCH
FYuPM8Nv+IAodUblVbgJUXTRovLFKm11sk3l4idDzWr8mODXwzkot36BPKfk7psCwqCUXh087ulK
jzjl1V0Cmm9zD1xG9KhY+3RVjDToWIKPOVPYFzqrQhiVJjdjPRKpTPK9RympG1d/Zis+h7O7euYi
yIoxdwuMLV4i6mENbVeR6+ChvLZoVf6VWt/4LCL6icVPlxn4N7BeTk6dslAd6lWUfIxnxk78tABe
4Sv4DOu0/4BnFvoGKbw5bJyx5tqxRJ8sICnct2lF9R876K3H4qErkTSjhXbXxLAMtoQhsM562Ufv
6KpH27FV+LKjPdHngGHcrVxaGb2S/KJ9YUdtvPM+Axrcif0Tr9h9aE+4fEHh+RvGd9ggg4rHXt+l
ADLNOoPWaeI0NlOxfqYpariNXK50IpXsHUQRZ6RTLe+Mvzkv2kXPeL0DcF7AVytgkMGTEwtrMr/m
A/rpQKSCkYy7GHtTXMgwtJuYQ+DpHbyL23EZkz9Q8n4U8seYA1zq4Q7C+5dxLrLQhZ0U9u/vUAL6
lkxSB8T5Pop8sP9FEfSHM4Ny9rfyGkjvyXJDhupqNtEhvjAAvWqVO1h4sVGtGdw7wFM+UnNPHTDf
iCL/WRFLEMvWwoHvtBLY4YpRTgoldp7pfWopSDrpYoP2zrqUtm77FzeXYmRx5gYa1lRjGp4pWkHX
LYiGvuENB3BZctmMHcbz0IPGRbxgfpI6nV8wESgUhDNEyb0uZuN+DlVJkCK7+SSQMTckfJi1Fwwp
OsIh6oJrb9sb2cDoA/lJscnJs4+a80DBpx/NsVdtewLTwZswXyLpC4rpvNLGgVGLzagadUU90co1
MHmg1gIr0lP1N363/5FbE+vyDYjZTZdaY6LxkNeIPkldb5ifDRMZEg+eLlAN/UJzs72cmk7DsJgO
GCeSGdjE30FoCZZ0/jD5to3g3Zq+t1c87MWctBZAWH6RvXfdQ0xe8eEwTYXRfqkTDIug4Bsn7cVl
728uRY/qfBxXedqvkYoGEZNQq7/YQWyZ67J890T1SIa5S1ERzMJhMdIcMOvu+nLVdc8TwJilmrEY
7uzdaS6sCz3z2v3CKti/OTJ2+HL+j6pLUrQyr6skgWv8V6Monnh6PacHq22IRn9o4bsiM8QQmjUc
w62xJTIFvrRszrGxeMvagk4eO914C+Uw+vd01iU4RkR87daxfsvqhtUASbffJQtddJ9tk09qdmaT
iE9hr53hNMIQrz2Bln/NIaTZaMVy/7HxqfaL0Ih9Ls7h9tCikfP2GFJJgXoxIixwGz8khqaNL/AB
MztXu6v5LeuEQ4C5xkNj0maYQJPJFm+MCgmHohWWCcxzBWv4X+8neYGocBSqc7Vkw+V/82LitIrh
tp13MzGzBPTaRNBxy8HxSRgvFf36ddd5WKChiX/aVrE4RLCyId5IPBroTbJz8UYeH2Nm1nS1cjX2
v1aPmdZK1apPwvhvNByexjI0EYguaJBH8AxR5aLExYKfT7xV/ll/+pZDRMV5cPZAop0/4Dlyeflt
RvxvBHvZs9CWHnhr9gQPi3VlGPFiMzgopb43M/XO8DqdDpm+iHI8oN9gjBVOL7RP0rqXkCUptwkD
r7IWL3jyhHPbV3doZ0Qbx5L2+OlxUra73Pu3cO0KlFocm2D7zV90cgLfCE62BeSwquehTQXlixVC
8Lds/fAmbX0fXrMGWQtICLVYhBpcBS02V7kY60SQM9KcahPkAaY29vyKyTFJzTYraPIGyRfjT3dr
FEHBLjZDpPpN3mTaPTFmlBSxZ0yHTpZ8Wwo0FGM8myFsX1j73m1pkfbaagp4/eN8OJ+bhM/gKZ5T
sTM4vmuBeAHsliSSSQuavsr2wGUSrdYJYAkGOl01hD/A0UfTb9fHC8VyurDKErLjpMrGAOrSifUu
8JJHtm2XltQdbXf7hUdv2gGtoi5Z8Ehnr6mhFB3j3V4UpPCCCbMnGPRY11is5MdksFMcgwy2FOtN
2gJpOj4TqnxstbBd7egVGQ0KG97Wy1JS8nmbw8dRpG+1cUokg+rkQ+fTyOykTxLUjGDTTS+9cnjU
am8bd9OYtVWpvBxGOOL/MJqvh7kuJLmHvEPCbNc9wV2pzkGZEofVepcHcsll14G056fLryYUVt7p
MVG3Ai7y0vjzlHqSglKB7C1dQJAsqVLB87V2e4mOfkT2K12zUxDlZ3DooPgdv+IOknJ/teXgKJNj
cgLemqZUdAHDKeFS6SMNFhE1kM0v57UDFu1I7lI4au+yE+mD3pVWblnIWmCAh7uZp2jQJsrTSPv/
rRbdcfrMUJyDtWxnd6Oovl1skP5DPJaEWH2XeCrRGN0PZy0zvrbyjHIczTuAM3D5W47Katx0nRPg
Y7JC0rjVBtZzM20txGbLpxvuyc41tU1lGX4NHVzdkq2esIL7qVmy6jV26MpO29uy1GENIl0gXmow
z0IjtDjth2HVjKQ/v2E5sXMtxPquInYQy//4WPzDBortmKOLIhrzeXRXSMSWHnDx9H6tmucC6hZu
HJUryPw+v1p0L8NhUyJOG+e1Qw3oou1hHZLuoLMHNsqVrvlMnjAcYpsBXkJ7TnCT0vKKeU8w2nTV
/8qv7VhQB4bsAOsSyuzRYMPu4b+0BPs1vJuwGe9dNYoOGB9HVgof6VwIY9IMJOmG0qJR26sRaczW
FRwPnVx0zDkypktnJHPHDatkoQ7dbScW5i0YmFg9J/2M7DroaU5XC1gPEIW4ZcPvD/pE78+CLz5I
2Cxq0SVXGxa7tkhWWXmLSfa5rctc0CJyEEvJ8HynyjSRvf7ZCd/0dy6qDmK75q0B/9FTLB4TdVzh
Cs0mLHVEC+GrsFBSip4fv2EwC1BF8pCCTZeCGhMyZEwByARuY3YymW+imEcUpn01O2pql9Lb6Ftd
9MK1XwvmfYy5GAzu/2EtIZqx663mcmRZHjo5WG1ARy62PaM+MoBI9hX33GIPSYGGujQwizcK2Ghc
6PmKcx3yvjwER8jOrJn743CCr8IKqR1exXZ9+gIpgnFEdNbkDyTYayZSBH13i1IepvEUH9qP8Uw9
qWI/yJjCNsktA/LehpPKawR8nfuDOwxiU1vmmEuDnwt3qLYIGM5dvtN0qv8mrdZbMuicWzk12Gs+
A+vbkOxbLUfynrr+SKcKxlKJRwyS252KPwvC+gf5FTYholi7LbdyvQoM15DafnMRjI8Ilnvma9gL
aotYJBlXMwgqvryWLW+tW1UdRlBepcpdzf9iKzHzYldb1P8X26d0gZSWKWx7zTR/R5csITfPQeYM
MzktkjbB7FedAe8B7ZkF/I9cs/gO5EM5RVJ/oJqi982gyc8GXs0R14N53dlZnVL7CNdTk3cPjC8L
XPX4AEzdlf7ujNtaQ5sGUxb+wayHm209bjm3v1JKtu0arBgcw2dD2K7s3BRbWfiyAYpy0MgM6xTd
pxOuqWHA1CnAfe2pCmDIYiGXIYYCimjlzt1oGNmNi8LVbcWAc0BRrYfjb4yLL9darc1RdFcWhH8P
QAzBcjX5ya/fkfu5fmtZzbMxvWxe5Bn9Ad1BwjRPREOkCwAoBrfi91iwHieKCA+dkO+1E79DPX+B
gsXqT0+3on+QNunE8Ma7M0ncBJLM3oy9cRgJvupgJGc9tusubojKJXtwU+IRWAQiCUpx96x+SF4I
Q/3Tue8eVw7mcl6GNklpY2L0HlVfN6uKTaHC8zf4I1WOCyUMAtTQd1vKuxDfhjFnWXKAzcCwCOg7
M+sAKMs3WERarpVKzQB1s+HI5UgIRUA6XupuBe/IhwzJpz1kSY5KhOrZdEaJKjoQ9ot+sIlkFfbI
Q6HWPhrruWIlXuxwYBNWT08sTWSFDLntUc2+554v8FrDlVYeYZMM3wqxUBosUJlvnqK79ddjjrF5
J4vL/hBOO4NWZWnBow2/TSn/0HBjsTUgK8pvW9pBe5OvxMCrvmSCkKIP1eOl6chJ5gKYIvQNjAZo
1I4pxkhvvsLoYZswZTiNmlT4/8rkbcc82VIJ+VCLpf0q1nhwEzf8/huaYybCcRAinVPxV5xSIYiF
68i75ictryHIot2hzNQ7R+MBSNtkkxQLogv/drQVPIQ0m7MjnLM0YCcPUQ/UUsGPw39DaPN54Ir4
EIouPwoV1s+qWaeivpbpbX34EYqPiS3PKp0TcWav8E/3nbZRtkuiu4BEs8up5Tb1zhypbYH4ivTX
BznKi1aid6EzR/cQQjB+/oT0cbsfzx5yH4XzGodUkPntuptSPJKW8fVMLr4/mT9xdRfMq5RALBn9
z/Rqgi2CKiSwA0aBDXOtYAoxroZgff9/ILgUaPgk/RijN8VnGNDzGRAJAZhTZOfcq6wZOEke0GgI
DMk8rD/n89XASPSIvEfMuUWEwoGqBdYL39D0TeRyQVriRZzRM1vJRdFzWcl20dGj/FGzeiKTHHhV
eV14ETLlSD/vuGytS5B4f//WfrA7qJLobHZd6mBk3yZ3SMPcHYAPMGJQgtIGNFcVy0RgLkLPwoVX
DZF0RspT6hSgKG/adVe+Ow5hKkUW9R7UUq+jPArlUBTv1Gqnw36edQOEfZcPNDAlCGAn6c6H0JXT
1/cleccnqqeqkjgKMj+8rZ1zYdtZkQUUHTwBbSRuSKlnms1tiAFgBp88F+KpIBGa36IOxJXx1B50
9sDw5VeCHDRv5lxLk9/BY57DljJGVecUJjPvfB9HVCM1WLikK8GyfnYPf6i8PPspcrOgE1wHSNPi
J7d8ougz6YuiysOwvgobnQQoAWqM8bJ/1ZP96K3qWMZlLCvk10Ue4TQz0Ltg98pkluX+1rIgFio2
+zYRtBzlFbULHENbDQ9LyfZsjJ1u1J5iZ+Y/SKB9gS5hOsFdX4LN+pbM5P2XFMyWuGO1d2fCdqPa
dAZVFOpj17agc8b6HmvJ8blR/Q4TxmgQIA0GX+fdLIXA3oW6JQdRZg4Mw2BrkrUKYAEF2eOvRei2
TpOrzemSfNko5TDVd5EGw/itcIbJNod1ZYGRoYJiwCGX/rCt8TG17MZFlRkaM5W6xX5v5krX49iU
ANisB8vU0h+6X9L6+VIzYK/W5DPn7/Haae3CyCIWgHlGVnmQ7Yk7OpsU4Tl3RsJKhnq334qS7S9g
jwNlxtWlxy4Fz5ymHa0zI9Sx1n1nNJZX+AGcOPEoL6722kEDGswNttEycRKzAhPdu9BLWoGXXqVP
Y2jbyDlst/LChokv7nVWuP0jtQGLWVmNGEX5qcMSTaPB/x7NK5Sas82WycpEg8zeJHSliJPJ4TEe
RB96wKYq1C49MehIV+Jb4PHFR9UbD7V9EwHb4KBVY6qHW/ZtE5iN5BCWas3HIKIH/BfygQcr0sQU
v2WyNKbN8lv2Hm+VDxHadLQDNByi3ORAYpPSF1bXcQWvoNtoXjz4Rd5zVOY+sGr5yOGauFXMIN7t
FhXzSIv9VbAK7nyP5RxlbxmjyQoYmV7RRMjNJEqTIlxsZzR+K0gBIK7htCjYyUuoTG30QsbkJxVm
w29JIqN1ZaoR8jbyF51FuUlz6Obnsphe1lL5GG+PfS0luxJ8/BCSUrnUNaeF8SJWj00EGtez/wWc
iHwZN3k/JOQrLNUq0DAdcAkK8gXLzmSyLU7RvRGewtrWgFWzGOUObNAEdb+pyjMCBM6yUg8vUo97
BQqdQL1ZZ6T4iLd0EmRpG9tOo1ePowywUjGDBHbEwhhF6ZNlSgMsIDYgeFLucRocIiJvnLUUjjJ5
oszJ93BcggNhj0I/t6spFxw2m4qxdorYw8ZtlOXWfH9BW1MuyKQ+QtCqY+ByHgzIfQVUaQhkX66Q
yCNgEBDk9pD1OTS3QV4JeyS4mELKgR4ieGX9w84dsHBxTiVvLuay05PFOwSDfsTuaIJT40kXq9XV
/ZXbYCuubjVBCdZmZpFu2FJuYXUM1Ocondvf0qBwJPRecG9vwhClf8b94CCmEj4LOGUGSWiaE2QI
phdTHWU0PxEf73b/CKsO/P2TzGj614sVHsMN3Dy1+L9FAWlBuTXJWc7NuzwsUdh7BGPbkkKZwqlZ
IC923yL3ykcccE238Gk9Y1ykztcPelPbbVTwFN9GkZ4xuMPONujK+Usn5es0RhOKk+A0BI/ppd1f
aHTDoixyZZSkPVaZz7XcvdI1B7y2Gtj/5xy7UMQ0wZR8AZu/88FRN/JD0bL0vCXfvnI6L3MTTVmE
+Ye4FdNaR34yM6OF2IeEXwmr4Fw9j8SHQccGKCpr7gIhfyROwo294blrvu3wuXUaHklifiYLcpXB
0+UDOH8vr6YSr9JTjKjXTVSAMQP8+PEWu0P0SBTO4t4f2DD0PuxXf5l+OkUjIZ1Dw+drY7UI1iBh
bOspfZRPzY63p4HhtuI31oyK+vwoUHAbnJ2U3Ymr2XSfftKDOz05UyJl2RCP9fquJ24oOiDHojVX
xeoT4ypMUsR0PCGV6cE1RjESJZJCMgWIfWKGH7ESkH1vxMdubNECFJj1/aNI/A9EJXCOxhAWbYLM
fHQg0OjnTXE3OmPT8Zde2G1LRsVqbN9wEU1kUSwx0mmZExOr45ZsRdXbscqT4NtqZNFcXlFgT7DB
B3PL9o7lO9WUuxJ2NBHEBC+7Ix4tIgfBMAuBG8FNhsrN8Uzd8l2hWkkJR3Tt396t5fJpk+ToTNAp
PYEfAVCtzJ0P3npCcQYVymbxdDgYHZNrBLtDizaG41+GRw5EoWQELjKJlJ/aszLN1eYXqm59eooA
MOMn0RBzTVwtUdIj7C9d3bFthwjA5Zbo8Tj1ImHtF5k/YRRMI11eVmIFqGm3rps+VLjjtlyaivcY
r59nuobyusDSn31npRp6aVCq9vB9jmFKyeZjQmaZDvlUm9esFOGvH2NWdG8rQTEioxlb80Mjq/Ar
mu/VNej/dFDHvqjnKI17QpTDLLsVx1exC0h4ljTB1hC211OvQf19khcCXVvFXej9+AYecWHKihNn
MHqCFM6J5bFxGZd6PzsAQbsFwJVNEy3N8y4wNzNLVhbcmF+LP147y6hBKzRHCgXFllUSMwTVuYYM
yDl+h6xBcWBVDT7j73FA1k4JhVqKIECPsqbaf2fS8DtsXBcl+g7cLocjdEzcqCUdgC+ZUMt1CAas
MWchCgcIS1nr3W2MTkYlYTZewznjU3sO0zdQM/tpFUKjOdor7S3naBf8S7ipfvBWtFediSIt0mIz
TSEFd4t6SeMwja8Vi1KG9LuRH0WdtJ5KTWMb2gQC1+JYkWvgqnqyLNyCAc09h954f3DcaaU4Jvwc
ckDuq9SKvZRpoq1ifCT4o0ylVOVAxXMhmvBA3i4pobMPG9flyKzNBXfwZLbY0dE+6wI2KFOrrqow
FzKEGEEFxZFxcEAfqr8up7n0yb8Om3e0BVy5ba3b7Tj+jM+Ss02v0Adqzz4ZKJ0R81qif0t0OxWb
ccWGwdhkKYKzMBN5Fvz1LBsKoCWQZTubAiW6wrZ/HR4kGK6jPRIVRy7qjfKgabnhJaStZE3tkrre
wHnW/aPjjEDsxiBxjs0u2nlggWyn+qrx5ydhJRsUSxgdmSUWnblTriYYw+mySGMPli4UOhsmYvDZ
Pg4ORvzRVZ0GkpJoM8MqFWTVpD/s2W0Mid3m5mSiRV/Hjv7ZUeNIP6vqedyJKLff5VjXx0Hvcu/W
sY3aCuUQ5j9Wo75hz57ZNRqcXaPM8wYS5aFKsApF0T22dLk74Y4V2fj5lsXMTTIbo0TcptNad4lO
5zGZygp4joJ1uoLLA0XUhtqqUICc79b+4FnmmMCHhyQ3IljhnjQ1R/71czPY6LaExz4taYS08mpK
VZkYnGqXFgRwDow/3osaWFZH3BEzUWEz/fsCp+X+k0+F5gfGjqtKkB/r1cpP0pNRvt+fF11R2tcB
NC84e4a2eSffixZdRzsQhgggNjxrGNgCQWaTejHKtd18kmZvwcJlOzv/wlpNSNgBG97E8DIMONv3
458hdCdk5snYEOlAxtOEFG7Sxa8I+4QLn4KvQqQrSljSZlI7hmXy/EF6df8YB/9k525TEEq8amz1
iq76Q0u64wtp9SA3T7FGWSuDjS0cSzsNlPkZ3fBcPuCmu90FdWkLakPrpiqoPBvThtc9LjwAUzP1
uKdjkEdjkZtyqua5QNOU9IKwks6zZED7lN7Y78ZxLsdaXQnXbfS9Pr2me8UpZyokbC1SQZYcm+4A
l8lLfwwqkhpXuO0siPZQfFGjW4Z7yr6nghdOIMnpnE8UlqTbEE7N6p2d0G4zQN5gxCwpciZjHRmw
kU2wRga/9cNgGffzLcRYbjD3eDwqwp2OOlROdaz86+/Os0cDXCGUoA3Wya0xhnBkAq1JvaoW0BWD
ToLPNNjPTEpP5dw6wu+r0dSr3+/py1XoaoZ5YP5+RgxLixJkg2n7rUTjFqS7HZRJxa2PPoFAk42D
mssZng4p0Ti/F4tNArk3s7plD5celc2WpT2RtlzL7rIhEogEOqgwtDVd6tHr0eayxuShBTgZh3Fl
OzI9B07+6kDOB4wJqYEfJwvySK6MuU9w8CpqpCPfR/nx6w+9ItSFF3AhbU5GJ53T+/oS6AQvDJya
wHtLAJWnkF45O4I3zBRgcaxywHJO3Il1N29Mtg1d3ZPOJWggmbDt8PxVSzvzkWaVDDQqbBq+O2fj
gquYWTdAcUoUuNyrZh6QI+zfNNeoc4khVY4mkwlVaJLNJxi3hW8wKzAcyIiVSW+B/SfC04L9VTLV
mQ5pIdhiUUgaudE+r3I1vq7SK8lPxyThWdAhRImnUlY/OR+Ar7x83m4eqeLp11Pqp3kdwuTdrQyc
1iQ8LyVEnRTdrtCGSpnEdS+eMLVgl7eejhJGTZk1sQfhLgFV1TJWECjZSQgeyISR4K4+JKAlp+WL
r+9B5Ge7PePj9mDDXRTdRCrwgHxNfm2mQf91nSzQYuzIVccG4sNSe1W3SS9nIlEcoHnE7V/zaGby
wkR+SLAgJK/0l5zIzZC11wJ6ZmXbf74sbuwVVfOL85y7ZvhJRP5R5XU/LIqGaWf9h9WGQd3wIyiz
FLn5BBdQgwSawPFzKbFCyhXTo4+lpTIJR7QL0TH3+cpy338daEACFxDFZYOsYEP4/XhoblTmTxAH
TvMo4DxVawMvJmPORt7LyQu7vBS5Hy/8vbyDBNQvzaD270dRpyfiCBwe19TqXH1u63TFCjChPqb1
yrsWR57zdHrLg5LTdOXOrCzaOB5txkMwWTTiD/j1/vsvN8j5gxpxUx8nB8rdev+uVdtblRrVGxPr
cY0X8v/FmHjXF5AJeQ+F9zgLUhW2brmUeNolGCDqK/tQB0MnrwbPDhLCuQJO4HRp0CV2TMNnXTsK
Gt7uY0rjdGr7nhygf20auL893dDUTwVEAhsMOAHPAotzfZxJeGeswYr/4uo14rJrOxlqit2Lmhxz
Edm5wi/bVVR7+i9sed87iivaevEytzbnLB7c5DNuUaqu/koizRHvGR0owCrCZIFYIm7HwFO1S9Pi
EvfmO+JxyMPgK1+OooKbQU9g4wo+W92hJua/Ppxv5DertSIW5QhK99jhlTloJMzy9v8lenFUAveg
2pN39rPC4ZcjIbqdCAY4yYc2am7zLqR4l2nup2vqYw9CEEWi3ej4ySXWDONVDyh3i4QGr2mzf/tW
GFix4QVyP7BZlF9zxlAc2sPppDp5odtkc1afhD7LHSxdafcaOnG1q98YOGyrrAmRDLTCY+rZT0VM
wcz3FhEkdbumWym1p1h+CNKUJHd4vNLrfOzaS/wtJE4BBOzj0yAMS6bhsC2/YpyqCJtrGKxifMhh
50UeaYq5NYCe/a2c4WZry8zVXGbu1NkpXA+zFkM48AxUM3C4T1xGKMNO22ypCQ1R3HFUvsM1Vhmy
yhVqtwsh2Aca062jMy0Ed+ksU6w2vUUZHoSBNW/Lmx5c5GO/6o7uUTR0UKyxXLyM1qNS0ZbDBcF9
XVwHycLo42fQdrDxV6a5Ncg9sD3N8tuqw2CnQ0HJnUIK39dAwYqgdtpVB8fm0URCNm0do8fBsi9y
xcjmc2kEADuNYpOTpRgLDj6gZannjwq64MXLEVONHNs5ONkmRcDE1UczF7GgYfOKdaaVBqeBd+vc
zE+n3V9nAv8gqgljUOolUgG9Ka6cGM6TUay7Egh8VOr0S736prK8J6kIvqqV5uXYVaj8Vk8BXB/q
yLPsdpzGxeWLP4qhge/Y+AZF1PqP9eO0Gfhg/ojO+JFs6MREiUV6L0AlcIZ5cglcGPmad55PxKVy
0JOECj6lJxV2cxuu3jXBqYEb3zLEnXBPMa2M2tNAC3MLggSPDUaRg0rKijJ1mAXZOJDO24Qa2eZJ
EtHX0jRUHcgX2qGxaFLok3H21u/28eguHC22nv2IoQ2/gT+kxHqtiZ5MlLk/4yypY347tGuWeTD2
M9rQn9yp+d4UykHa/5tmtehJoaZWwHuQz2yNIYWH1YQf+uvV5y8/LLRyK4d6AKZ9SjNwnz3trcQh
+1CF+lcLmURdd2TINckDmiiTEIM/1XWwgpmyb/Ee5UHo3bpm39evQjS0NhKiamsTy8eeXLuo96Lv
C/8nLvo2rGsB2D0ZA7Ld8ZNPXs11ty3GvELYqQGfPqUg7y6UIHEg5ki1gKxtOmP4O2ADo07oYFR7
Sx4YOqsVIKERpE9BHsa0GxBW+kIbk7paecfScCeW2Bz2MQFsKpRp6nHF5Kns44iXqxVPxELKWkRu
1QRZCqym9976CeVucfm9mNRUp4gLWPHQpYdtEuctuxIUZ2DhVLukdDQLP/mvs3dmXhd36kapCR1s
2+updUNr14LHynRWVl7DeOlBO/rMIew2voSENgaUAbO3BU16zQDUBp93IfPHkxy78zxzjS+poHel
VK5Z8k7YDdnmOxAaxrKkY5lVo0WAuxh25Le2XHnHpmGJLiB0AgXQ4y6yUirBR8c23wheidlgYMeF
8NmvbIvHVR9C05dbA1lmk8Xnm2EVx+YhON4NuWvtaVRQ6hUsLLnV9Q31Ry/GYdD9pwLqNr19su9D
KIxGBMtOCF8DF6s5kwW8K49qdNcjl/nG5uOMvXakH6wBgJu8/T8W23moVpMWeqtoCPwIK5iGT1iv
i727F653XgOyR79BV+D7TURfF+moySHQl+eQspHYdbXcg0pc85eMeZkt/wgLA3pGtAn8m79YPuas
PukfBKEOm3/icuoZG/xH/3tbfEHAjDgz/Y1pmGzQxG5LX59HddAIjWvHanLNZlyY0N882yE0eH5o
VJWAZLvePGXU84zMb9T7vM8po9S9xpwgF05KEKmwkOWiCAo+kj5dYQhQEGn3AxuHrbEOfKflmOq0
uVblhlfKfwAu6oE/F1LTvPgYxLKjEgN5k3W+tlMFQgorqWj7DzHWEKc1Eas4dJ2ZELwisphcYQHD
G0GJ9WGyr+G6Fc+wjLJqZcxEnoDBoHqP+YQWhU5FqE2lrGGsj8hW2YQIUzv85XLFvnVKk81+Srb1
VuxQ1U3xivY4ZYa7B/FyWq+qLO5OwNcox2KdECc/pZNAUQly6COZhf8dhezzcwz0dvLYW40KiRVP
JSpJPEn6AShoZHBjWhpjqw6XSOwBsnutblJDH4qhQtlCK42Uf3P3ZekphdS7bD3dq4XwvZnn2xPm
GlKgK0wBXfzwWnAa6mI0SEizyOOgxJaDiZxOfu6vlZCrHHH+rsgePKrGSHWaT91MO28N+M34kYsu
ZljdgzR75cN/rSKbSiZj5V8/nhE/Fiq93yag/lE4MMqfAg9EqOo/dsakLmUWttCfGFDgBVLkgo/d
KAbbtB44oUCKCEJChVAKKnPARXIzWtLCwtQGq8PYefwSopczK+QImw0n9bAtaAlJQuUJZOg+tc+Y
GxSmGoyJ61Ed1QI5j1AJfv3SXBAjDyQ2L8zPwfcskaeJuIPR2WbTYwOw72Py+8FG1KTg2KBdnTGE
1UcNvD3kF+84yzvgER7nAPOhzbDMhj4RCF8QW07Cjq9dTkLe5e36b0mxqEIBbTFjghjZxWWgI2S9
o79er5q8Mqmb7jGswpJR38tZmFefMxzEvG+M1Omcm1g2LK8HuYMXaKkUjsD6JWT22AkG066d4NuR
y6FLM+EUlkK95kwQ/Fnx7vm1bMWSEGQCdJ/Iocw4hzVb9PTbtDVJ5sle4pM9cyRZnl7qy6zMQ7M8
iGtvcsXboXLxH6nclX5LZjktru2HdpC7gNLbG+85q8bj+bR09qVfXn3pGJK4t7RqhmEDmmPysLVv
Da4GfVq2vI6GMVbVwe+U0t2IMQLWzalDLgCZQEYPOUaCa9Fwf+BweLmDth3W2z4CuyhjnL4j1+0Y
DUJCq/KOfsBs9H32q9dk1IInhAjfRlM2HAMSqZzmlyYh4ub1eNqJR0mgAqkyY3URAnvDHEQJuXtr
c98C3Cfe1+gOfTbBwoNHjDEJnfRNDX8d55DgHdddKspu4ZIb/E0StAq3AYsgj3jgUxKE2JpduZ9+
D54blv/WY1FzQPBMzYnlI/gKUNO2vfNwO4gnVLykAlY3NQooeVlO1mkuxzXyN8LOvHsDCHPuP2WF
98tccPBGH5gv808UFbjNonSOlVcILPDpBi+8mcRmvsVYBfWf3tj+LMON+kB2uRU5RzEv1nYzHzRp
pLKJEMi4piOAZ/Z0itqzcn8/cWxcJ57zM8P89NaQO6e9faZprijr+DYP62445507qzW6fqVE4MGt
Imn4zIROgssmUiUe8iEhUyZcIBJZsWBzlifwv/oPYmoKTyUro5Out1T3AtAR9JVpU4WVFsai31gD
PkyINUWPLKA6D3pxvr50arWPEdLbkZ7MqKj4cUy30KroA3JT03gxF6QcFL4XO6kVdU0A7VabBsZA
qdNC+9z58luqQy2jeXpCqduTfhbmP9UyqyA8L0pLUGR4clb1K5jTF0M/hDuzDUUAuuo7o41xYuy0
4pQcRW2C8c1tD8wfA6fAlegrGaOsCIwBjuPay2TLkEvMdy0L9Vu/wZfLv1BgSoOjLU+T1ANVAAQA
4GPhtEop4/pteY8z+jP8hnKT8tm+4QTs4cdTrCZB8o5OxRKtRvwdy2I4DW8gClB1HfSj+A9C0wz+
ViRg78a7o42seKLDhwCwGkJs8Ovz9ODJrJXF6XxibeV/EAtniYT1jyCAaLa+KFWzYNOcByIKmMo8
tdxWywe8/c+d7bZADZjjViMaDMFMjd8c9jj1IaocXqh82Ut15195YeNkRMJH1G0Iaq3Pk9XOHusn
SxdZyS7AygRWeZFA/b3iwlFp3Csb6pVRIBG/ByS4vDOlDXewvQ101FHXNhHHmhK0e+BQkOPsI/U9
wl3EUFqzSgullacdovaftmiIPZPh71d92vidrpGbyDHx3rU9mY5aqe6gG/8om/pKqeOsTQ+EbrMk
6qQzp1g3DmtUotmsW6Si19C/dxLxw4YhMR7YXpyTrOdndzn0Vvci0GX08NWaTJK3XikXocvS6OpV
WEdbhaXJX7+dKA8J6O1D7tq10A3mK0nTC8Xyg+i9Wr1vOfUEdEwhmat73YB4A5jbt6IOqR+ClY7A
K2mxln/TMrHLmspOC2OPHrSU0qE1KEqpVLL19epPOaOU28PFDXcLINlICapupEDpBw/qHgKvNxcF
0v3bN/v8QKxIaUeYURbxsu0E7e59POEB0jFvpM5VcMVvBICOPeWZjn7bNNAm7JVRUYrr2MWCpRz+
6fLpghROIQRKDEihGlKy6hiO/S+gZKTIIpSgNZ06bWhPjIX4Qi2TPZ8ZDtnHcXl+D20f5KF+B1G8
RoBnYoFq3j2UjnohQ8UlCYr/OWXuKtTtx7uKQo/Lx1dqkTQGLQ8pzvmourJ5qyRMXv61a6P0MLXw
Y9OlW9ZkL4FX0i8tL0KeiqeQYxABKJk+BZd17Qs4xrhXXH6DF7Y5QJK68l8a4zeCThd4LcXX9on0
GUVF+f+yKydm9jDZNvvCjoI0obGFCu28QlXQdGp6K2rWSpmGdeMr5W1ld8zxkQAGE6WvQEnbwzc8
l0XhnXRh4k2thjLTkaCTZdfSfpeSufYvJlPPND/E8h0k7VeE6WgUWPHM9i7breH+pGedDmTkHjy4
QJiyv5G66LAZ1VeTd0cSqBFpZN0sWH3VKBZH7Ou5+qv+KOWRE7bjytmC1oq25xymtnNWbMIdnATu
p7ixAPCWVrRPOtsTm4R+ptzlXZ9tL/OnSf2sb3boCCToRNikxE2mYYoQtxXtEhtcNSsHeUmlHgy6
D+itejApjTi0qZXBor59ccMgxpk+iWkDlyxIPzEIlh3ZAx2BimMXvF+iC96Ne38pBZGUjkly25kD
aIFV1/qfDdu0hrpWmeUTykGtU4bDJCvs5pQKPxGoaWyAF5MA1FJCstpp+6eW8tp0hoDs4RfpW/aB
Nd2e7KLUfZf5dG0EbiLQJQfMUoUy0YJTa6sODawrbtl3+8/6HuQskR8OSPDGQf4aRjQxeemyISNG
nixpy/f/szLWYq+szXsTEvGkP6XsBPiBGo5f80fFJnjuHlq7/HsHohJEu0XU7T6rZQkB6P82nNrR
4uTDV5zNmfjzxq1WPshkBcAAy9oBu9VFurN7xMCqQ9b7xwzkyHjQ59+rnYS9Y/VKATByLMn1wS/K
UteY08sJcr0aELHHpixxIfdv0hPYbYnQLAnYkMJKXGPM2fgStpj8LQT7sTAad93KdKZEp1SR9mni
3rFjieyDUfnLuq46m0aYP6hUnuVfQ6GYKXWp0AOqLWuuj4iAdRF7Nv9aj7glPMxd6lIj8H9Yz44S
+XptICq6NgAjKvgfCBQ55UspMkI6mWA/s7QczPDgfov9UpXa+QP8Nk1eKAc5c13bXOD0qW5InpgG
kZqc/9xTkgWniJjubskx8L//dQ2bLcv+fIx4MprYWOLVipD5ujvj6JQ0JpqcHcjLqNXeDO/U5p1O
nYm0hkdcAqkeYTuIv/RoG5fGWf4KtcauM7rhAgS41To5KRg0wFGG7QkdxPzMgFZ2qc3wE6+OW7HW
VDmJX2r077kTtTcYf+cMGzruRGnKaj6KVr8/fxqmI2m6SzNupttTpV3l9d3dyT7u8yT6OJmMP1t+
4jWgbe77mUhq7MtZYSfxNTSsR/7Y3tpbaA4PIOsg72KEdBZRRqh/SMiThr5CQpJ3FmeKxtb+omCp
o4AHfOg8hZgSf/F2DUsU1Oip4B93VasxaXNiayA5LBAo56akvWWnXTL2ZvNHHgKbCxuh9ljeU60x
uSsPn+tXb+PeSf3AYBvP42+xPWIK6mqLsuvvRFrCAs69B4LcA2NSOHhe1RjnaaMR9bJc9O9ONgil
oTQAkJjsV82s3ehte51k4lFDtknEWr5cc8eR8aQWxilKO4Z24hL76IPbWWjlPlVBkCcZaNIBjQ+F
jhYdRTYD9aSANR8s2ypHkhIH0DOCAY4CjMzyNk/t0mZlBDgXDy4M2Uj8knPy60KAphIVPdGb9XKq
wfMbiKOwSEpc4EboLI5/Q0OuNXt9x3eKKyHzD11eWfbHhEn1evOoajteEL+e4nUQyAWPaLvIchfy
wYokNaS3y6AJdcCGjkih/EKv7ofLEKAs2sQHBdclOUgX/x10sfBbZfN2kc0O4Zlz70j4wqI7O68H
Hr+pBWDQMbwwrFelVFdEXYJYLpoOu+bQ6hAJlhM1FIvZSYQ4HhY0VAuv9e3Loed8dQTxf3Oki9FN
17CAK2xFBfc5oh339o46LxZ6fsiaXw8B3AFKoxBOLQe7zJRoNmT9+1YyKSi2qB45rLHAN9w/P399
k2/gt5hPhyBSIx9n1ccg1/2bHzK6bILIZp0wJZ2Mtk6jTJ69T8iFWzPUf3qV/sLdtH5aaSkZHPj8
Hm02ZarZlLMNEWApkH3bGOanA6E+8v+73Ci8QHsr88IdswirLr+RTZuPJZ6jdgYIiq5cwN3nd0n8
RXlZq5s2uJYe3a3gCmXkbTnFVo/DC1MPMJaZ7Cex2ILOBRYnBptTVx8H48HDzVlW322IsXiYm0Rm
vEIuT87mrSuO6FKGVQr1Gg3qm0Rp9SK0zS2dhdzZ8LOBM3ZXYzBaqgaLsSeCjclOnlyuCxoui+Mt
Lu4K4kad7MrIkA4dC8ndEhFITvxAA9mZfMyggiPMV6MC6ZLerZJtoSDGumQZLp/uOufLFi+oBRLp
A1/kkig9WZyqYwPZsGzOlUyB9EHTs/pN3Ev9EYhwSPsgB8d2BwlCGmq6XKXpu15J3ps9exBKJWmC
SMVrkFfrUSW1eoXnqSUUFQbYw0Q7MyahOsKNgB6ND8P4CoquXpKe6BU9mltK9hDZ/aigVleRYMMG
ESnoaN1C/il72IqGgxsTOu1Y2u36azuSDMz7002jR4UaR/FlEA2ONVJumbQzkCZReekbH4jHq1qh
TfGdE7p5BmivMBmP/vXR2BP3VrYQjnntVPaSm5oxqXQ6ewQGFSm7P8veGAAgv/+ecbDtDymkvzIX
a88mdqJUahn7xRIU+VH5rBU5+XZroYHMNetgfGngU81trbI9Mrh0HU2rEzS3qI6OMTkn5fpPYgsX
3gBZ2bzld8IIKZuiK6ek9HKtSb1MLm+kENcaNsnbHqArMjzseJCLtQiDaIxIlO4BK5Ftxoom2TWm
j0uzxpSBpaDYbqtZchSIspSmHWJNLZQyB3e7AjzieRNRxz+1Sv+2yd3JEQHysCLYLoU+em2nBJ1P
lbYjiDZNiS4jINt9gGQwBTB+HrsEOgFc03BsXyFVHxxD+Dd/8JqSRo6SrUgy1KZOFHjVDx/Uf0K/
3I2ZAVPtqgjrhPv5/9O5eJUeH8Zxs+UneUl42RMeo3rXB8t3EkC2HU9rXmE6D7V4pWDTzhUfzdjc
nwngVoBJ7qgrTCyKITpNN1hrnJwjR+KjKyRfiFK2Y4OmQ3yNtmGxBnlZ0R35lNoVUY0lzMO3g/19
vxQchL00upMqi9386H5cb0IPUSOFj9Ix5bf8AbDB91SRF68bOIX59oUpuuILDpsPOUiWcqzSClgq
H0ExUJAUU0bKSUYklvDZI/t9nBqekJzija8p8VuD0omqJgr9n3UyA6Ugu/PS4pioq/VTIOnhMISr
OzHs2figwPbgn3vXJI9tIjW5+89VAQwxuNHB7LXelDcaMqJji7PXBqFTqTGL7ZRURvSMXflI9zBM
brub5HlxY5BSi93u9l3bu7Um6oyn64ZJzpyKk3TgIj90lfSxVukKBlRQ0a91Nk6NnZXo9OEaLGh2
sdBfLWnxIJqQAFozafIrTo3ZyQVmIJ29rncF/Iyc9PC5cZruEZIFLW3EPd22paUsSlw+ULqkvRD6
x6vMU0QCrz8ISeCc2WnxR6/KnLWfwSvMC9VEOLmDL7p9mSb8+Xt5rVwXJ0JcSJuWxU+9E1H0UwYH
B1BQyRM8jYGmSB2CqOtmxqLAznOGas69U998vXASj8cnFI+Le5EX4mdtXLdfnhSPW1+rVwYeKu0Y
qHg0NIVCvcul7dZu8guSL35X9ovsbZnAMuKqW06A9qYqKcUug7W/+7gun2asbMYWR2E3kkqXhui3
3EQO9Q6zXRb1fee1VWOyZqMyUqDAtJ66yZpPi1Gm05I1AoHojudzGgnATN4YPXcIdQuJmpyBRkaW
estSj1/sESlbuMwAmoI2Ga8yil1atqiXIC+2dRYtyC4w4QAqN3ijk6J/++H9ggKgWNacXV7iTwQK
yJPN4J17bfzgzyE2U74o94HkpS6/fChYokIsdKkQy9ZwM5haHhBSjvHLaedOTA+galbIUG10IPmW
sIPuTcubWFyjghnBsx7RfEt7fmXIvWGTr8xhi2hxGLO8RtlGhLwRR8zZ9osicxsP8XNFyjQH03Xb
wWE3XdCDquPuJhTL/VHL71wByUkqe399qlJ38EVcuXTulJOp7UxbyReqzoDovORG3uy6GLILzPp9
RYNgHyn6YwzsWUNJEPL231JhSoJobJb6v6TghMiU2XS0+eniLTy4BGP107AIopdZGxWt0W8pSco5
D7TZynFYsYxhwM/MFOjykfp2zcJsdtcX5RJgg8iu2hw4Yt+x0oSel0obt13Tk7NqfPq8Bgf+8G7o
S35Mqsl8RTAu7j9X8B08ufF2xirTljf6J4g4xHJOEfAfMAGohYSzNsrY/kDa9TgJ189XJ8mPMHWE
WMxEvERZ6DRfc0FzHwpkRkr8QnXTjIJJrjPlDr3CnLUbCGKvDFGoenF8pJl42KfsZuYla9gcdoiK
bruiVw46qu3oCRcuaLPXtRgcDBAlqL+CkCAvOz6IaBU5nZDZXgx8wCXoEFK2ci/nYz0sdpS3aX0l
Y4REXT9yMknymkKxBa0HezI7nfdO4R+Yid77DMUIJB2IteMB6e8vzlfE22Ar5SzFhHTtpuOco3sS
LtoVTItyVLpFRLendVV8tZEsdCEl1DiBTAwA/Q8DPE2XG5zoRUbzsXvTfEUWQBZwFV2cXA/Wsxrd
un2ZOeP22xElOD7Px1gqR7K5GmidqeFhWKGSZtFRmtzdVTJVfZLJdN1Nc340F2pQJBpg0jEoqhcP
ZQwr5iQzF+0DjyklUfVyiROsCl9/x9CaEuas6Dw9aXVjAvGM2C2nV2+nKnUnDTkea8J87GPKQj/L
JODptCut4qVWRVgocn06jjd6l3kTxk+OUJJnkUrdhtckhQhh1/lRJHgBdGYpdOebglTKIQf/uqh7
fGrA2kJ+FdYZ0R1m8gtAv0Z1on07ur5EoCje8qvbSGVBuU8PIy/7dXbpx3x39CMIF11CzVt3mKeB
6EzyBJM0vZPUX7xS4iEmUDoVCTkVZaUgQhTFY4gY/0lFMiG6/mewJA5AV/3tk7WtHIqqdxFy4/qy
ikMYpefE8RdmN6r7xiLagmeFofJdvKJXAayZ46vpig0sDA8FZxLI6IkS3P+xNKoZ63QyYo4i3TdZ
UZGDjWFOSTB6thu/Cv0LRVNPeiICGw4iGNxt0T2L7LcEETkzzGf8ANJ4l6mhaPcPIrL0JwjmZrrs
qIN59ACEU5UEapk31pI50gJQ7M3UJ67PCLtHF6KlAFD5IKYTezAw7tFIfUgDr7G41MOPR0PTLxJl
9W4APBz43fwl7MIfMpcNXNQ4oJhyOfTYMoGMdL+9fJ6Qc3wsRZjZEgOfCdk3DiHzm4dejHXulJ/2
1DJwP2GONbzPe11pXH+XjEtoMafDaBlImewtBF9x2XvgyZFuNXfzMsgxfcabSTrzLgLCLxjRE/xT
PnTk5+ikp9yV4K59Y94Md98GmZrlkrfwL0NuQLv/CCxhzlj4++9xUAV/PXrJnfMNYZzHSqdhGFQK
sT15UJ+D5N6hpUJCstZ9eIThi7GDQj1pbdMu3nvFydj5fyTm4rMxCJETntEYHwR3eeDlTyhV3Gjh
NeGsSrz7pufw1qZnTzvgwEhtNwIi6VHJdc7DHFswS7ufwKKkehs3RLHw9b/bIrzJ11xGml25cDID
RHaVmX10YyYJKYtiO/nGG2ydrVwklmFG5QcmZCwGPWsYAP0a1GilybPw76NLr/ggZINhCWdJQUe/
tWWKkmTwR321vfnQTQxzKuRd2FFL5hqLfvgEwcDDp7QWXyYWtaJvOAkBQ6hro2pqGVyuevR6cfM5
uWuqZ+0cazqe32XWZd5IxYET0ZJ67rFNfaeTYmPSe/Nnvb/Id8FaJ7T8/TlX2M58ZGSO5f9va9cS
PqESF4cyU9+L7Y7Jh8pfX7IX73mVR4G1B0H58v4n7Mz/CTfNs6O3WwHsEA+PByQW+VJTn9kr/EBp
SVC5s3lWFBRBgDIacKNYtWaxsGmlKjJPhq1UCuKNrUNmHyVjbpINnL+HuXEU0lat2GBLRFK9aBN5
CxQh8V2wKiE4rpHT0qYxFKUd2zzaNjlT+p33P2soQ2J2NTMzLetBQuhaaZNSnwZKw9MeBdPXcWQC
+j3dR85qWxdZ43nc61owD9f5YWS2hsGezvm0IRrg0O9FwKQrczv2ahFCSGKDQj2bthM5fH7eUYWX
slugDiOlslhI2Da8VzWHwcxdWXuS27SucUXixCEvyevwJ7Jm3py8mlCffhTKKXODZl3PYJ0beosJ
xUMQNDPvlOgdJYMpm3zIeM+1t68SlE+O3Rpe4uYsC0IbzvHUFEyteMUeTEi38MF9s9LmfYYmJvFv
KVNJC+DDotVF4fo2VLLGDVeGXIGDYvIXfh3yhcouIlt+i+StYcChZ2Jwq1crh4rAs1hmaBCo48Ak
jXa5AmJVmqMaREfRf2UkKmGtujnqIkZMtykzRTf/kQEsUg5UDesdxfqGGB02sbunp3pdjPknxTuB
zUJtg1MIIZt0KyezRWwm3XAtBq4H+sTRAN/xPNPMMEDFcyO0F4odoajUuKPFui7GilxdUGOKFgY6
29d9S1+O58t3r8xddOpvn/6Mzddkub43B9TFcscIs3TBh36Lj9eS/E1HdQ52o/UCteYx0p2DYGQD
SGpTF3lJUtBnzuh45k++UIaFamXZyfqQqFQ0EkGSKUwb+t2WHopxkhpQ73U2gNoxaGNxGwANhMx5
BZbEsSXFJZcvb2W12zEOzXU+KN4mk53Ikgc1EZoxhnKgc5nBaN3ZY0g2S4KVlS/GkZePBwULWf5w
iwyfqOCUS8/1U6ijtAJF5EW/mrtQ/EYS3ipW4PGtZWqbNO/ZlPsxH7UX7x1MfNfT9IfekRdrq/zd
oZGc5lxZfWto53hRCsUN4wb17VD+h6ukuZ7+zo839MEuyIOxfE1xnNNjlRYKJAis3KVEgy8llF3/
zgdEjcV+Gp9EdF/qjfb+FwhTDfYzsSDHc3R3OW5hnQH8TWmlfJCfHyXphCEBBpNmoPBIu1+0rZBW
s1ZHZCEj8chOJ7/PKkQTkFVT2JPQl1vhLx8l+lBclSosIwYOMvZnvlgMBZ8xNByvN+e9NOP0h3uK
8/VLUDB6Z8KXPtJpuwYGtVJDwgdqQgGnsnayCZ5ajFwKexX6VdF1/kq2LfxDNrhcfFHJsktxf4kK
ye6FYJblz89PWNI04xF4fAJZSxiv/JBxJQR8s1h7gfxmSR+4PFomaYv6dytjepDQNYFtldVyHLuA
no9AQdvOlH1h1AOA12bogJl9NwQx+9R+tk7j97CJLrbGlWn0Sk0OeBsErpo9ck2UW/NxEjfGvcy6
Nxp/KIYyHN8f7SkV32xGbAkyL2HnjiCe7fggTMzzlE0zeeKHXZiZghrbMPD2L23yLx9DOph+6It2
Ewpr+ZWRba9U8qqij9+mv2IBoEtBi6xPY1zoUxaLFDH5ioU8eX47otvuRQwVbJHz8XdnFcC+qkSo
5mMTG/EHAFmBaa2lRtNzFfyyKLpxj+5cT8S31rc71tdEjOFhzywvgRLB4wJHQ7EL2R/xO+o+Fkdr
BEfgAqoYg5nUZKG+/aU9GXCWF2ppoIoh90xJwjHFyikIZ4kslAkahS50TMOV+gbwGqr3yAPDrk0L
dGF8T8UAJoKVAMLEhH2ohBfFd9+PiS7qX+qXQfFv1R3n6kJWicndij0nDP1pRpBXuaJpPyGygYV/
OKUBYlD768DTg+qWmfusjs6a9mYl4gl5aG4sNa5n2R99H3EbEKb5ij5/rwPBhhECHmJIFd1zoLye
SrQJjNDccNjfF6X/fAE8hjv26lSzH8fIbigzlx5LpeAeaiG32fegy5kuJU78lzl+iNvWFoJe8+8w
NPdh1ZVoDAMM6wZY3u75WBpXudVM578pokmTiFmpJB2yMV0Zsy7fiHMmxoGii3SCklwcw97pG5Et
VHNvJZ/XjsGKbxEDy8raoW7uOxyvJxox6J66TbqfqwXtyXloB2nUe0Z+sznY0/mmJp8fUhcbOXcC
eMOur0P5F75DX5qQwPqnKspdoB0U/B6KKUXmLLktN5uVTPGOE9IK7623oVJvK819iG1+OQ6dGRGw
ra/f79SN7T41MyWw0t0ML8vUQTCwlaJ1pQraAW3UFARzn6JptLoe3y/6bcVV/6LRphZLLlPXAGhN
M3rGC8uLJh7/RQyBuuEsOllHNdUCmPfstEwHN0BqiVunzSJ9wZc5nHxT2J23s4S5VaJftWJS1GLa
yyHdnYa/QcB+ZygAxokBc0qFxQ7c2Ec4FrXfAyW8BtLr8mrtEXDQY7sOZDjp+BLJhdEPTnCv0hY7
yTCNj7AgTTHIP7NLpv6wFEHrayKd3EWl9aaEGePZdhObL4KJKfyZx/R+thCeEY+kIJu33c7AssKP
UzzvbZJ6tnIZIpDood4IgoEIugDeORJtiQFwnXyPtXEPXrgF3a06u7Kp/OkG5m8tOMLBh9zLfP/G
IvJlfW4im5+6pHNSM9xBKPJMIf15ViLy7KtpYxGfhETJdJY3OY4H1qaEaTBwyi47rYz3G8esEt0/
ZWxMF5MCqs0XnusRW8dteeHchXMUUgKw6KFm1iE6CbPZUg2EYAsJ0YNGQdJDQqkyKUeq1u5U9eJi
MvHb5yjxJyzsKpfFOB+iRZDXjrvpe7qB0I5dVZtSkmpuBXB0p8w7W0D7U7g2gdtChyIJqejdUoM/
GbP9xXxBE+D9YM5gQ8l1+8CZFHKyELaiOxkI8/nB7RU6k7Vyjmh6K2S9TcJgePKboYA/ZIjjrWxK
FKNYJhaGgUMGnUl/TYsLkVbIfkeg2WEqHGxGyiOACWI69hPYZ6TWCLAYjTucXfgSd+4ZQlIPJN9W
p9lttNHncRVDCe65EnI++TjMAPDkiBbf3e+31GQxdww/x/1+dPkzF0EiixI22ZcjICMwvyDb/o81
KRTj2eTrZTNFT+fwHfysv7cdBPkuyIlumXe+xcj+WYAjpjE91sxjCldLf9XIt1XXNBgtHqJUdnJ5
NoLjvWEOHcGy0GZsRnpY5ANqpCY4mCw1WDi+6BsrozucK/vLP7vjnbyvx0ySjsqZk0qaMTJR1ZDt
1q/HhMe61nh06BmV3i6rQ72ft4RIGZjzPwAqGkSJdy1SyYzg7dGhQ0+5kqZyvBhadfXfZXUm5t5c
aAUFZNi+FiB0/NM06ZsmAnk60vJBoZNjf/RspTgW4KJ1MeIe5KQrIOjQmaUuJXmPcgL4q9Bgk+9p
iAnT6sClE2uxUutoNiCDs131VZtcAFXvml2pDy1koR5sRD6c+zpnnMhRL4tO6murtXNOTrDSH0Eh
azmdFD3uEd6rNnVyW9+ONXjsHcnw409wlSJfhuiDDNmBR7TrMceQ3oYhZH0J8NBWEY4hSqp0+UwV
/CJDOVZTbihrpFV5qpdTRcTSiR4hEW27+8APWdmVCDgX5v1vKOoXJq8HUakyqjo7e2KU4TqNtd9O
zTVFdh+dy5dWYxNis0RFe1QtGQMY4RNA+Ksojsf+RmcBzSgirEu8hf/IA1vvPXH0QRBeCR1zMcu2
AE0/9zfeOlrMR6u6HMQ0qAJ7iOv1CGI985dFsnw49fktlG2rkY58CqMtFEyovHxBPmvkmB83Ed0a
Vbm11F0WwRPzz1BmxCROF0+fjDSqCyuJva/NC0W2wXSVXf7vwcP+1T1DyLxk6PlTh724wurXHXaN
yVUKf39bstUBSZfWcYpTF+rfOLCtljc3acVMZkOT2D3vSuJcqR7ijUzC0HjDBDXZlkFfAmj4Sqth
F15uRzWyfGKgKy7eLbbgX6uH7p3hZ4Qb6JNKBhx+lz0LhyheykR4isup2pTReUrvm0PFSHDl9BUo
SoQwA0V017JtbqsXBXirVS2lY8nz6uZKWYORdMn3G0ewjeSKm2kRZTgFPSNjMSehffzQJ4Tp0zjP
sWGndAWAAr20T5YH2pVPMbL0dp5xLQZLNH0ArnGQqTdLmu8U4UOxv37v0DZcBjmpg56OmYpt6yfe
Q+UHivR0+VuuHSk8dHjKtlHw75+exxw6TLh/nCOxuISl95zg0x1JNRyst8DpWFCzwK2WEsDpvW+D
/sTSm3/K/+n37lsi3eGaP2Dt/8JWWlnVcvuGQlIhht/WKf/vVTPB/opZWq4HWMzQEs4ZeUtwBU3c
nHkrkb3EWTgDIDVSjH4LNKbn36V4PbZsg9gNTp8Qjyn/6CrY1JJ7S0qFnMtGHpyxZAnCYBrv2j5p
mjHf2t4THfiVebwU9tkh7omnbqnaPERdjnFCcBXuTyAzIJVB9Itw2v2/n6XBOYG2Dq36tAoWJnEi
DDleHmoOHYxnMmGo7hLnSRZreW2ovClZ9jmVtiGYJawztlH6nEu6OxLjtzlUVPT02EpXNaVG4k/b
ucwk4TMpc6G65tXCSva8d6BUR59W5qIcmrq9tXzF82yY0Rz9YV5VZ3DaFJw2IAShR6JBTHxRjHx8
RqX/MOTKBbFqpEfeGqsitSd4blb8DYpOm6hN/K0Dn2OGGqBmpofAzZ/IiioIkulNNUrk1Pzke1Ia
fBjOBZDEWZTQRaSaPaZOtvixPrAitLnO42SbNnfmvnmLspeRUdDj96XxP6Ckybr6hFiU6fZ1OcAF
dUHz4HVyVrGj31f4992k15HALZASfPR+JPuYEh0VaPzhNxt4/FXahBaRZkygQENyWvNcFadUilST
mI3Fm4N08wW34MQPn94OnRp09UhJkrr30bXHA3uHaJpiQATLX2bXHET+DaGQZO6NDzAL6EPEMTys
Wk2+Jlh5IPDvr+V2M4kXhN0OY2AY1IQVljdNhb3xnpd1FBMQy5by6m+Nz+yNEg/LMpY/BVucUpkP
/rPqPdOqFmKiPAyB5pLyFasjhUtdRlVkW14rN/ESYQiBTgSROkv/qClRS6aP4vHEwun/LH0eGnwx
xYZxb2y5ZC8gKqYYBMKyUHRHAmUhGe6kAS2IQAjvDvdj+xw8/lnI573a8qzUAZrHzk12pxaxw2Ms
HKO1k/gsDQv/o+l8pmCwDrgkROfWT1C6NDQqnS6vCMmEBuGWeRQReTqlha7kFX6nZ1Ua4+FyYFK8
e4Q58Q6LpSyXVq1bD2BibVUDOOwre6TWQSix0oV9i4CsUk5TvbuaitLPSNq/SmqSqa/CTiw0smNd
kG7GGUCokRtmR9atJo8yzJ3mQ/PUrw0a9SId0t75Jd+niGZoV/7c+cEW+HhiqL/Lj9wId4477FVN
XZ3PJZZXzpbbMYr7Tvm/8I1OTLLivJb2vQnMmOXkXiZJdvyFH5Z3gOVP5ZujKaHl+4jnUXypKRoF
b8FyTE1KVhMJLJ72XSEjcx+C8HVdVxm4JXp7yTKhCdMuXr09gefHw4GX57c5hlYgEhgbS8jixXFU
o71xx1gK5jhIiD8+X+sArJGJI2DrWYStEreErM0LTaWnouv3tfqfm5HR0yZKUCxPsGFpklsNhvHM
SATO+NlDREwqs64Vj9DM0KfhYK01j+5F10MXLNIQD7p1lRAOigTldn4o408bbg5O5My2O3j5FsAV
JDch/dRVvcUYA/89APcZpMw76A66oscgqUsnuwmLtQoxJpYUrlIDx47lIgmQWEWUUYQEQ4VhFDfF
F8iFMHgUBSdBvSy5vfW5h7o0pjtz/+E1pxlj0ET/cGpNFn+IdUsWu94Mk72pdsbGdq8/MgKRPzaB
lsXZaVnS11gt/5rITxSrRbxkO+JIOXgvEqEXmoVF9IfuL/DL5H71HUQQEjaqK1Fne8cAsUQhJ5bW
wnUL3x4KGikJp3VQL2PP0+VZEDR62GIi9DHoQNRiRKbDK5c+jlptL6Exz84km3eTgZZjWQ6P6I8d
iuyrvK5ToXiU5hxzAOkFk1UQXcnasp4B98qSB590Oo1zAVTJ5IEo4/MhrZy5/USbIVO/U8DsSQp3
1urKlWXhYsZbwQJAyvRyECWAKTX9zcKVlgBugJCG8VrR9cAY35qKmNaP7KsOLGPAVPlxh+rIxgjv
4k2pECKjl1LyEhNceVU0e9qVWhL8oX3cMUY+p4k9aEIVia2hStzSbWmSmcXBogxIhcf39og6bbfb
7MZXRhwgPD2APL0uOWyhFEkNnC7d8lNdJXVGyGOaoZFgyOHCarSq+3/wSnUvorxEyu6MlOX7tdQM
SxjotXqvHX51qABO0UcoIMmdeiUavWlQnS9nk969VREGlnt1vPZb0G0r19WS/oC0sveSrKSQU5jT
7VaZu128fOhYgW+0Cgs3q0im4bHlKXhx0x2jPi7VPyOjMNUvj3FVCeAOrzK68e9kHuMbb3j1ZGBP
hVBRgP6uhEahTcEyFoJxvZ0/wNxH7hJykaFmB9mK5QbGQm5EpQOW/f6XFPgYYRyVETYQjTISBJ16
LeICZdwZN5TYHPhQKNDyX20Y6FBbAOugkvRSrQ3qOS2gIywNevOlLBbtXRDZ+Dtjf6y2GjIG113Z
smMGgNBc++L7GzOvsqxpXe8ibxQw99DRM6rDnWLFHznNEWNBMkmXJ4dX1V321FYQR+WrcI+aUrg1
/WuMTMRnYKEzczKQk5iEzseR1TTHeGyStOIYSz0FIPQjAEaULBK+5YTI328mMw1tpvH8ewLBRCQF
uOnosJqLXvxYKWQ25x4XSns7QsGXZCPmiZ5leYbWVUJzrXlqtXlEqiQEPM3OjLZMV2YjBS+vWEiC
FFZVzrz2nxBFrL/8ZYLE0TEtoZjs7g6Bo430/7Uni7G4/EneLr/yCetlodqxlzFn3WtIwT4hBCMI
oU1iRdzNmcwnRVCfZwW8ST+zNDqTrHNa+DDKp0cugE2YwzTlDhQY5iGo/8gx5MFTgeLRVScjBIzh
AlYOj5QcuOT5WNDtDbWUueqw/tY6BsvYMkNX9p1lyOpGULOhDgYxmuDkLkwnvo+CLMw7mxnvbazE
QMjbyHjrMxdzIMAXa6IfYbos/TkdwNMxe9RIvznkZj0kUWgMQHxnJquXctuZi5LC+1JjnL78hZZm
UOSxp6drYcHrgFFW2FqMhhDdUZFqzqbQ5aPEzYDgKPmTmyHAVF+d2VGV4tLqrtVpygNsoefsXNIR
KjHyINjzFUr5O1rQL7htfJ2w+cCVf3A5Nn39FxOOfRemkAFbqkRsbI8GHJ4iOUPMQmCmYsV+nwj8
NVy+bDXByixBmOYJnd/xDhcTcCYL/ryEZ08BHE8SJLzsH5KbIqZYzliftQ4QxcCuDBPiAxK/MdfM
WiDuAT8hTJFqQglkMzt1QTgOlg5L4O5WUgjek+oURQHOzaHxVqVBFcWI9IKgrRGMyrPFceY5nfHt
qgC4mk3gVi5HXaW1oGCCxgQ7R18HVFl7hxJLPsallpINTwfJ44KlB+5vUdTVjAmhciW9hkMOw6pg
67n5Lf7Wchm1UWhLBRTi3Dd3nOfumDwf4/XdvO1mPqJh9FFVrluq2TFPClpUGbFVrYykv4r4TAbs
XPHhCLNTbk1Y9VKEnrnmyGo3bKn1xMbaLRllnqkboWSEz9+uxxo2wH8piRBip+qHT9e50zLZD6u6
TKx6Or++MLkyUtQ4Mmc3mVgmXK5cA4LhiTiu7DoLM3QE16Ipau1r5zdg+0Vx1Q+D4hNJxQmAlpMw
dmxjGvojRmNLWsKhtuCPE8fcDifAtzw8nlFp8mM+hn67C/gtl8z7bcqjMDVdy20KtzQ3l52DSmVz
KVsCcbYpK66a8rM+T7r0jVxbeYkqQ/9HSPXO/AQD2a7hvPz/zVCqh5frVZDyqp4X4IyrX0viP090
VRpU1yQYIupHKSRWkf4llJ2X/r6ZX9Qu57+/IQYtijbfKhYT/OMXOkkhgdbO55Bj+B99h+31BroQ
d91L08VQOtMnCj6BRUD78mFAxXhijTrwmKRd0QCxTHcGRCUC5cLOoAxenxn4ZCdMyDSQAaLAjk+h
+IWXZQkfhDhLuQqX3Vm/C7t33uX6NfY1K9mwelVPPQRPSlijne9JkQlmkNIccfXoHLUJIJms5EwP
UM+YHLU1qKY8F6BzA+T3uJ/LsQbsCCc1OE1tU9BfIGBes5KtCcTPvnff8j5qTg3gKQBPar7J6vCI
ihJWuiB599Xmpif16+oaAJUWU1yAs9LCA1JBZwKtBfuGGGIES6xPkWFBNPMOF7VdxEr3VgV3Yj+0
C4jaEnUEIYyksfoUvy6IYOL8QKYXuTBkNCf6X9iY3OaaKNl7LrSm/qgccc15wbFehbFD+/oBahNF
D4fyn1MrjSRXtjbMvmZSoaBe6bDRaRNj/XVNVSmL9wDYbCWNIKlZZ8OFbaZ5IN9a68rcXjZVAD1l
zzYsauo38mN4jrVUjbKwQfjR3J1sFPPbAFrCFdUgXVDCw67/NqWyL1YpfyH6yVocL0d2/byVAu6T
h1ClLVoWY0O3i24t2FTcqKHgR2D/QcUmucGuadAznJ3lamkqQlCGX+QHEm0uVLbbcHMutwXLgM1W
fUvy5THRAHSsAmFwExNFGoKlnvuiMP25rgRErLbOYfR22S4it56CikRKeHQlWVnzj8fbzeM4pZHu
vtnA8WyTTU4de/2J09ll48dcJ6LCTuNCQL+Y5Y+zlfhUplMm6pS6ax0EKwRb/DdgzEeV0cOH4dbd
GSfwQQYI/LMKSWWR+8vdPBAw4jngflNo7X01bLiF54uIVENv7AogXvvr2jfr6wSI0UT0pzCxDguV
xy5elp8FKx75TMt0SY8apynHihwr0xCdzBkqQfLC4EQUeXTPC6+R0i4utaIiV5K4aubjgStbigS5
2mtLuCJ1Fkoyxk8Wl4+ED2sL8rYzihSwueUm+fwkVKYCS+2twV67XsYQA/IgZpPeV+YUuIwVqXiD
WBoltSj3w868Nt3qYqKdYru93GtLHJEZBktkSXt9txcxm4m/YDXd6SwGBNDsRly5KgjdlrdUCpJd
WTOqBECDdteYRtppf//Ob8Vp7ARvDo7p+9s5DIIdPlhnl5e87E7La5o8dkPhantvObvDCNrBGwWl
vVOoMPUfmHaWHaVNG9qPze8wuHOI4eNvEmKdLPQQ1YKPzirNv25ghKCeBBlOBrZWsjWdIIbh2iWu
kmrv3gPqW6VcsUV/SMaBrBIICVOt6bVwyzqvTUhhXFwv0+pBMulSI4ADmkudSXaWDQJyN6I1ls57
QWUWoEPmoT9JCgtbYOXCVb+6yrNNSWMMvsxsGO92xNoOgL+PcigwRzvuOSeRsEJXxG3JNlj4KYng
Vb+vnyH6l4fT5c2yJM6MLUsbmEcgVXUQK/8wtQnyrcxDO1DC/PUZRwyMa6eB1+7c9oNcEm0iUgg9
Wm1+ocvAy3XvUpMM7/9FlSDEv7AP3OOgOo6HYcF37FgvFshaviQEdRPT5CcEMGiFvTaFgmu+C/Aa
U7QQJfESAcULtjEtLqyonS5tyRzE9k6lwmOaRuxkNw7Mx8Fe18/ODtpDxm1YJiclsYGcWBL3tJOE
7pLH+fF2ZX3BMFl9TdQBJFnG1vvx+51oNN1g5PXZJZxKUe+2VQMSBd2/8w2P020NCloiIN38WU/A
Fc2Wf3mzCjMBnNF1ZqBr+biILdIHHUDZzZkp2izmtdSTl+z1MxS6/N+g6W0sRbWmwEDiPcs8zOxN
KGHmJiKv3JQQ2ggyaZxInNA2ES7lMmktj+Z+c3pbUAtIiqfhBGCUzsktj7BKCZW/0rp+1aZSaqrs
NPjhudAhtt9kfenu1zeTEA89Lf9lviYOg0q9ly9KPBhC/ZWxxXXA9ND9aL2/CYhjjgLGkhQX7vdw
4zTxH59Y6e/EwpfwLSB+WuBQCfhWXt6nbnBTmbxLE9Z+IwfNaEQiOEL3eQDK8c2oOv7uhOIctM6h
uFWOrucijq/FDYaKEHVU1V/W0uvAfPKv0nNkyHANcMQp5QGOJa+n1hx2YE9+0rpHcET/xN3r6FUO
GzUVX3D90rHAm0RwuEGt+E+1ZtbU9ywtRhdPhJedIfCx3HBMKTMwX5oVDgG2NFvunaYrsW+n4HGV
L5vLRsWMsi2Xee85EoyZwfswOwn/payMSMVYIL7GvWa084GuFA6fgo12rUYOetr+XaWGYdgg/nc7
nbj6Bu4P+NW29g8oQoeb5c5QL3TjMF6rzkOYRGClJdae6jiZWXHz59wBCDx1qnfji6ckgZiN083o
oF7Liok+C2hwfeOffQnQrJrb+fmhX86wq3JsabfmoRD9j5hH3FalLnV6cZYjIPQL7J2tGSh1fQyG
V5Mj88NdImHAyB6prHF6hc3E2vmx3UZzndVCVayr6wDawJaQf97sP7GWvj8qJ9tNQq/+58T/YViX
4Odkr+4vWb0ZLPdcw+a0g6gnigBB1vY3V5ckYu7AzlCmtr+T3aeaa2UkRxz/i3dr1h61BholdHf0
Y/ei01KIGulxCF1kmIjljD00lLJ+STg3SGxNsatH4hOzLk1uv+WDKB7FE6YqcE5rv+FT2j1tGKjR
GXYIkKHxqabIucBdPWDau4rSU67/0KQyP223SJpcCQ7Mt59Mec4M6TPu1j8h67Ap9R9qROQKYDNL
oyDWV1fwxyxVNKNwg/f+RMXhSO38OBlqCcsNcSyvVBw/NAqbsUakL+pMaR/4yJqm9iXKwAePA7HE
Umrd2qhd1AOoSsEcFC33T/ooHUsAuuPH7ro52NWfls4k5R+bOKGKOnHZYhLar+RMkGygcFFWYjK1
99M09KL/Re6HmInigyYW4LmOpSGF+oyJbKipVueEm5slHypl0EhOWll+pKXkaZUcC/8TezxE3p+N
DIy0hSLqpTPQYu9PpejbH7cZsA9YfnYnSFnmYHp5xfTD+GI/9X5x4bsCdhZfy5k+Y4L6Ud+VFiXx
dtgjLhFSvouqJFgrDo/BB4pXYNzfCitG+4xUxFnaKchvOj6ZDKdGrExBujHUY1/sPLzNB0QDSlEx
8L5IC1BprkBOgF+GnZ+Tuuw++4RmLHIDRBMp1oiJGKFFmtQJmoX77XALJ+C2H+8nFtrPhkrQ01Ak
By5+WK4p97kU1uDLT1nMWJGVrzW2vg9Ro5Pod7cteTTVLq9+lu8ptgdSLnrWoynhPhsTtXzm5jMY
tILICnUw0HkVGJE+TaoRVk3OPAn+6yTykBYjw+hFn6M1Ys4DvSygU9AoPqnamqvy8F3IXGp0auHV
dLJduyMJJ+vCMtr4ZMnh1hFj9QT82lNWJwK13Mb61b9nRLKFEkAu7XpYAipO9ezoNkD4OqlccZwU
7GZp8530ElvGlVjoRGEETDiYI3sqBEV1RTsG27UO+FW5cwQSps2rLVJaHkCiuHRDd1r+VJPHRf55
AgBeVC84T0kv6T0GiEd+zD7tqnWSAU1a8mbVCd/SkeBRGe/0CQkgrLzz356pym/XzR9YqT7qFuxt
X4jyci8PsflxEIzzNzhfymHKFjYOPSMOq68BC6rh3P4YBul4DmiO6cc38AR9zQm4LNuBrnJcmlBb
62+K6wj4JKPWfMSvGaeRaGN5tKtiZ60xbVdAXy386I+m63hMaPmqrLjzYZhfg7h1CQnXxcDd9vvS
yT4ams9KpgSSwn9ah7iuIM5ih6hZ7u9UrxKmf4scCM3K3RMiNqQP9hPw8j1+z6OY8M4eFxB6QXJf
AKME85hKJHR8JzrkJ74a0W7G+lNcrc8UGWioMD7GJmYX6wrJWyesP9u6C0I/T8jJkURYv1ZA11U7
rQCo66YfrKH8snVK8OEJciijBEwtAsT4JEYV4TLvpmZi97sqZ/fGd0iam9It66FNd6B+UOqNp/x6
ZHiHophFGm1ERk0i3y5lal0bP94vbyvdHsIErI8U3XgnUKo4SfDb+iWW1NXJvEyb4o1MNs5VhbVF
4ipg8V3vnBJ5ocdyt/pXvkq4M4pTgT7/bRuF5+m8OXYRrgazHnlNBqcoRq8Nl2X/TY7V0RDPWXhd
XnokolYfPWA8dmKBcv2hg4Cdi6bHWQVPPmB9dLav3IXM1FZ+YTUyC5XtIJBUb2V59zbNNzjxqLys
g1eqlMZvhFDZK+cYCNcXNhlM10kqN9D4297pWGHwVIVl4WpJJCfwHgUJ03qfV9rhLcKk/KqQ47JD
xJd0N68d5IajHATb9d9MSUUmeSUoneIVpHtWcq8phC0z5CywPPYfwjeRNTRMQJWeTNjDMNr5N0Ls
rQdlh1CYHXTMltcF50eyEXnkXXoGqvZLqlKnGmmJ5TKKkQmkHwRUbuMXe/SAhURWJg9AIhhl8NW6
6yNrnxzT2tLAFtIYUeXsSH31pDlRFFlar57CTbNJu7tE/MUvP2H45h677SkpkOceN/TkYPPE6eyo
IXtqQnZc5JmEdo5JmbguVVuv22c6OVAJOPtoi9aFknqGc7L055JT06//VpCyKH5gcL4gyttcHM3q
2aB09Nu9gVUVXZXDBAc5X1d5Xjw/k+3Djm/RzS+6zw85t2QUi1NX3DjVmrml8Fq4w8KMytBfqQBI
TL0osdA1X62Eud0ZZq93PhNU7rwmkLBzKltaDuBQ20rb2dH6EQ37GUuL0BhreoWRJexnWVNsaERE
PI8mVMC0LL0SQ8SC0OKowdzCx4qdMmmC8WgEkGfktzl0JlGinIHUR84VOOTQ2lWr4q1iweZgUjgd
7Uvz0JnQmY8Ik327OtMRu0fl3U4sJBrmf4tu5U7OrZHaxvs1qWZizyq6kT/oOJdgdt0t2AiIuvjl
cY7Og5ax1fNdwDI9rrbNJ2rSJZ4wenOwsIxsIFqX3WRTS0XvNEgFaMRPTzBTabgJVwPvJx+xL4vW
Xo2fU2h2/4kXk8A2R+S/xnOCIqFZUtjY9tIo4tis4BOwkxv22MuhsZTiKI+/uDkExqAvYKa4npCA
C/fAx5zyM5Gjiaf4kgQkSrWnuVHMTo67t4Xo4RoJdIgK4yY0E1d0Sg0r6AQ215ge8hZxWZG+G7vL
rPcw9k5eaFRKyf+jwvRlAXZ7MX9t/Ydv+OWQuSComQpMUvfQeUCUHNW0QgrE19pZtscO6Z9jFfKK
qU5E5SN+RzC48Kn4gqK8VLPDqt/m8n66XLIKjW8hr2svYAkH9onQWfKulnSHH0sPnj7xnw7Pbvdp
Z/yeqOIPMQFoayTA++u5SEyBm7eHgBCQvzqMQQgFZbf4bVa8rbC34SI1Z72R+6niVhWJs05xez3O
idSZosxvHPMX+hEZ0Z3JcDyppi7gJNYmLlshMekf+eMNMrCzgcEwYKFvAq1LOubNJIHcUfH3gdPL
umgU+cSZbVcAc5w7FtOwaZY8sprQzTxCxNbACtEA7M001wqp/H4w8ujx/88gEM2LMtbd5pA9zxe3
siQZUnvYhuL6WXw/5u90pe4e7q56FCxzcRelbrZ7VADKhDfOJM9YRW2V1i9nxRGL8H/4ONzUah8F
tQZDFQoGwG0N3rrliT6JjFnb21MeLjlDlq/fxrdo/wxZEV+vk5qFBH3DDkjQTdsEurw823Q4unm9
vizLWiS5jIMr79YaVugAhJ01HaJ4NsSi3lNpbKjPFhDBsfPiiF8RcwQcV61FnjdnET+1eWjMoA4h
hXfcA6TewBhjtyC4P1BbZJriWoD6DuwwruCa03qpgr1EbtOJFdOGNSaD9i8tkEsVO2W50Rniu/Q4
ruL/03wDYeDdqNbyp3DDo7LRQu8Pz6mVEVjLVUjeV6xQ48WZyg1JPm/D6s2WqM6qUR7A/IvUwBE6
2VvWF6eFXQ8MZyTKwUfxLen0rtpLi75xu74jmmVtxotn3J75CyO1FLOUz/Yrzyn3cnv8Cjq3NHwP
Nd4nc4/tH9zTtrfwCLwRkmzvY8dCHE3FyZ1bqX3vYgtiXtMuhCtlLI4KSAaxn25mSsIYA3y2Hc9s
DiLs1ujlQkSe8qDU9EKfHMQauu+9U7sEUYXWeYkUfUxeKlp8zQEP+xlsMLuwcRhpCaojSaG5Xntw
ZW+WclN8tq2uyHBbCTnT6ydmLBiWJVP7gSfLmcn+UkZ6Qm7FHdnkSwhhQ52q+Ghez/tTyLHACR4K
hZS1DjsnPIr/H3qhYERPopWPx83O4gLXPt3rJ4EOOKjeDYx/9pq27Iz+EsVPeklJ7JngpvfYmGAR
9d8yohs+4h8S8cFOf8KgfiEcEwXz4bZIZrreXojEa6SWSF5gzIHULBfjCdyWb64/K2cChe8t9Sfw
unqL7Il1XhFmDPN/3ArF72LzGQVtymt04VgUwlOTA2VSQOC2JHFfAWFo3bPTKzKglCMPrexn0Aex
HE7cnTVYlMdL+Lr14CZwbTnGdZCuNf+7KtDaMMztC/YW0nhvOe3aKaEDFh60Iaa7erRrwyqabXBS
vlxBb86Pziah18tmFdnhClt6H7mhFAAAQWoGzPX0v4aEbtwXHwdy1bkg93oS1uJbta4CD4/qLZyB
dVJiv1Rt30ieuJD9AjTSc5axWtcjUszsLnpot5w7qdLea44DwACl3Ze8RP0ZCqS7Ua89EKxs77u6
44ePdfOB0BFWP3kcMkmWZJacjg2/xSXBuG0jzbhJzHs5XHudZBYzoEj3q9rgvltAIv+AisOJ18Jb
Me1PRqZxiC1MUmaf5BeEYGJxGL2PedHaCnZLxH0+2aI9MrQDXEl2Vs8GBIhPiQNdDtCcnxmsW/1S
R5zE9GTy1UeujKVsXHs43+ctM6+cATDRVoXMdGT1nt++AAZ09UfThjGdD5belQ9dRA10BRbhFXzZ
+ayfAruOxpl0FYK/789hYK95a1xfo6kBniYNUhvxB0zoYQB5s9NABihYbrUkFvCDnpKNUr/GQPnm
QCMK8SjFMvdhMP1xvrXFIyo/5w0Mzps8jd38V3aoHd7PJw/I6Dw91Z3QeQF9IxpcEKf2v5WE9tks
pWUDA+cy1a9IVC6iOla5WumrC4gLVHaMpBHdf0dR4dZgnD+f0UcHrMruCn6t1r7cKio4nbSuiVBe
WZAUxBq9ZZDyprLZ9tS6mchwTPPmHQPXVZz95TBKbVkxh5CNj6lw0zS8hyzG3oJbj93OHEf0Ouav
6xDdt5bCxHvCaNPxYjQhdGhBuo4uj75dT6NyL3TdsatTEO6V8MS+s5YjiDevWOc4UVEuW0t73iFe
6vrsTMXuzZ3NnN01mGIbNZSqFcCLSv+2NCei2nyaKLaOb8NKtY4VGz8+g+itpCFxp8sohk/UlSc6
JAPGnW2mRQx1ubeXapQIHWFnvOjTXfsZrLBH3wvp3AysRbZG8nexAE7io5ZGsKriOw+OtAgO7Uq0
zOKxmuI3CetDEHWBGaKqcR5EMxfvNvYzSOPt/niVVtpv0Yu+UkvvVmaQM4tntVWyINZFhlqeqavV
l6EIdbfpJbujH4CHD4Zu81UpsWItz+aMtQTj7sjt4IShrdc6DbRTDo7YBmj8s6GyYhVb+m+9LInU
8HuAMz2fbHSHKVH0ztImEPKVaGBexG47iSpqKxHKn+XQM1l+JU8E+G2kVPtYckq+jrbv3ZPLSXk2
rXsFjxbDmf0hrbJ0VEsYLn+V5YT5kHby3jr00LakvEB1k3jjyOCHJKZgoVKOPvq/MF9Bm5LJcmOM
C2W4rsiXwkOLqs5WjQKVQv4VVlXYGnnWnyjpf8HWRG+gt111QV2Xi5eMoxCk1tgwczYN0RVWd2m7
THAI5kEJ0tL6xJdYI4k0UlsBaRMq2rjeaaP10blAXJSkfZ1zcjqbpDtdZXWy+DhbCV0KUuVR6Uh2
S+xQh7NUDGXz6a6TOT9cKuNgmnXDe1pDFc5qLnen8nNpUfEoDuUcgTggKNkROeruuihhgz5Tesr+
YNkpUoLJkD2L5YT3XgRKQGg1RjzceFvZb0c6eIh/FdRvNbS+zwt1bz13naqKPHl1j5ACVlwC5W/0
sCZJmCNCmJvsAOXdBJJcd/57y5deq9MH0bZ2TLNgGKzgOtWcITxUqmnT04IQDMWA6U3pSu4ehVTm
ObuksjMdmzQzdi6XARItmX5adLXXgugUOSfZ+0xv18M3sUMm4ezuigipjZBUD05bammiTGlJr/9K
GXldKH/1bft/AWdvtUmevFWvW8r6pzgABPxKKtV/NQBNa7OMjkMEdPgNWYxbScF5Y9dNl0MB51m4
CWHQRkt4L0kHr4C3gc2R7MeKsv9JxGMXCtTeHi4/5k8ObSx6dE/ciaqLHwx19dBTN2H+Ml1KTG3z
ewYTBdfYU05CcqqzW0sUZaNKklDV2gcDmFhDVz9HHO9LZTnXy5U8HBYxo4v8PjKQCqj6N6+jFLdG
ZetvGs8+4boaMqtwXFOhHk+DBVGOHkALZzAGYETuBGuyO8ec6gcuVah0C5utEPAEuBvVfEaAWcla
ZVd4HexM/UzTK1KRWGXXZr2BiDgSbaYWLNuZ+IhfqBTXEeamj9f9Y9z6G6xT2HrVmZ7rgMiB1zGI
ieZ1BWmI6kvVPZEjXkwPzFmhFMrS9xvcpCi8iRtxj4hLps71aq+xB/+fcLJFpfn7+Vs02OR7/RS+
69RkLmPux32u+LVfvJpO3Qn+lSrNSTfaq4NDiSl1WcPdAYZcQTrVk2zxSzeyYOBUSLd24IQ4i38T
32wH/vQxEu2Y4zXmst1ht58UG3aKYnNbNqMi35bFCsgV8ViSuOLPRKBq0wf1NE8166+9VpDM2Ftc
1yadiHnTQ/Z1ncMMU4SiIN7qm2Fh+tVkCIuZf1NXqcjAFLyzE84n2JKWT6G+xvaMjKddRqCNjqwh
lMP1z7JdiVjdiOudka7+X0IYEVT0gOIiYG7xiWaMrsEuKSrXo/GYUTacHY/gSUgCUAkQrBx+GfGv
IFAuCeqr+KF8WZiZMxDr4YjeHMw4yUyME6hr7mGgpt1GIqA4/yPySJGZ+fqJqYQMhqY+WSJSWvID
vqaJrTz7JE/UoxqCwrIsqAPRyvH4t8dpwPIaTsJ1Lzm9wqBUMfoRFW73eoGwa8GlSaGNM4CYcEiy
G3aU+wHExrMopHev9cZnYtOtD55HPBDsmqMlbGWwKBrLNHMmNWTSHR3RkLJwL9FU+uaczsY+0Sk9
agR+RJsb/kjRD/+hMtGjAIXrY8PlzfkhrANj+6QE6vT4pgM/GJ1Vw4blIrC4+aZQOrGqZsPDD4gS
T40L3Y7Hl2DUP883COZIMlihSYpVeKc36XeJX5FbkeER8WQkBJ5F4uNK2WPUGVAuS8mge8xEWK11
vO5N+fDa1Bo2BrtyCEKiloVyHcAgOWYsXep+JrorI7efMU2oBOHehRy3QXJSsgyWpMWvN7Kgujyh
11AZ64DtfbxPrAWYkXbVc16pFNw7wD2YOWOb+neR9qHoTinQ9EvRlX28J8Hl4xI/fTyLSIl/34mi
RHVfcdMnlWmspytYrgOHCHbw+iulfGo/GKS4560yzX/i3FYXN1RLbU2M08W2rvCcy62iw3wNfaCx
weWbB6WNgcMvqIx053qY2ldX71v795NaVlS6p2/2rao/PjPgE0xGG/HU0WUoYYPhngV3e9+1Zfb7
bOdBr4xIT/MaT+7OfOUNAVj3DG6G2KMN6I/mlLtF1oSnY+8Bge6HmqKP0nqfvPDfG7X+TE8jgfkV
3IiI+YH/XBjLiaf17U8sAhqTGBsm/1hhnWFeKqHe0ExIlvwL6DgfNahvXTn79X5wcC2mZlu9yhfD
0RVDpP3zgz1B1o2WzorZld/qoR9HZ+7K4BsCvNc7RttE9lXD3iokEoQr3sKY2QV8t1HOE4cp3sdf
G1mIlTuyRtHo9A2I1TsN1r1qGh4e4KoFLeJLQnslJlS/neSm7GezYYephs9VTVpzmwvDuqLPqLTn
1H0CGbmeZjnCJEJKJOYSu3bHsGi4I+lYM836l3IL0wyuJhfVwirRedOK1COGNVivP64YUId+fcBm
6Py7VT6HBfwMtrKQTidBAlm05kHo1wdLt40U2GCLKLyKDAxGAds/S/4ltWWlG+EoEIrszPKSkzxl
2c5OT1JmJaN6OCK2TKUSWL47K86BJJtx4OgscZAqx3aMgAPie8kuJm+U++jUGa+iqeyj9YBA3tCR
Cx5CJkt1sRwVTdvYI5O4ChiwS1kJAuEbtT9++WJ/AYe5ZCx8CR0HCpxyZANRyEO4fEVAOoMzyd7B
XXNNummOser+QWpR1stds5BS4aegxZcV7uXj7Ff/R9Dqlm7+VIrap98YYfMKCaKFBiAQAiRNxN6O
G9zgvxeKC9KZpE2v5t59oZXm6pgl9cjBgrWmC7qDzYSake0uute5PunymTf5bKR0QzUkU3tUDqZe
IMtZDhZA7TCuRC6CbGWECe01fpuLzuDrw/W0OJF8kI9FBdUPuTRPzRPD43oElMTH4fZfb71/u9pr
xm93B2IPXTNyRH5O7bcECUKeU6V37ghOF4OcbHhLXaK7F0ii6xqsNBqoduVfNmQYkGJjz41v0rlk
IvW/9C3GDAH7uyDxJyC5mhKW/4/USN80m7Cc8FuhZeH+htDQ6xFIBxXsDrjg6Jnd63qNR+FKLD25
s4yVOxtJhgc0mycUp36DMS21/mWWY1sxvqgHaAS2CNlbsCxTT0isvfHCJsgH1R2WQyMIGjHQNebl
ErRifshKS/uByDvKZfZWepSy47MhUWbvyG3qfshfMM8WJG6Pv0Du8QKeLizbg7Ew+9QYErUMrlyB
CRR/jh3vc1oHS9FmoUg4fG87CC+ilxCS71lIk8D6y/ntgxD3e1JDyka/R0Kju22d1mkl31iZ0oKT
O0r8Zefkxx158+0BgcPE2ajbWHV50qHybnY34UMA+p4swKux95ZhUG9J4ftceQUGMEMrmL22G5bG
AM3c5giTlxWdDOReD4Pw/LbeUoXKxU1FbKk9J12FvGw8vlo6nNUa68EESbT3Gy3ZU9NOMorb/v6n
WjjrfPTsHMKq/wGpf38o88LHYEMcGoWBA8/MFc7g3pCmLyqxVsLQy2cVowt6xWvd9g+sCPpVfYG4
vSIt1xytUVhLxS5Ip6lFSv/XZBcz8iLLvpniSKrf3GAz7wM9dWVsJ9CD3LN3sB27QfEbhH2icJ6E
6vgeFDaJ7mETWWkjBhtk9KyOissJRz5+MiWJoHnV1OllFAKjaP2iS/bD7XQQ6/E5mLyA6Vz5WfKj
NaFJNGf4jasPWGxdL5BWqu+5XirEBzkQqNwK3B3iUS70Rd4URKTgfGdzwlGDN8wLsidtaL4uiJB7
xokl3IHzXQpiR+7cD2IOMVxIQ+YoncNHBH6H0baV4pQ+EowVESzBJao442DWnidZub/vKQMcUHWo
djXsAbcY91itaKWvPIr2w00U+vvQn7Rf9XIVj1og6x42BQse/gvPR2pz9ABwQsDkgCF0TmAtlqQq
QReyIeapdOiWONantNkO9+kGEKYxvUYQO3LpyaoQePitdt7qsseiTA0J2JS1d+ORePt9Ln+qjy4n
mDcjJVz7ZnW41DP280E+iOVggETXPjX5KH/GgI7X4KJF9DE7jkSuxohGDdVI4MDUJ7Zi0MAHAqAX
KQCOd6nzt1SPtXsQwLry8OodM0M/M1YLS4T0E5oDfT53Q0h/GVt3/l0Olhjy/DKcntWDdML2dZCJ
H6rPk+pRaGtRs6L2pNhz2xv5TskI5p6KBWddU6v5/EnnE5DjxIeSKm3NjLhKCuzQnxSMFIUbAw5D
vUWWc4JtUpYwPfYJF8Xu5oobTvp6QJyNQLjGSAs2uVDDdJYA+55TkseI3YCveHwSv5kncg9fHSDG
Slw7Uax8IDXTUwD7swLTd4FWyKIByHOS8Pu+6+8a8fo1+0yIeAmS+VTRutPp5Jgz6PcNt55RbdHU
525A2C5BQRsPFp1kBShiISX6Xk/QobiqXQaNYL0o+cJWi0qayx1BhpcPLM90gZFRyywsNfbziXwW
eRgIiGo/ckw2MfjPgvXmqxG72Kr+5vTVl7s02tfIt+QgBHJ6zcFt69nADSNFwPAUcalwuDQ0iIIt
4a8Cuhfmv1lkrMNe4UVeTXIG8Fwk0Z4fwEmq5M2V8xP+jfnR5LK+L2eKhmGtAZY0PgbyfNnAVkFS
m7m+xsMCs/+AQKUdkF7dfKedoMyG3rOfEqC3AyJdYb7LMQnP2z6H/tXSKidOvGsjOl/2nWw85dZc
dJKRnAYVhA0AhSbTLd9xCEq5wzWX7mdspTTdipAt/z+Vz7jiOCs8KlBLg23zbngQQPFOJXVu9gQA
o+LlQXaQGx/wpt13IEOGyari7TZl18qk0zMfBMWIkvHJfjMI1okHrddUuYhXy/T/vHcyj9v+e8z/
HHjjte7B5NP0CpmQ3cn6AkXIidYX92bYZVItZcc93Re107wQ6+H03jefIm+ETwLXG4S248Jlw1Xz
AN8+AIAFPh3GKHaUNWWmObuaV9uc47TNnN+8bmNnShtEz0vHDOldZIPQlhTHlrUSCOzU3iXeye2F
x4/86AY1YAqIArhF/2fgetUeQMpTWY7M6P9RcWpnP483msxsrD4CZFKz7yFjzYH+TM4cmk0YwNw8
sVXIHzBIpboxBCYX0Td7B+4FykHBTDAcDjlA6YHvKKKWakRkArc0eIToVbw7eRy/1AecquUoVf+b
u/WfN8KLBDadeZtm8I3/TDbUMPdMkjjBTrN4Dlq6Zf9XbrAw6tiXNheUYmanwD1uvKaysFkx4iEX
HOWv1at6DebynOPOXvUXGS3zzcv5QI0G6hV9p4efN5c1ka+34lSWp2tRVKPeHUVoVrjt9nLGbasj
kLChzJOBKQNHKcqH+t19ogCjmjXgrCLJc/VXsYWRCsbHfT4vZSgcJB7IovYW9Zfffvng+rj8Kn24
w/IPZn0lVGcFKh95E8f1ha1PiQVwKSCeQ6OUIGCfPOP8Lc4n9KuIeJBsO1urHedXtaRdWzmFY+cX
brKbdOxgmSMNNl3J161O0i+nKWc5GNZB0G7AURJ4o1mm01QSHX1ZkWXeEQqF6RU2nRrwjm0Aznv/
kqDBozQuqinw77/DIowV/AU8M45sFKKT1PTWEtpx9c77ljCEaJMpzaoYx3vz9+FldTNujapmzRVg
SjMZmQ96zgRpu7L+eEs1P3GLXqLyQIXpKTfjYRnPFYntPLxmoy0nJ+TopkqAWzlC4Ug79qH+YtX/
PMx1UCq6kl3diLwxYOHMOhcKHG8GYbAqS4vkUrS4c57CEXGMirrmOPSVSszY2szaYHQg1bT5nj9k
W7PzGL2br9QYR4Yc3nOLKMHTqdAe0Z5o2L3GfYoZsV8lb2VsSvfDQbU30g5Yrp/qBYwdV2vexqP5
jt8koZTCywSF57MI5QhJgDw8S6x/9LUj0gPsw2pSlR5Vvrn+GFvx87FfanjAsxN8dEsCZFjDd/tS
8PBGEQahRoy+7iweJQLMguO5phSDoplGLSSJLvhLlkA/XAXw9xxkhAO3KoyvL2ErNv2BCUjAEgBQ
bLrj61TFuGrbiVCuANIUCOLKuglr73m4UTqxFYuP2AAjkunB1LxlgKWWxNpxa6WL2tEbBZ11Zalh
+zb9xU+RmnyswteSApOX7BfZ6FxDv7ZhYvnogXj4KnYEhmPAHqGX4v1u8ZFz0de8LTgvkHssPgT1
/llWwkXkYybcpD4pN567ELYhJBAyJL0WvdWnTH5okE0NKDew+AdjxPuMwGXxBAHpJz1ZW4h7N46H
XuOO+gr+M85DXzyMMElGKHPinOPimY7q27HM0Go160CNv++iLDp85w/aGMCOnivxg9ljS3SmMTem
CjTncdWkvuIYzuSCO3MAzLkcADib10RiW/WsO60i6Pbg1P+jy/DivEKkb8faAUypnM+rcPKn90M3
iiXbH5N5Xu64+xmF/HR8y8BSLOn/0UkD6vkfyRuRedniaW0UvSAX09fyVQlyP5jqxCz+gOSCm9kr
jzb6EFf0SpfutwyNSSlengIISFQ53DcDjT1y86GEr98zSqYc0AcDHdmjvipR/5Lso6R315dR/2se
VWTEaHPl0qWLE66kXV+CajqtQpykyxTIZdz0HBYg9oeFt/gSTySDoerKbTlUb55726GkcQ1r0hC+
deGS1s/Wa51/sfx5rTzEjJbv+ccVKCzqE12GDwwgD8KfkKFupW7/FavpL7I+Lzcwl4KjEh70GW6A
UNj0cnZ38w2o/NxlE4gJza1IucIYFjVWqgKDeH8LI0GbLZeGdgEa3nYK+BAi2f3sLJzpTCMEB+7g
pklkWxuu2Q/7MJbOWfq9jhvNpzxuzfFskj6XInwHwen1ENHdTQe3OKSaUZB0q7M5A/W+Z0D3uss0
L2cnBmZpivQrSWW2MCaFnNdQ5y7VizutFN1z0XY3shLbf0NP5b3qAfElRdzOKrdOE2AMNTDLOKfd
YZAbJZHAf3JGZkj5BlCSpPz8iHxD0+OBjhrmSyeJ7oLrzWq6IGyOyZSRii9V4L65mRK/8ATkziTx
dIWzXXGwdchu1ooB3amrIAMVJB2EmT6RLdZrwWZ2TeOg3T74ecZS6Y9TTe0fAd7jXYXFV7icJaMS
eqm5u/mMO7d5+Pl2F8sxZUG5NspM1ES26AL47NYpAsSO41L49MnjYSsdXKzx54+u7qhVZk3Qto3b
ssXhvlEcE16CJi3zdTZRnAbMTW/nQj96GDzqiWn7/5jdFI6eD7A5+obaARg3z9AK6TQsBtElMS3x
CCK02iRTQZzsbDGlzEQOMC8mkBT6rIxLwmoE33nrBPMst8ejpkerKFufS1Bo8CVjvNCY9TrWzLux
qaVw6+2AkBPjSeyZDhvJkJaZoie5jejt3P8tQIdnzKgOo9MlaRAuI1QcdH9fiP+SSTMIze3v7Bk8
XV9hWGcKfzQX1JJFQfnC7nXZ1P+h9pxCNeOpKdkZOrekW0wbHCOLw9diR3+l9ILg0IOlEIEr6zKU
8KCb8oVou/agsbxe+OyKQitYPoLqljGSk0DRKDQTsy1W3jbwPMOeKptBKSoEtPwzkW5QT+CnnsAF
YwVMKGfdCu57VXir3QYpuK5kUJ8D65/jdgfAdujbQsG2ko1gPQk27wc6e80D8gOBuXIHPqhCeSbv
t9F/NHGMbFa242IZTHANn7T+vtlFMATMdv6El0MLnVdIa4gWdBMpgEY6NVuLclPBN5Ww9yjk1b47
qOLbv1xVu2EXp8S9VdgrAD4WmnQh0hQ8UFATkfj7XQi3UFSy/RpYtNHudHewV1AnfhfHPAE8JGwn
wCcR6FX+7q1wBac4uZzZt2/jtkqOmV4LSGupa7YuCrSAMwsmsZf7lDTPPPpqw33LBQomh0l7naIb
U7wyZgjSzf+c2y72LCdW2HLT3YgZhZCAG06g9i9MoUIj9SYg1FFlcTmgHORxLexw8B1RqR4PSjev
4EvF6Y3664/u0CAZeUWIxXYghXc9YZjAohgca3JfXGmkYdourjZDFtmJZmOA1lstxi4Jq0tOd2QA
Z1IR1Q1PcNZtbjJ9TZqH5vxFIxHDRowS5FWysmximPgwYvJOq0mc72OAggVs25Ay+QniM/YTFRm7
ELn+f439Ftb1KpSqpL+gkoQYgC5I2xNrUsXXNgj5T+DVykdO4PPZHOqLG04Fn1Cmm+IC7tk2/k+w
6K7B3qyHhL7iOKj3WW5fCxTvEwIVJQbtjfr8RF45x1NIqLvMxXPclxAgFRN1BsIIMe6lvftEM2Gy
UNly/ezbZf7YfiwmPBZx/AItRYPT/T86LPJhj+ZJZCSkpZPaxoa576Owi3C+r+r4RLNYr1GhLZda
jMxFw1WZe6AigoqWeQ8h79CwYp6MHIgknaf1NbKHjr40fYq7gpBEcxRhMCHZN2jfNJKjWhPu++hm
6+PvMHkjb5AAq8AgbxyeoQmylE549ob/wGwAks9RIxCt1iXXFKRLwLgUnXGEK5ei2cxrzXx02hkD
g7nbg3buYmWLoo9B+RAk7oH5WAMFzzbDIJSCwjD9DKzFdlJ4Z8dhxp5UAeFyI72tTGC7nf9kAlIv
HfcAFXfnr7UMwA7HXEI7jUnNBsaeuRmNiqDFIDqJsbcsWSwjcisNON41AznYUR6LfXDm41Awwp6I
vluQmmz3eYZTuwEzZjVGULqBRB14hvre+WQgHEBdcvi3SV1y7K2EWZnEUpz0TtJwhx6qMANgyOMz
BuefwgQ3ggfEL4C1ZYGIp2HP8w1WtmPPTMY8vYNv9qmi1vkfcsaTyFHHsJidsCFRA8A36HL0xO8P
6ubSFkwco5+dCtiJsN6Jg+5e22N0ABgVkJcJbQG70iSlBffRVSlOWOIP6DtPgbhIlVY7u2L78iZ3
RoiibblcFdffi7ionXHrOxK5x2WUE0Xd1gYVv1pzl8jkOU581AhNKAPFgx54rrjcjsEvydLH9/OR
vVeU3i9br4FQ7RlFcq7Dd4qopnybg+b8oII2Z6y9dziy98f+7qaCW8nG74ryiEy+3DFTS6LHnguK
mxhud/LDciSKvfYIO25k6wdPuLs6CbQHOyef/godL2qcWfDz6pYBQRaBXxZU27eQVcX8WwG+4HDk
7kZxLTXfTQQ9ZJqImRv9oLpQO8MjCTrv0JUW6S3vl4YtqWZbHSj7NcJVyPraN6t9u5lv4as8bm8P
gLkW8K/6NWQ18S1OOL1xhMMlxGeolYkzD8VbXISo2VTnjln00tqvbPC6bfV5puUf+Yq3V2i1JkNi
GhbqKdGmqMBoMmlCWHWzA0+wKTvyNgn0I/A7UJaRE3Rh+ScB9p4vpS7xEPRF8bfOotnULa4is7qG
VNTSDlrfQnqDuFwGyOjMnNi/nEqmzRnTvHq7crF88DmB8oLLSicd5H5uccEKj+cBT3xFVaRpoX1b
VCDDjeoNAKxEXyMglWGkErixzpcmB5G5Piv7p+RZgTAZT6GOXQNNQ8UG6Vu1OtNkcerEhwLL3yrr
t7cafEu+RdwHQUWe+lxTWCWM1BPBZCVrDNoMpuziGh/XcRIxRjaByj2L8eHoaM2kz8k4emEkeImh
iCYPvwPVqyRBdasnLTTT8T3R6Fz4y0TLoeNaLKuXEaTcLKeWPDMqOqfS7tQ602wdWGTenjRsL08l
BB/tiv7z6bOzZlJC5dJ55Ve7YaJ3LBeQOeuqUIK8PYLUU/DY37IgOAZN653J8o1ptGBuldBppmHP
FCwoglmNaBJ4MQCssr5BQ4JVhvb0Qoq4PKtF68TzDRTQe3IRMNWaJuYmyxtKje+n/6b/+G7nAFWB
mtQnnNL2hsI3UaIo6mkyy/I04FgTNRpH4WXPsJVnxFpavc4LQ3U4p66BL0yQp3/4bCn31Nu4SA99
s59GDSgkObDOZIpG7f/yZP3BFQw1QppGuK3o+tQFPijATtr/FihIB+QZIgJuteM2iX9az8m9m4LT
O4uMERCJjanwLPeufIjkxSyrblFkN3UhAumS/3j3Ul46+0nqra6aV76hPKGKRJ4G2Y4NlbTgCYir
LytlmeFZhW3L1H4KHR8HL9fFEJF0yEZkZycWz+alJELT3JA1ZW+VkGW94fnxNrm8MKKr01qu0HkC
sH7exCvc1lK30mv2p+eW0bN/PX7eIzxfA3i/GbZVY4uIxrFsC0AhNcYdMQ7gaNZLSyHYOlyRf0Ky
wUCRxH1kzX2uBxY15WCn+mZBQ/ReN6UP3RnGaF/DPzSMNSwKfUgZF1EC3xyxlwMeIqndRo89LYSa
KcGHC0QYnZkhp3W8BCPH+Hy8r9ksuTVooj9yaavixagCDS1c70AWkuR7UL0aSGwSPy65InCGbGDQ
cUX8+Q2ykd2V1g5sCn4ox9dap8PyzzTjUvpdS3v6FentGL1nypwXtw+Bn9L/ZKdgy4Z3TLIDSty2
YUk2zHGAn+/rDeBDVA5Byyr8QFww9P1cOOYYg28FyS1E92Aa0DIKzqVWKH6G+zaOFMryB1T8IvcW
NZOetjlr42AqFVQxRkS8X7kbNsfTJbS7eKQGCEIlmb1xALTKkBC1tD/GWLEkyBTvk6YAtpVJVgTq
b1akswSCObM0tBzan935nj6uyd/fqoYIay6P7l1z5rC9pgCpPR2eBD/oRtPR2Upok/6U5zSZYn/V
vxFOmrgaloeZ15B80yzpDw9i7/89YNlnih+gy/a0Zvykas3NMRlu3w1esp5YxBwxy4gZnEfdIx+2
5fBfCD7FM5qZnOB8djqxI/AGYcx1mF+ibXSS1j8/FfNLfVMtGk70o220ZmmdMZDa9QIgGDZwRch7
XFgq5uFNS6vhGQTrn5kJV9OhHO28TJGIG/ya7zL9iTE6WVe/UoIL7XGYp+moTdgRQ0YR5b9VFINb
8FJaCMzBjK3/kN+T/Xz7N76dYc9e1LXHHspgUu11lWYZ+UXnnwOYBsX6wH5SdNK7gEc35XYS+0FH
JQJwG4oHA/c17VseyuxETqxsUjvqRUIIb+Y1/IYMiANtOPlZQhprF0F5QF7un6rgLIUKwmPx9yPC
Nvg97wEgxnM7DEr0OkbTMfIZtD9d18SZ3NRsZXpOG1pPCiLVPeKTm6uFHYtdN3AW72IXoYXHzSXh
dFNFqBsuPke1KGE5h1bxFNCM2cqvqP005AcLVidXWSSY5tJWJRnNpOAJr/w24QlBEGbeoBOt1bFN
kHVl11abUyJJrwo7p4i65yWrwfj/EQiIkpr59XSxIHb+Pb6ymMESqknwGWIMQt9xfhkbUMQhGZKJ
Lc8mGj06ycEdcYCdYpxVCxs71Z+hnXSHkE/5T3JW5kA1PWBn3a+4+XHQ/sUq8mlQicF936MmIl+k
QBll+pNUfgytB0N2QAItqqre4Eu/G3PBc/btOuEeDS+iB4JSAwppgEbPRIQkWWU2vsKH1VQq7pDo
O5Voi2EFO3PdMdJPmPx55LZWNoFlmRvpc1rgsmUNUCKiAnlG8434+QyNAGAE/+8AYq2W+9xdtCz5
zzWsB7jbWUP1AdvduIHrgBhYnsG0n5AAdwxOoCvNK5QuxOHyJS4X2Wxj1d1nan9yLXDbs90wf4OQ
jXXwbYivsio3DnEl0tww5AqLv4t3+bDXCXeue85ns7xJmNd5JNppjIcHUvA4jw0A7PY1/TLm+ARE
RPSf4ZV/kvpnMCFk4r6wqab39s4W/O4WwS9uT7hNy7IE0hMeAXzGh0liy7kdK3UB1GKZ7MGvvR4G
ykBT0gp9rEFEjlTecG2D/cQURypp+QSipIHwGT3nFMZ21xTrmqvZwm3N9s3lGgw8fCybevmeylhW
EJSsmnHoeziyfS81KqeKI2fdnziTtDK6Int/CAd3nYKkTpNs583lH/upbn0me2HGA6ZlAqdg/THx
PEjBPezDJh/H/dj0u1/vJAGgZ8TtQXgHoXrWDSZWLAW0EZckQajJtripBYaQGBbmLx1j2NI6ve7P
tWK+LO/UyyAE1w1RIO2A//2x2sPkIYvO2N1/gP51HkDXCIIcQcPe2fJn3u73/Hur1HdMleonEVOG
rE0AaQPqrjRuihGdIiy3lEZjsyXWpTzOoWdP4S+x960mmSbRkwPd6iNPP9YY0r5LoQtKC/5kzioL
Ur/bn88VHueoiX5oA4hhXeiPQv5451AhP1OhnvDSd7rxs7PKGQUA3U3bT/+QOB4XrO/DrDux2CD8
dX6p/7ItI2Ip/pHf1soc7gcOONLh7UPoECVmfzY3awQl/ZL0yI1ZVENVyHoNrs+pc1mvfH1zPGHu
4Ke+OMBNL65F4RdaQ4ZVzf+mYxgcYUChJ1Zx2mwj08X9zy669ip7XWF35WuT+pbPyoGDtaMLxb5S
Y66I2ZxYeFbwWOPNKz7Vlv7c+9Z9R0AdirDNtre9TzfXGkTVSga2UGAnjj02Q+ARQLBTpIjkQ/ah
WBslyh6AxT26px0hd+9d6Z9eBZ4M+UJl02yIFJaATxYzycECEvP0391F9apCGdh1QJNIMcOGYKac
1c34c9zzcdG2gdgfx5XZSSVWTBTlBR8peUZoTshNGLLeYLHQE0D8NXTF38ki/4CMS9AMjcRUkyzT
25gViZwghTFLgZY7gxyoU4Jh2jkiqwD5kWIKRA5SWJ3I1vF97A2z2NK/vT8ULuTMhctPuRUxHTAa
AwsVfv6pRiT5d4qIPpvnYnDAGGME/mGCzP5u5NlTbT6aK0pQ7PH55gHbYAaQVV14Q6QCYMtZorPj
xAYWBYc8cGr6+BdSmUa/S/ztMQSLt32EtHpICAybTCUUtr+lpzcjkIjyiwbd4Z+Vx9xg9ZXDQ4iU
GYyTr04r6Mj59jbLMXRiK7VW81sZQLg/X6fV/wWlgPzvrlnell0Ccc4YMDhEXDQmD3YwQwD3w9Gt
z4O9rpNLWByKGLWNbf3otrE7qKIPsr6fZnlGyx7qOJCsA8cyieiB54TTyzvxfSr5yKlI47yYJE+R
W/cr4QaMJFy/NW18h6gVS/EFoP/q+YN8pJHXNzVbZs/wlPpvDBWFQPA3trZjWVkTMzoa0UNH70Ob
9sno0+GdfGC/Ua5Kxk50ORKmHYA94YksoDv+qEZm+ruj6AWqdGJxK40Rv/1W2NN5pj/KVLQLaQcs
sSbsShlmkHldsUr4KFSIGI1uaPCr7qc7SvU813IK6wCPcNbmXU4MDxWrAkvWIyhd6wnMevR0wEXU
6RkeR/D0jLrJtSXDpwmp/h5nM0ik1M5Qiwfd1LkjlHpmh4uIAZuJSBAo3V7BPYMTTnPizfJBRAit
GaPfyEplLzb8xoqvz78GDdO0DqnedBC/9UuFijCO36qcL4UzX/33rPw2QbAWfNQhHcpDj8BMMLR3
v+dsHjRGjZhq6GjhzpYtbM4TrRi25nmOZGwzvCytlHkryG33f+NO03u8AxCC1UE9Ny3FRExJ+OFM
lhb7c/XJjb8JDlg3dwZTjKcOu1sjae9moym2SjSWC9wnOcF1lDiy9EKzz9FSw7UY8A1+5WLoplNg
Lsug4HrS0yUJ3hIthJ0f8rCwLuRP/TFemKktFlwYwq8IYs5WcYMdA6iXvqTWtgv876CeZPr9UArP
JwPKmeXgDxGR122VbH4yOCdqSYe+dCXRsX/vMDUWtVhE/VxQvsGZd8ThlW0dzxriYYzChDXLjCKA
p4HIxyeU96lkGcsDitYPb/rzU9lGOhGo52mmDYbrq5iEAtaaVwWiuDlel+s+X+/GkqK6pG0EQR6u
Fq4rLW+E+eU7uBatlNmWlRFmFDGdVnYa0/W+bL4q/6bPF58CY+3fFafAP5bV9NP4OVw9kKn55zmJ
H/nyesnsrUGqJphcgeARcZhuDepkotWj8dNZhMhjMmc9N/p38/2+N3q+vdxyhYBIoSQKp1liycxS
UBSQ4LrMZWvG2pA+nXR2g+ZYaDd9CYbXudaepgT6jhmWj0ejnoVHsMOW87uhnfwrqnieUxTbwuEW
/PSLtGy7tedzudY1iKfODhzYDyKhyZBb1LAJbE1GsXo+uadIhLM+q8DsOYcMdPfDfF+Cv8dKilyQ
zKNuOdDl4t1hrWNwdlwJa3ToWIJA6fc8yA8+xeUU5MNrtYw8PWCdXxJsbAYdZI1v6jcLG4Vu4g2k
gRveW5xIvAN+iJuzo0XUjoSMUUJtW9K+V0VZMUGvSbEJZk944pbVOCWoiJvmfd2bdXxCx+Mbf54Z
lfnEF4gy0Vw8uAb1tn7X20/AWSHyLAkkK/8ASDS2u/Ca1VLdRcochgieY6BxAiPErPoiUjrZY7r8
m4ubj2mtatGSdkLiqIFA11uxoItU6hIVcsyZjclbI9h7n5tq4RDelzWDpur7ts+DialzMkO1GiX2
A9qRuJAeESipMqA+HhLVHNc2XrNa/CCYAzHsEgHXb6NZEi2CPgrud4BcgITCrIzihxofbpQ7aQDO
ybttmmOth3vt4LbEftS+me0JRM0JOSc2I3w9nrZ+dI1YP1wOkKFRrDXG1qHZuY/nd4Jm58O1jH7F
GeZTArfpxnYviQxardVbDWMAz4F79bCS8cfWbGpSLfYnuWwPUhDNAwLl+2SJYSKkvhDxo2p8jRU4
2bWZIz7lefYBVdHqQfH//OD7t3DyKIoUiVYjr1VTmd53rH2YBNe+VGSQf4tW91Aom8pEmrWRcN9S
91QZYzm5pMTRdhCrhH9eIrd2otTyf6nJeIkGa1CNbJnvLL18HhT6nj+fzwARCl3BFUZvAoLl9WIv
4/2pCw2byQidbVRYbTFhQ17ZDdx4cRqwSAaGboxG0LCoWguAXY+KfX39LxhFaYTMapJ3qSrZjYtS
BCMsFc6Zxoc8hzjqy26mIgO7s8icYeigbNxLENauEKXHNI89vRxM5q2sQ20kZTVFmzvNu9SyQ0GK
fAFio+E8MMc/WgyPrNBqHa3+c7ZzLMF50zFGl9ruSrZyn2wQ5k2acL+wElRt0zOncGuVTBnYRo/W
JrX1nCXFy3iAuveLICsOru9v/xwbq2Oj9l+En9WxgZZ3419BPkKcJDYhDhBg0ogk5ItvTA7M5pxu
3Z+tnz26CoXn8wVDyTRrTBmu9nvULF4znlnG2QyQIUcpAeqDTtrdFz0IMmpzzP68qL32sFo92VS0
bxUKUqtcrJ+Ut1Hw4Hb3IwCY52ncay4u6RNwVIWkbXpTQzpGrH9pPy2+t9pW73sEC0fLgiF5jdmq
cwI0qGR21LYAXOevvmMQ9zw34XjTyr4IOKy8p3u7UdNO+ntYggJMmyxAXyeZmP2Uzd8DZqD9dR+H
p8f0uWFXUlBvrriFxblvExLCA48HduYQ01PILBwNiPFixSMIMwpXijV23rLRU/l8Vl6tkcwi0vJc
DOKWeJUiUPtfLAF0SDR6Wg1WLeP1iaKKQf0hntBVptZ1EycvF7quEGuYbu6oiAqIPzT8do2MmvAx
V45T/2s1BwAICclxs9cY7XV5LD5NZ0eiZvDJo4bys+774HU4dq7TM1ZJ6qqWfGBhUyljEdVYm6Op
1e4KUP93WmaUsEuj1rHJyCAuJFTwWwINkgRf31PTBQI/Bj2HDU5fy+F7VS/r5FsW9mEh7utMFd5s
TrPv+rcIjCfmZyzKe5EroLT21oQegbmYlVV0TAsyIchVjcMTGKCcfUokuo+ns0FWhlOraWb7uNDo
Ftg9dyNfnAhDYZjh50zO6JCN3iXNZe0DxX1gZtbAB16YJAnEH3mnDt93Yiik+FKTBqOO6ud1pElS
T3cStFziO5qfBG7H/f4oZzQMRjkGVhj+kuaL9PBjoDXNSA7R4F4rGtYI9/DDsceBSll5ccgReNLY
4/UGLp6aoMSpY+iX+BLZmAngTiLV5l2pB71XH5rK0sjeEgw9JJeCn2b1caemPDiteFQ3TXlhynIA
Hb6VA2h3Gkw0X7fO92VNufX/tHyJnEkpdEU3FMcZl5wBMccjD/wPWumyAtsG/mHqv/hsVmwVKLHf
grGYF6bmNfoQFzgX9tKnDOSKStXI9EpdPCI60hM+J6UtGjxQV/zDqxFn6oSa3sZfNlpra7FTMS+d
OzpTm8nvhOEopUnR+KX+P5EnES4SVj4h5rzA0N/3GA3eAzf7MIHiDauKmbuQ1uRfctP0Gt0mysXQ
XRQeWI1OD4Mr7cEy/zaajWlGFvF8AK3EEESUZvBAib/lWyFtdv4XOsJcJUJqG+11U1Ep6GGn3WJU
CVF0dSKFDBchCyFODed0A3jAWGg6i5ZRrLlVPFfT1zHT+mZ/oRBunLhG85SxjlKQCx05nO3pdkAk
6pbUlB7GVLwWDdxEIw0d46bU9wo5d2b3QODIyurxOmTpBH1G/mUC/uXuYCpn3XnsNejibmXfa7RU
rgRmCqL1w3wDsW716HCot4s+2qSBX8mfL0yr/bcFcktXGCYyAi1+bwQAfvnpQd2F79sChoYQlmW1
T/GumjzBsRR6MPx0avIwYLao7Iys1tpwNvy4VMWXYdb9kI/t47hHXDIbAAa53DMKHlWRy1oAmfTT
LdHbDU4egQlwG1Jt/GlcWy8H0OxqTtssHVKFNCPn88wpCUz7McegeNNJ4KBUNscz0bhmoeUe3K0j
N+7Bi2bTPflwsEgB7TQiDSB9DA4FuVzLRdCczPKK5mntuQX/9wLk2a/sdaPzd3wo3Yw34TqWreZ1
I1duU4FUaUVxfanXOCJJpESXdMF86zuBsLGjAXinMPiVkvY9MKTxDsnjjiaeb0Ncns2trjlQhkEH
AR1bMDklnO0fEoijtMBVBsjq1/creorOBgdPpO20Jjm1cvQPNAzIumsUhqoMaLSOSO3tzTsQOuiJ
/mlLWQeCi9EvUlqJGXfZ9hb0NLdGEpVlCqonAm/Zs11rh7KkrdF/qKvHJFq12r8zdt5bLZ/Hnvf9
1Ql6Le8yBKrnKR2Gp32oaCB7PelVpfdOEUx7U73LaAOgB1DFZFIj8/AIqvb/DOcApNxBngGzZPYr
Zq+8JFRHSGujBqgGkqjOKWyzXe5IzeiE50dJH8odxlwudwPoAHW2rhyCtEQcRPflQELZoG9+wngw
dQF0zp7mZjOAsXHFsSQM6aASYNpTIZqDieMt76bpbOP4CorSBemJYV51a2I3cMmnwmrBtY/lo9+G
pwZ/6df4ZDbU6D8HvhHMRNGOKcgBKmLFgPQduMehrRzlpcyCgu/U092NRb6efYh7SIXS2QHSAG/1
3ck1RslOcDkUpgkQPBb7InEatqG1DJ2QVvi8pDqfQjMAlxXM1BS3DW9Gp9SU3ccYbES+8/itWFFC
d3vpHHKprB4Vvvc34pMufNYhDc6JQvAzo/3TrhYdPN9MmY+9N6MWZ4L/ljUaMWXge/FgSFnQQf0z
9EBrBeNeH4hAFVPDywPpqYvIjLFxtLdhaI9PNFzHTJwjoajtSUbrdfmdL+FK3u0yrUHEsVgjMcJs
odwRFruiEcTWTlRYt8OYWpgddLc6wMEed69a9e9uWei37NVkokZgAgX9+c2ml5jzvHHppfAMQasW
vwS++iwdN4R2h6GTfq3QA0I6BvoCOGX+H8hZmWHaf3U2i3LvxOAzT2odmVtpgS8BoRXP/kaS50UO
QX1P4i1kpjS15Y2NNgtxm9d2K4P51rUBP4/WFPK0gAVi5jdBLqli+f6kAUonPtYjYZQNZyqMTZE7
GBX1yueEaIKDRjMZQsz1KCuFApV28mhDXEK4YyMLuduhBJneoaDDdmVta3KmR1ByFH2W/TXKwP50
JzOvVUTbJSKgs5u7fo1C6rJCtO2Pri0Vdof6yrbsg6s5bTuGdHklokYPggytAkadX8yZ/RqHyrVk
fzM1cZwCi1QiGS5/XeXq7UfLULleNEDE6XN65cxOAtfvtLhsxnG9KwILELGxuWUG5PzN0RfFYdgc
uLwkqR0idhSw/thiGZLaVhJXNLBBrvlCxho412XO8GBTTl+G5tiJHpjpxihD8EGM94C2etMrlaS7
QkDfN3EBGM3XlscstN/3l7u5OSvBYrjNrbRE1gbP1ReskMN7pjDfwQyTGPHfWOzSZhx2KputX03i
TR780RJ47i9j2lshqW1M9Ssl2AG6vbru5ijaseLjL5ThVz0K5QV6gLsQiZ1XjMu3t5sAQcY78t1t
NgWLH6rr3iBmFzl+RD7zuC6EfZJdi+cmrFVZy2ZDXqF9iTGCzzv2iVE/BlvSCsK0eC78RnidjTA0
QD9F9FF7HmCgm5D+2/xytqTGvHfKO6dwBAVNSbjINrIiH3QhEXN+jLPGQKQJ+KXWK79dfvQ1tQPv
+4nIjtCGik+RsL1HaAtzKHHXpfHyjyo0Ip1OKf0x5m4vNHOXFhnKxpI116nSYYcay6uCq6PQPyPx
EvATRZ3iC/SyoPW7Au6gyQIZXkpy5CdCmuiPKJiT1uZSHNR47SzayfaWUkBecfGOOrVmlVYKNs5i
O0zfo5/j1GVLNQ9Wtb/2r9Uis5BIYdxQfqGAUOzGeDW3RIMJvfuTco5RPXESkQR9o4Pzu5ZJFCxm
LjQzcdJ7QKZ2CfTe/s5HtBibusmoj3Pu5Qq/yXitJvjr7gBzl40Tvw0Yjd3rDFOMddK09vegBQET
S5edIk8PmQ6FWDjuu82Y/DK7t7Uqk7VbBy/gsPWHCV0OtCy6QsORFd4RkTxKQQrJR2N83veeQeGr
DNgxXfHPGikm/y3wKha2zcNX0ofNZiOa6ducoY16SPChZhJ8oGLZRaZUBgZWclo8CP3kozEZ5L3+
C7USEGfFQH0X25TyLufZIG4CWTC73kKFYwA0Tfbzhe3zKwhv6nVMPTg7nHFKWi3CZuRUdZyxdogV
u/Bosy33U4BYtZDJAxXdbL331J1nNwgkzYgIF59i4tet1RpdXIasYu6/xVo748TLyBefSOTbEfhN
0tSlT+PMsb7Qmg2fh69y6wfyz1b4D0kkC1y3OCGtT1abRJ+gnthRfckSKbEPewZV8ETHuB0ZnEOH
fBsMUK2bVqqMZoZK1eB2VUttImT6el3gfOLHsDFoHeegHceEeyv/tedkcJZX5juLwoVlDnMLZiqL
RewZ1/WjpJbsXqXf8x67yNAHuShqpXsDBNDCAabT7O8OU6Ui/QDWeGo+TZk9EJPMp4mwiD4uGYuu
ngpOl2KpH6ASivo3r14pyxtHfSa8izrKcsZqeveNOreupgg266p43JokW1B7NEL4XdyommANK9Tm
oQgGex4OzsmqTrxnQoqyAU6DM4DVnbWE6Q4tDRb3WIr3abNdxNhF/U0Fr1uUJ9AxPUzOtugNjZqV
8heVmf24uAtokEOy3kXD5iy7cOPMJAW4Qf7Cz4JIjbzTJAGbv8Xm29GcM5aT/vvg0oWXqp+FBFid
LxDED8IS25/BK9X7hG9Aj/j0hGzkipkSUjpRBzBt2FipWROXTqNIMyPim/dckxruvTYTc3QawSMa
oOqJoMpsE2q4Knpi8ekQyxS22RygnZeH46mquLgxmILkrFhjemjNlJSEPUuk1cPO3YwRCIV2uM+X
HAorYmFEPYHIurfzqOGg0ndIiRI/oWAjiPegVItWiYJaah2QnhMs43tGnMf3KUfhLguPCDbKA3u8
9lkhW2NSAM1P/kmcB9LtMrujg//5bT6QPhtOb5ddnsEhOMm6aLpwvwNUJpdJC1cYOQ55nOqTeWt4
Js2ZckZxxyUV/uusioGyskuHjCKRmsz4K3H8C+OZnNHlzVoqKeL3IluR0IM1fj+M3FpWOnwhSpp/
esXM2VtjWV+7yVHlzXgBueDUfUSvqO/llkwfBnqhS1OqEHqCI6VLWj5jp8qv2FEdSNVusFJD2HQx
39AbCRCghEn0bnntoO4WUJLkIXBQI38Ew/PrVxBR4UFAym2TCPtqk+Ll4E1PdxsgyjZu2QneugH2
OirjgAgJP30ju1wv4ykpvpLqjNrcfUZrL/gGj95JApiBo2ZDY7etxJI5LWzPT42S44ZWJ1NU6phh
iuKc3KxctTQ9qGc/ZUgI7bbZn/PewqBD8PyFtL3SZROHazmDQpxVPrPyUYhN7tKIPm2+GAdlt9aU
+14cR8hFlaSUh+XXbLP3VQM1QEejqLevni/HKomm1P2gb8++Sl8wBiDAEKDJ9coolhk5xLKeK6Ul
VrFohptLosd0JomQIAb9V3hjWLRXtRy9O0EhCeEnuvH87GuCBReFqQ+ajQFtegDqQogIQXOWKYmb
tsLU79VTXPkor9A0J29i68AYvTqRKPgh3T2o+Qqr+HiPLvkUJPo6kMYRcJrHKvCU1LUaGoAf2sa+
C5yFzJkfF7VDi521uP6CUAJzE79eV4OVRj9aRBD9jkcFkPO1I0UlyDyldb5MrTpd3Kv2o16HtF7y
nXlDLc+tBlBd1JDEM7Kmw4hWCXXL+Fu+XTpHnzIMM4A1mzRIVwjjYXErEr3S2yYiHDl7IvELB5KQ
I1h3kS69oMPkpGtxrn5nJr6TPDyfS/+KWbvQXVpWP3LbUxwTBq8AU8SGeeaD68gw88eIUwhRsQRK
4bmic4EzHqUlxUA98epl1+VDHDBrJmuVc5KNHB9CZCV19Tv6k4WHnJPG2qDXXo1293stS94q20OF
kqNTr2QdTNhwRQlbNJFjp7FP6PT0fKhzhJvy2HRhdntRD3Gf/BDnP3S3Svd5KyRklFk4SP6NpSpS
5ntn943zTaT4RB6LC4Ne/tgVL/OYJXRXz6UFlWzSchEXo16oBJRMDmdjeDfAreUuc6+NN6Cx66CH
vWTSxZPkuPh7F4ohUHtKXaqCc+JzJLo3R2TBtHue7UKHpYGqlbNMJn1R6D5rdfI3yhrwFekhM7z6
lVtTpRteAa+wovnqcwFUHhMzqBze8gJ03cyTbu3xoeRAap1Z6am3Zx0CiBzYSaECDTKM40Llrg2B
yiUqV66sVfytakoCwutaHTaIfqo+IBZX1PhIdSnlh0FDXT7uw6kb5cOSK8eCbKZLNvT7ElB/94PH
yxe6oi0g8agSf43sh97FpIu46zSEbqBK3/7k/FxYmAvuNYPylbuMNI/4nBdb42LQJYb1UdZ2cI04
cENEvbIWHwXyHio5TxIjhwUYdIbFgax10nfFW3pCh0bvMI/6z3XOipRuFxSKHgvBfY1nvfPMoUQR
Gg5KyOaD5iugfgW/wa8xBTXw56CfEqHh1Hy2gTfbWgQSFuj0lANGJ5C6HJXxpmizLDaG+GfeLYlz
Ztpt+cZmWl+kX/0QfNBszEDBVNJPg6CinNq9hYDmHk9k8i6upmFUwlJhFSxAXPwTv8etFseDoOkd
CmYW673DoFoiFFIqDhGzoCKMJFL52Em5Ae5ImAbOIk8ZollVewvFfAVp+zlfWlqHzTqGAlD57Br6
1uJ++H3yUWm3IIlJyvXXKTUgIQ7w4NsgKVmp+kXmtZdaJgMNvihK3GG+ESQmnvienH1tz41wS9Ui
B9vs7z7zd0mK9KiYLXR294BJGQZn15cQCmP3+kG+mRHKFnQPLleQ+q2lsdEeaYtmFwoI7wm+1h3c
0h3U6sremgwPc0L68vV3feAbmX8izOL6TXL0/2/nHoa/uSDfVd5wLlqIjC2paw2qjvMb3H+0sqh2
mFgy1TbepqG0W3DPQprLzXSojmS63xyx7l39f/jrt0wIHuUdgGGJS2Skd3UyHfbQUiiiK8PKYflf
Hc5sQlDzl2TFM7R4DrTW9tMmQpjIskClKVBYQQIP2bQDUAMeIIwH9l7x3xtidXJkIZE1f0A571RI
nDUxI7n2zpXPGWzdWSc39g3uIbU6LGmde/imBei9jKSB/T8ZuNqAGGJjD2eaKSFesCiDc06q14xu
jRO6wWQ4UzWGhFPTuNON5uZYCdE5oGc85n3RnjJ7glHvK6LXyWDoNFPua8AY4AYSy4JAziv25sUl
2QbAJnjjSvt+d1YHpiL7UlKVqKmxGS9XU4qFxYRuUKo/zX10Yp5ygYl0GOM2vOGcby+5yIQXAV9j
7Vhv9o3VXh9r+Ml0dSRBiXr0CkN3AM9i7HkopHnYCEoM2Oq4/Wj1Ms96e0oCk3AcZZvJ301U+6wg
pPrt/6HTqTJHXk5e9H7P1975H50mKyhB+RZG+yAAyZmF8zerB6i9ky7eiSruhw43LpIwrfcOr18u
89IxTB5lrZ/8TcUbc+KLoObQxXmQYIlMGHeUR/+m8JLZhDcftbSK0kMK8Obt0f1FYKpLh7enHLiX
V9EJeJ2cBCCvpFrJhJLObNjh5QFwPBI8PfOKYx8j93fzgMhyeYR+jomR2ko2Kd+FDhFbGYWgg2ud
tWuD45nUACJ0+csKDNrZq+5NW43hUWNVdF0YgrprOmZ7L57fQIHu8enC8Pa9ZpZaT+wggAilmOhV
2zbx1S6PKFOPRcZGCklN6bl9IIIxVGGipM7WIPrae2WYTBr3AB1YDfAT5wzsxqHAu+1sOhrA7q+r
RA1zVvSWYvJ7RgFGrBr3e8ph+sm14FZmSIQwegZB8/4AVPi/i5bbGK9hOfUjYxxb++kERjHLoTcp
LmRjS3XVTa1rsabr5gV3WVNJFo53IDnllFbanWek8Vgd/lOv/l0UiEpbU4YQX3AHM1rOq/aaiabf
+jY2TKlPO42UiXIqvilGZzHOlLDuUmyCIyWUEehUdI0sUoy2YvlPz00mIEBTloedpjKjALjuXaIn
YWbGYvIRltorsynkAOG9ioZzYTg931B3bZMA0Z47mzNQy8QhbyDNK3tv+Iozsdrjx1IKoziQaoUS
W3scu9tgSkMvwOudwVhksstyi56nVqcVEGjAvfzlFUKMC1nkhRpOdOCHrsssWQXunc4/PySEBGNq
LWZGU5/XPjIm/+Qpq6dBiNTq5oD7TgOFl8tLK1iZgWHncfLynmhFJaYRP+i0vWSPK5LdQZ+uJg0c
m9GHWtcG+uzq7yXlDNiiTZW9W9X06x2YkQY3FdgJXpnoN1UtJcA4QFgcbYwo6LozD1t1JnoAJLYQ
OsLF0MMcrMLz8idmBQVSks1Zv+RUAanhJyRW7fCQWlHkO5kZWSKb5h7Wq2+oCiPvEefDH6me/aEU
5LXwZ+pqBlHK4H4YEck3RMn5axdaTAJzEP2bInFQ4dp4Zg6gZ4FVwF1PaE9jaP7DYoSDlAKdpwAE
qNAF9sRaCEbv66Cy51hag7c/CFdC8GWzk8rPVL8SyepDUBE5+kdoa4n/+Ea2ggdiUW7y5cAnHM0q
In1jlBANbZYgAPtULIFG/aMiRI7o+u/5uZkA/APcOtAKB4gDlttp8B/ZWrAPs/OpK4AfIwOP4Pmy
ZAvCQUY9XWx4mPHH26SHSLCiSRkql4GQGEixVOHeV4sXINdHrVNhlzF/bXPxOA8DZ55HpnJ256WY
5Dbo7Q+SnBk33koHpWhO5TtFZ3LaPZfV42g7W645QOuCeg/vi9Rv+azw7eGdCPvJA+dOpY9ThpdV
0/+KylThIepytq/ZVUGEGhAFCBQ4UoVlgyKeeQJ3csC1hziYD/2WMa+g7345Jv8vhgRpFeWQ6o/v
nB3qN1EkpUNBRHcYfWcTTuBT+vdDw6oxmAON0b1qhirVRo5FszOKm3+qTcihiZxGPTqVkXIUD+zz
cKeOTxc+rQwoo2ijQpQqWI+qJaynWc4I4bUHivPQYDQNxeqKIkMp+5VemUsxN3M6NgSCtf2norln
8iSmEEPUhrs0h7RszNfGk8uZ/jpmp8zQZ151ZdbTLoIhnArjwIUbHEcDumgzB3uVTc2LUbNc/5vR
7zWzNn6DxYAEsrhJcEJDSyELQ+NsdUtz8LDvt+7rOdiAYYiuqk9lfnC5I0fugZIvKQ4v3up4f4es
zxIuPk1rGHkE30DqUydt1lF3BnWCsfWYvNkb7m6eMkMxKZ2rEcrWQxlITJwZxl/u+Mq6IvMYrOxc
k1QvI+nVICp+uP6JmzvEByoG6bxVdchXJmfO8qP7CcB2bqd/sBNh8zXkSg4klyBhPQXhgSGbYdcO
rTOsEKnaazbh/fXIklDlY7JYRXtF1sOOGENZ0y9Sbsu93caNIfKIlZH1WI+mdBS4l1t6ltEFNWzi
84HtnRFiNLNTT4Win7YKjlptqnYglJyuF+j8rOeRb9qLUCgDMVgLBBeueG0ewrqo7lGHUlU/28/8
QV37yNGrqMY6kZf9DmIobxPMAV8MZ0fk2e0dFXApGW636nkbXNxEb1ZaFNHAdWKFLg+TiqjE/wQr
MSUBxKKtlprVUU1plLh3TMxH2nW9kdoBw2UtnFF2WRLwf9t9bK9aF1Pmq/l8YCBi5CTtOsZJeTMz
ELFG2lpDJmlm7fpenFvUAodBSLdMUrWm3UM9rbrtNNBw2q1bKy4ZOvCxLCx3CXP6A93ft2HD5r0D
QFzTgcOOAm+WZPdNxqr6z1GS3SaIQS4OuE1lba2WisTu1v7Fb3/pu2SpQIDGA9p8SNKDviwsjDg1
Xxa8r+yRLberL1B5otZI81tw/ia2fvU7u7PpkYnUlZIg9tAcx9hphV/jaHqEx80zox9eHJKD9SvH
BZwe9ahreVsI6p/vK4v6AOnUKYYOleLrCySj6Y11vHZPhd4wO7rXdG4Cn43vUSjAm5lamkuV5kqZ
6imzTVIKm5MONnoOKEcAye+MTXrVcudaylvi57UbwSR0uMpDjfDOH5OuFQg15u2kxXLtJp40DgTH
MwcQuzFJuhNoYU1l9zHhVXsp4iGrT6CvLohmCWZhkzVYeRTV14+6JoTrLpCkSpNggFn+7Ma2MQ4H
1jdZKRYeuGLsIf4KAdKSYXWpkHbEHHSZHgek+8jWuMp/7b0jUzJihQDqWROyVEqudHA5FbtilqhL
pQlUCXI47A2+5u72VzBjY85hHukdQ4ibH5iLc1KS2ARI/NqnGjvkWl+4w+SdVH3iEWicOPszrum9
mgR+YdbT6PCgA/a2fHdtW5HBSFNiAeGh9nqZreeTWhluP+VA2A5j5tNcdUjEeRc672dN51xLoARS
qeoKVNFN2oc8Q6WRtUClG5hfhdHT4hvj50+s1DMPTtBnQ9a1Br8zjNc1cczllxCoU5lCdfreiTgL
lVm8wipN7llAC+uTcgkfbpuAmamaec41i15c3iRzBAEDK8VpwFCtkAANk8chPMCuHRyjGGebRigT
WyZP/uCTLkzG99IlSCqM24bob4FJxH+bgKz60Kn3b3yCQpy9tuVr6UkOa8fVgDauWK7CClCkezHG
NEh5v9p602B+B/deOQZse92z61aHb0KjPbNjb9/SwJ2V5Dyrc7iy7N9bXYaHfElEX+899wjI6dHl
AyzG3a618cI96YzcbYCKqiZSpxLxruLREhb/f9no1nX4VVn4jsv4jzhcRtvNqA23ZpJZLiDoGO1P
YlshCK4ZLIXChzetE+3uFeGwMH4MCW9cmSbhRfmcrzC2vECTYpufCHlJbupyiUiBoMDWpfrFg2p+
NHpk7g3hAb9BqD1FwvKztDOcWxM4Vzmecrn4Gl6tHiMJ/tv+XVLy1ElvdmGdR5D+3w8szjQyLD5o
fHSLhQViFKl6CdoOqeQrXfvkm75pMoIqaltGZY9AC10MlAxVIqeC3yZ7yP8X6RNVHJLH+VQJI/ne
90M8xT2Q4yrQlrrDgBAGjOAjBrMDobpytCw+48/5D1H/OH7A4AKCyZQZq8fgI5pbkHplr73enj6E
PZ/KSfyZBHH3P6d+MePA0wG6xuz8YTzgWcw+boOmKZ7Jl4yFKsVJ1oHZzcdKygWPZ5QcrQimgsJ2
B7xHeS5Wvcz9rBqLIDk0UEBJibUR5dNTDhswWa1jYNfFuRJc3lda5xSIBtr8Y3Ma6683bmUnqM92
XDc0ScSLVHFVpLTeHikKzmNHcL6EzKBDnXmV2kbKpVfB9a3H/JLf5JWcyBrgXZCSyQSVomLK20cs
CB8tm1Cc5qlXO8PcCo57lZRlBt0m6zdtP2BEB7Q7QxjrNW6+Grp2PoRevzssKhR22/GwPindTQaQ
wb1fkfr4SKQ3vYGfhfvYaWr68tS/ml1hzuZQyYPMakK9Yj1uu0SbgEYYa4x3dkz39gXhX/12b+HN
bsUFAL9uszKfKwcIQ9n69W1DtoRTwcGOk29CXW61M5H7NDGLM6fBpTN45Lo3VbREfIo4IpvlqL4g
t+O8CUnXeq2bCSWvCSBOew4KJEl4wPYCxEMoy1bLeskSfY2MsL69aQMSSrlX2KTeSxf628Z74BMD
zvWmkABPfvHMyriMbltgQbICdXPlt3YTsnDiLm1PfWmuoo/rORgleaxTp81VKNvBXrkDucf32bp8
18QnUpkp5zG63fXI2KHL3wYTt70tZDXWH+4fre+NK03IkVGIhRaPLM7Qr5W1vnWeBURTcZEsVhf6
yc0LNEjAWupyWmq3bSKXnh3KIZB7AA2GUMbkEhh+vdT4XtTYZ+eCeyMiPx8Rt0fQYzNowcV6hq24
6jFazWszplBlIYNxX6sRWySq+tyr/CHzlGneFQVnPvK2r8wtfMNw7M4Me6SYAKS1CcKMRWbeHIHG
Ht/xxms1rhB9GypOuJitTTycZZ2CuOhrctNsQgBTdyS/6n+7lWLk5dkRPXtUb5XmQNcHXknEgE/c
jmFvh9/u+KGKbEAvNe2obFyhF7BpZ47yGWQGpmYgyzEwRI/6wVf91rupeSKtcKwqF3hyn+uV3m8k
n7vJ3zCGD3wubi4Z13UIj4lzmqT6fkftkwqLWmwj2xw1SISF7rNN8wB1dhfzRzpd2u8QKGR1QU73
U/joWkYp6mN9jApTsDf/dxlPcd55HJbAYgbbNviruErXiafHimWRmNnT4VhCALplNkcggu8X+JPY
OOtdFngIt1DNKjRR9ZzR2o+1xliiy1gTW6jM1OMoP0kukrP91vNu6JVDCsqNzHDasnxJoiCbso9/
I369qte1E6InFbCe65e9/hPEruiHx/QjqnSLU2MFPJf1Jej5bLTj6aTrZQplmiSdvX9eoKiH5J/s
W+M3gasNi8HTVtNFp9k4KPA3EnTp72pA+YtdG7gSR1yJ+m6m0F/QvCi5Hj2HOgC8p6ty3f6+aK/0
Ig5alQmwdJkhY6lm/pbGJR7G1aWC/xp5D1wVh7VR7BpgdAISYLa4tWnaAa7uJ4KajfCRxHsGeg2w
tu+lH1vJ3RLeMEBucnddwqwt/FSxN7zEydzZT3YHhJ/L9NCLWqrzXoa+PDHc0IU69u+EEqO5ugbR
UVbnwQQPqFtfbmSXLix8NEf2RXGBUOB2DkNTvV2w7uLBAY0ngRxMJPf5kAW5KzTocr89Ngo25vyQ
t+KKuGyPiPjmKGaGgYQRHvt6f5C978hptx1319qs7ZZXgdVWn+5tdrh59wURIJvFqnWWU+qENF0B
v98JvlxGyXBRUd7PGZcYksfKed6+GD2bEm9y9770HY7y+SCt23XmV3lZvAx5XqtO3GW56zAB0OEY
+CkM7nkWwmgkDN0A+TNAh8qGmkguA3dC+kVWrrb2hoBhtqutNbwI069J6nVRWuFM/trDSjAQLXjp
XO96j6D5/73ozYm79OeYsc1VxDAFnvmaBY+Z1iEYy743Yy0q9a6z88OGnWmzEL5jb8wAUjkhptwG
564kH+IFsUJaRyLNKIV9Og+P15MF52Sp9ilEsXODA4b5kJzOPF53SVyRYN6pNyRPYGWwj/KKlebT
ZEncEk8oGixnql1RZ+sqtQhsae98bRbGtPom2eZjXeXnEPq3yxyTjFa1YL9IlcrJUi/7XrgHwFkK
0IpyPr5dIj6ONPmYlAuPaxxVONgj5xbTRHyIGGyLNeA8x8aBZBhfRxIHDSrT+Cy4wzwETp1Zdjzr
P3OaxMJcQGndU6Lsrv7Uf9jexjIqZPFuj+zp84U8kLKeoNNsK+QtmKKVAdHpVLTnsXn/ncdQgrxU
ojIGUi9j/Vux1dRNEdIVaVmM1MLVRGK2C8IXlaLSKopYtDjwRUGhmjeCxMSk2xPZq8+VkqnBZw09
JZZGIsWhl2jSFySDTG+5RK5TmRjhgnXT2xu9wy+61ZtJ/2OoHTpDQOiT2IVr01q0sRptk+BJQ9qO
ZuhSMLnGELQyRgartHWFWi6zhJj143Un6no3KfOPsPkW1s5bFD2yEEaGgt536uH6qaRbIr8UbaFA
l7ElSyzYDwUBjSBplHuAEhj51ezXA0R8aM8+JCvSPXHZIQQFNuuj4E41Cn8IWliGkhV4u4hEPjrD
s6qajIX9GLpDfrKvKlnOaA+1JgpJPuC2myjPJ+ZxDcYZAut8UDoMHDpvhROLdGhI7QFWpdycaxdb
os8wds5hKURijfI7YqMxon+IduoXXUWUIWWvqIOBsDQIFENyRxvDG13aZQeYq8l2moD2P5fGauv3
n2wPmTjs7IyzC6wp3HF8aO63Z+JV+5FZDD9ZCAXPmiJ+xlP/M/28g/zSnfR8mKz5e7SnmUhztzFJ
U2ZQzrA/mTfsAN6jzyuYlg49JeqZHJNKKRlWH4etW4b6KRsrcjqL/gQgoaYgTsN3msuxMvR7Vg01
cjsMzIWM3tP7Hw4Al1z4OLsHvbxH9S/cXIcbXtSrhh5kMmmyIjqQA4ohFNntBAdY0xsQxoorA6Ug
UMgZDepmymbsVBni97NSDD0nkJ5Pq9Wfk/m/vN76InRbNLexw5uzlRC02BBrX9Fs+qiZEAp71w27
xi+MFTSCDYKlbfSkdILWXLmytCfiJRoDO+25S2V76Sj7POcJt4a8r5q+7s159GHFjknTAiiRvawy
hkc+pOLOwkp4Ko1MmIQX1D87B4mLk7dKx0nZu0CmP2vLye1P6i5tpXuyuUHrYjDup+IG0/wFMM7G
Yzq2If9OHIfauk31ZHj1s0PoKq4X2WZvOxPdlq3dgg/c/FUFFXyaFFj/jYQ9QaVlhmOfMReVETNQ
NHZUNv1fUr4UHDyXMNqo2805dLpmuaM2yWL4R50p4728N9p8kDGFcHocXjar+gmGRGscn85dh+6l
C95cHb9uacpCsXD3YoGfOZ6zGYnUhSDF6dXuBHbUddn145ZgXnlPdQoSEOQK7/qmPaf4dJg76gJ0
t36R74sJVXiUIOyaNdXQsmMF30kA479L9qYHVruvHb27qnfuIhk7u1z5cTF4zzVjnEal0fTXtZMW
yywXXqR3yNY+Kvq910xBQTgTpIGXF4tY5LYBQvsh5fEWTWB9HiokBUidUHyQuWsoZ/gC7q4BuFOv
puVzkpFFmPLtGUJFueuZxCJrlcGHFYi7MkW6qHOQRTK+E85neOuSqkoLDUA/fUiSdn7AoeFU78xy
4muqhFc8mX1No49TZpjPLjwPtK0vi3UZ+YHHYUcRXNlBr01lRtYPcrN5akPyGZrzpxhQQczXLga1
6Ftplc3XkqmoTEseV3z4INDyWgY2k560FKaJfzPN2XbFsB1gwEBBcVlU07Kw5s3Z2WKkKegMXPd/
psBT9FQJ+MfNT4s+uhbXCZc2E8Ctzld517ibA2D2szBgQ4Q/2G3r8y+TV3XZb5+RKLEdPzQjUp/r
bLF3SyLpPbFsaMxqxnmYn19zNcJmrD6HCkkx5Qd2rRSOyLJRZpAJvcVVw1/hR/pnLyemKwBIBC4N
ZGPHIwyoICEC2p6EjyWM9VfbMDM2pR7iryEIkNx5e1lxqNeNsqNC3tcUcF4O+CLYTiEc/+0YQ1O1
w/RmBx2DtxM2+1BBwPt689ORbX/ZUQa4Bo0k0TccNuqeW0LaaRgk8L6Lcva2ZLj8bJUUzF4Qbo5M
SLwyUFWkb1eT6Bkmd4bOf4R0MW14A4aP2XYnta7unEJBH9Ur5HiOGxqQZ3MCTXVp4P4B46mUJ/bf
yaplc0JAQAywYliv0/3t2hyyGAYypbQ3/d1DmaC3s9/8eASr2LHgu44IMLuOWz0mZzXI/TlEQ5Qj
JYzoFlJ1I6tZQQBnWVmOnqJXxfEV0k/RKix01ruya3Y0ss3drdNB0zguolwxyBQ1V0tHBSFrbYr7
hro4C4/pwXoPFhhvvaakZOQ3/e2Pz2H4cU6yoWE+9M4mUe9oxL+zbD+ws7LNMWDmWmAB2dtPaQFc
2eZZbTO47bSurkt2D6lLy2Mg+8hJczcZnmnHM1qNHHp2RiiVeBS++ZQ4466jG5iSoMZptme0LHcI
wkCyrTH76TRbWHyw2jQ6EpnFQLkxyTWRcPTlycJqUWH6KJN/mqK2cgnX1cX9nRGoqk1HU9L5pKQN
lxzDMH2RydKvnUal1r8Q1vdjHilxAM++QEF5RG+XG+MaHqYTGdFylQQ1CgfpUOmNJLf8PBd79R+5
qrd+Q0C4hLLPaTvMJ4IO2Ad2skkRN0zuSwIQTkuK9Z6+dN9DRz/zcWa7+feVvewr3S8U6bteLaMe
4fBWOBGYasFN6kmkhRBS3JwPojeeLfSn8BYYAWkZd/iPaNzny4XdgyJ/C9ekC7l0H1r3xDvUPdLf
bVBnSbeYEbh4PGPI1kGvvRdB6QHEkqIw0hKEmyL0RYortPCgHac0yMibLPiLiAGbstznHp1BzGEq
bwFJrrECEv2uscMCKNMXddOtMVTwxT226rar2zIsOxdO4UZSsrORlhooAkq0S3pkpueMgzBsiG9w
MZ4V09LMt8tKWMNWHLYk6TWws7DsYeSSdylthYzzRTKunDjo2fXCVJ/PgbbM0su5UdiQuhpw43df
JwKsm3nF9ic2JgZtvePRFCI2bkRpuKNa1xKmmUdf2c0feGpK6tG62D40kwk8ya2DtPDs6MHYkdOM
1zcbxZwa0nB+HRRjKyZD/y/1BYhvcrC8gqyqEm8lTFOXXYCHhSlSq3PvgXKDChMJN0NWNrqwrGvS
bm2+U3F0ucBy9Af8wLAuRU4z0zupL/Z6LoVC+Vyaxeutmj7lWTXL7+l2hdwQeYSA/iFhGFOV64OV
cw1Fc4vfY0Q0RunSdkoglt0TtntIyQS6VxGixWv8dR7kl+EfkpsaREyn1/0dir+6opM8oJqhswMR
OclWDv3zhyrjhmh/Gmx9YuTY9tUdnRhXkBt8G4YL51UMmqvpUq3jkU0TJs4AZGQzLtYyRBWiiJ3X
+a9cjjSqADYMctfvjjIKuL8oK8xcD2h+gRjWiRMz2NeEwfv7ADjzFokncT6QXrcwqpkWywE3QeLJ
a0XiaDxO9cBY4XzZMIvNwmCQe+1a8xKkZeh2rl3oyWwcv54AmndAGWW1R/677hUO4pNfd/tQVGMQ
imOj4vxft+VB23ZviAKwdXueXZOLrFCI/Y79udEgNAZ88TcPkROeXqoKkDXuZbUz/j0zjA38vjqX
R2yrMhRoQbBBJYmV4WPs/vqkhPlqbsdEoLBHjmbmyzx/bFpzk5MMFE7H8eeGdcCA/QIJNzTdrbND
e/weyZGkincuHcaAjdzaBrPxxN9r9Jo2a8Xbt8Y4aj2Nh/ecD8353vnFRljyfqaRu+bXyAUC6mQW
sJHx63QALIMx44EMtAHuXPHs4WXeGj6VgweSpZUgcJMgcKbq0gWdPslR1YLgbk+HD/swGdVL8los
hyxvU6PX2nBzvz09DFOA1/1b1BP0wIe/i1J8/3J63Q5yrqr5T8bBN2/AG0WUgsM1crdlBbruWC0b
2WCS4t8A1OUQW7zYPrnqgMZu9NL4Gn7f1w20M5FRPBF1dfJf8Uj1HtkRefwXJpz3mVzmTPzlxGfx
IA1D8uy/Rdc6BY4JYs5c8VORqMlw1zEnSFrtuk+SKyN+wxHJnE3MIPg2Xq0/ALEhIHaAfRynC/c4
zfrMCcM8m+Y2r3K31g3MR/tDGz1udLTuO7PP9CTJIv7hAKSAFk4OEsDcvyNZzVaJPjdguylEyFh6
EB9Bo42JqnWihToG0kER+vlmn6Oz7fQ5cRTbAxcSu2ycLKN4EM//yLjZQcw8nkEBMBOQWqtw68zo
inXnHgn7leBAYME8FTugOgBFbUOvkLscpV4rQDQsNPf/Yb6gVKf/cyOqr9wwkE0Twaz6wfWwEN8A
LSea1kge47mK6eUqTq7kuXThnExz+Fy0nBKjWNYkt2oULQOL/6PFPkLsTElpbIbajRq+XNtQdj2s
Rh7tmjskdF9BY4ZhclRi1LkjyCYYNmlNeyqYzCDKdLr2Eezv4EF20Xaootn2l9IZfrp4+51yY6ak
ng8jzbuIx2bOJBzod3QVYHV6pcKmnFvxaCIXL9a1fU5FzLpsAHplLCsZYMmFh5DfYLym8+0cTTn5
TlxbyNOvtgcZ3YC/fob5ie58fyojyTLBJ32P49CMVwxS2u8LaS6Zd8U+LUSr7+qWzrVQ8F/XhHpF
NxhZPptFjCpoXTJ8i3E9jnwnyWiaEC3HIfgmoUA3ZlRbeRJ2BnF5uzvZ+dLJHxizb/XREefWNuJc
0m5dfYASN7didMRovNL48IFeY9ExpN6Qg9vqqyN09tCZ/utcUFfwNAZP/0Agh10b6L1Ufo2oT0k9
lKoMt3wd+IN7HAFWSk96FACQEyQV0DpLrnz4V+z/BBWfSnBAPVWd7eAFgCbVeDaA92nv5iIemWQc
woZBcigRF/XXLMYS+9715Tg5SfneS91nMnSDGBj0DKGGtTfI/9eL+PJIQX0qsz7F+WipkflvO7wD
qA7t/hXeto9SADHtyWwGM52H/6RrX/Apv3bDHwv0ebesIBwB3wfh48h2NYK50LAGCsXDdH8D5Xln
7BQkREnj4BD4kDzpZQZrvzmuTNEmtU0t9VT96RZ1zYtiEqI4lyv9rr+JphnAogVuHUZWfOwQMlxS
j6jJYEWYkomv+o2N8dnI09GUlHA0EylfTfuzEOTagjENiKVMGrAHSOkHWHQpA3J6YLfDDJOZZ38Z
MKGFp3fz0RgAWMSMd/J153irYauaiU03S2smOaWDSJqDTYdcUtGfNdu77wV81TUATjZyIf6IwX/P
R8sIrCsmPGD+SJ+DzmvK819OjXmfPLQBV3RwoF4hcBuH1X3j792AUA0AA7ciXOHg6Rclqj5pXtGN
oiftr6fwa/sQxcnySJxm1N709xAywWBgm56Zm1hY8L2bvtPy3Gs8Bt7HPmFqZAP7ABNvHrU0q/8d
wxv9PG5dgjB+BM0pbBX40BIGC+9bHWFlFhFjVMKTvO/0OspPr78/ojgcxnrAhW5rv/zrZ3raFFPB
9BuxE6ih+H+grLaiio+LwfalUd5htcb3skhnv29nLGUZT6VPF9tDX2EDva3mPFWKHVCe/iNdZlaw
uFgScfyitFm6ektC5cIHQ3DZCEKLpB+BfIkThgVdeHYJMYBl8fWbCXoOd9DimaOTXnRJcqJyCRMK
ndZZIysN9+IyDkGANIecwyOLnc+mbHW8RxExjdnrAaaMSycYdOODjA5gkSoMNNgpFK93sZt62Mlr
+Rlsucev5CeLtENLV3z1+k0CiejCNChIW1DGAjfZgvG0fE7EGoblA36bR25K/zFNbWNbl/WEVZOD
XkSlYQ10nlcbsHCEADIeIPn+/YkKehPVUBcC/jjbZM9taDaXhqVOAu3JKDZ/Z3rqJyOXd5/IgYF7
/wgRlK3LYlmcoS2KE77DGCIh0S/a8dAI4nnPl+2K92DI8UqCBBb4ePjMbuysw7GyOr/aVtWDVwjL
p37HzCQl/qu1h/D0GuQGnKxggojQHwnhMVgE+odHXvMEsR4cUAJMly9sGG2XuMptRVA3y1dJplbU
99MwCMGmsMlopiRjxpxJkam4H91gWCxwf1FIDF8QZo0KJ4QrAnv9Sd+pLfSzw4w2IG2PupzD3WNR
gLHMCjIsBeLUInwuqFtXqGuztN/dJBfM2k8lUKrDDTYQlPlVNYmfe1CtW4htd9iWD9QK0K+kfBum
90rToukkxJnXIxPl1eqyvU/JazhIoFMhpLWz4zTIbaGl2N6wLiak0zg0aOfK4Ovz5PiDoD4xO5pv
u+3dLQuCCSLz1CzVGSMZY/9tgFPjeUvjsj1thJIIX/vYXKxaSsASEJNK/akHyPA0oOdHoQRzRtyS
bYWZ99C865QxkMXIJUVmBdXJ1xVCX/+EXs3VB94snCZXZMfzncp8HTF/72Lt3Nm5j9PQTU43vVm9
9HJ2uF2pqiVkdexmA2fVFvYBjdSlW3r+YWJz2TS1SfL2QFdrffkImxkcb4RP00P38NHRpzPfprTj
iRRjx1YiKDRk84gicpORDZQ24osGF3/ZrIEgWmrwl4hEXq7uFNN5oddE/bQxIBw3rSDIDMUX//lH
E0gJYq+a322JzCl8rSkM3K9dBxEf2bGL7Rf3YriPX7xyH9QSm/x1lpABg3wspZPb2xXfdWIZIYh5
Y7iq6RdV0mwK3VKlhsqDJ0dgZIlRUdud6ERjt0obv8Tbep1KXn5mgYeu44Y5ujKIhGkUBo4PWqye
TTVoaOhEtsEKfYcFkdM0mx1oOrkUz88hxPYE783vNzbNYrlalpqi2Q21QscrLsRafacjqodlzF7h
4HVuQGwamLrFcG8IN8CVTlt89azpRKdx4DE8yMHXUvYh3uEaYUTZ2+nrBV76BU1jXLFfrpUocsn3
ZBBUUqGbwM/kAPtkUaxO+qocoV0n8KYKvNu6TiQrg4qTpua49bvSOJHDmZltyCiG21vGV+Nc+3t1
dtyjoKvG15Mn+P6oOUV1M+J8+070L3bQGU+NHyCi3ex263vnX4kyHsIVsKp2IJhlvT1tIfd+3MAq
bmbTC2YLE+QCJ8+iLheZv/IPtv9e9y4ICiF/xa8G5zM12aP88u10BAMjlJe1+3uSVmfvWKQULtFl
zeGPWNMIQ+yehRtzVJ41qji5++yen4w+De0211yibafR6nKuyVyNujCIFgiPVj7BdcRnlrPXBJK3
PoMI6TY1bKQngj4bRRYK0NoR8r9wCGCkzVdEj8B/tmCuRp2fNNsK+s+bsYxfusR5paPqCY9t/XEk
c7/RtTk2jZYldNdbMc/MvUQ9hdyU0cRTNoumdT6hwcJ+RBWQrA8feOYiVr5rENCtni0DQ/vmvy6k
AtlWoO/Zd6sDpK8Kfbcwh/YCwxz03+aiAvhhJNPLdZOCyZhN13wzLn+m+TO2nX7Sba93FahFimqt
Y1YIQf8jaSS4tw/qbZvg5wc4x4Vhr6HCrNS8bXJtOgGYn4WfOnVVCMf25dw2dIM6SlViogU5ZJXM
bNjxltSz19qnRkj1NtWmdVKRl/CqoiE4IpO1AFFXrhy2KUE2PTjoc+YAXV2tQyQhKQQ8zsYOCvNV
IsBbeNkIIoD3QGS5wgjriMcEIMVSn9FmYkeHB4P+eZyxlav0nXlZaIfjSM5MHihRPTZfwcQMXuJb
xwziSItQAmk4HKL/hu3wwmdDgFf3olg3R7sODPCoXr4bs19WJArKYYF03tL/el0oneUS92Fm86/2
luA353EsYfZG8dibOmzY0TJZ5Bnya5V56zKtYyuEVhv9hSrcWoHSUg3cDYQHo15bNBGW0tuq/b84
ZHoCoNdPfp6ydDtfReSwZHU3XLfBv90TZNufdXTneTAJItfG+9r/CjxSqdwpOVibOu+AYCPbErEr
yBG0yM4CYFR8acsZ6P+o8S2NwNv3XDxgpGL8RfSphf1U+j63mBFJs3MjY0v0GQNuHQXNDeENB5ra
kaBDd4fo0u05kNyNV3/wmD34G54kijrEUp9VpgK1Omct2et9pI5a6bZbkNO0A3lNvYN2ojJeTiQZ
kqkST3pZaafcRdBDpT0sGb0T0uCfFiTrUy6IrctArMlVjHkfP2oL+b9F7W+RuKQDNwI1JNh/O0n8
OyET2rincwZ0H2oyLsSvkbOc12Xt52Ptmu/wdHvvHX1F8E0cqD8HnaE8xeji9OTCFxHl7cDUnYRC
Cf48e2SQTBP0IUZtWwSIWc+cG4MRvVer5Dbq84Knc0pvRw7iwrp1Ldxt59rQPJ/QMT9EBtpc77j5
Ux3ZBttKhyqoVHUSdaW57B2VfIOp7wnu+2vRD7z82n9dpNCW8SqD9ZIgCYkG6vtkKhHgxOlgkG2e
dSBKkH5y8d6iIT8qorCdSst0iiAMdaVoOEDmAmrh6xehb3BvywubtqgkvK4CiVqHlucN6IT7buq5
zW8j7m0TDYjJlLJrHKUvfkBX3+SOXb0RQ7HKR4//jtxs+5ODDwDsJslVc1ZJZNd5q863JyN4FSoD
apDBpf+55hvbTdUl03QKppJtX8xKlCo3BackEN8SmGbD7lnPg2WXLgE2T66sQpfOuBpHhvgVzC8/
S9s05i2c/S+xlFWVeaN2yleHkDjUMgkGC6fqIxh2ei0cqPGdbtz/lp6khyEUYZgktPA0x1EHoPTM
Onlk1HWExo3pJMMgzcR643w5D/vA/eVihcUe9n1tyrMwxCqOq2TcHJyNFlHs3pUyN/cie/c3W0D8
B+xl5Iw+LH5dt7ph8528fc3BQiDN7MXcaeBlBibujSdvj5qNBB9MsOwXaCc+nJ9zjWM0FvxCUGZB
yWFITQccKvS/cdq70GXI4WKl55jtT6d1K4kCSw063ekUYlg0H9rENicH43LjZ+S3+VP0G0wDC733
74aHAqDRcp8mt4yfBfG2oL4QL9bSgwNfc0ACOu53IW568TNub0PAh6+qBWOiBVJwcxqIEiJHK0Zr
ovA7CfZSxdFujg7wSuNGc5JXy/nw8KY3tp9ajnHJyeaAZ4bb57Z7O/QS+BE8zrDOZTIo2Zx9yPM8
L5Ia4UEJjOzwiLuyIrtlhaLMpRbBkkbPbemiJ++qllJ4ZVvRzqzFJ2Z8JI20n06ontAcJQCt4hFe
VdGdZmAYPp6L4lOciqY2tQi2X147EdptAVXt74daEdfHHGM5ZU37ZyanlcDEmybWp3PuOUYw2x7i
EIubifpbyGlO7+IIFE8eq/w5D+jtMLCMM7DJL8BiVMXcKyxPAdEK83IShM2pw2+fRp8/TVcOk/eG
Uu/nS02W1E7JdjNS2y+H0Wk4s70qpAvNhgo4BlE3uBQ6LIJTSiJUl7ZUIsuczWCgFlFsFMGMX52L
QQ+76Aq9SkXhg822W4EzsJOzGmOUtAkPF7sXU87YxUD2lGIbsG2KpE1pb+KZ65k2jSNOmXwkU+Nr
s2hPgGiOZiAImNoysX44yAzVmb5+uv+1Pti3rTcOQazDgKwv+ycQibn5D+Rg7tRtR/lzRflxpVaS
cMd1xUtdqCv4f5q7UR5Z6ZWgP+E7by0UV+lMTmbOIL+pvsLp9FJw1DCCiG2ETyy5OsHDaR8L5tr6
hBURMqMDQKr/5ZqsSC97WA7L6gnwMkG1gxUoMwmcndyE/fY2ihcwaNWG/4blWKJovtfnugyLY4Oi
fYiqUwm2QN1ADYGnFU1cAuAEb1+i3ke8fpbWh7dWMbodcYZkvzAg/EdDncjax7wQO9aiK7/wkj8F
uDJZ5d8m7xG919hTLMQ456qh0G+hbtyI3PSgy1LdBwkYABEugG11WCMgBf0gfjUZWP+GZARaMsze
N6X4dXc1ti2dQl0oO6cY/eJOZh/jBmpzFEpjvuaqKhKgwLk3XSxwKfwCDVCwdQwoMRsL8TRcsKuL
pJAtPfWpCBFRq1d++ardGd1iOGjghHNHJpaeQd+ROkALp7up7PyWe74MEch3sxT816wvwW29ln1u
2aY6v6g4zRFVjIC1eEsE7SdLpMWwoCiNh8+AxWtia79qUuczzyaCljddmbzvNL+j2SQAZU0m7iZu
qv7JijmUCA7sJM3iHrCRLyvoUGNs8IZMnuy2aRLaxC2/QEB4sdLOfNiTpoXFVxdYUQtq1aSs0zTE
VorjiRrxWQBB57Nhs7R5pbNvFrXe7T4MQQLC7C7rG1yL8V8cApDFGm/2NVFFh7wIqyabgbJPAiWx
0Htw8syjoONH5Ti0wkQu16umIe2TLHediZ5nq+ZLeTl2PCotgZtH+hZO+SrVO1Ke+FNBVjNWtBBL
iAPjt3gQkJK+e3WJgHGhHQP/O8bObwdF6RCDVV4L1spUhCWQ2cw+i/E2AMcSxTm0kZuw7MDMzCwc
fehRGzYuZE4yT0JgT5oi8sJ96Pd6apLewKnQg96eojga6TLJg+HpjkycWkRY9v4Gbyjh4ScfbNPq
iYCS2MaH45UGupHpaME1TprkO5JO7G06di8eYMbOyNA0Mok5ZpGUjJWbvS6461ZTwRYi+l85YfqB
RNNKErkGKQtTOw8CyPak/X8SVgMcSCC7ULLacIAXNEJs2QkgdyB24mnQw7rL1inmUN9l6wwSPysv
ZGK4O+uGC5/v/sC6+J3YNJ3v0fRyDm2sqD+eqCFD8p7urvNduz02R6O2diIyYJFK7lInREx5tFdB
p1bC2/mBgcLJkJRytGqvX97XWgZqlbJk6YehtYg85EMRK6QuPcXFY3ufNK/SYFVGdp7eaje19IC+
ZnmqoZlj7/94nFRz5zugFpZrhkhugc2a/fcnuChyVoSLq4ws9fbhwo2rshvbng/ONa9Dd8Zg7Def
Vkvc3m+/MAW91erDQSEPbOFW27NkgSo0o8pDYPpngTgVfThvxQFgFycoCY3XtvhiBh8Vm60d1kVo
lKDQ/UTmmE5XYrNsbgUQ3R3EahTZbMxTWyxmbyQFh439sMqyv5PpFDmV08Zc7FVr4lHh2v7xIAVo
F4A8X2YsRG+vrBYJuTEo+LORj8PiXO4FHA8haKemLUvXUJ1vRZaDFacP8YFCVFDPnVmxpT4cZ9Ss
nVb+TN+Dw5A7wznQ61b6pjfgkQfX7I4oOcfOfAdHFMiJMFaOxeA+JTDZ0CtrnKfBfuiPBHTU7C+0
Z7QS4+IRKk8FxVCVUdGZHV4CgKAe9n6sU+QzIBIxtZ4zdbDY0kkoGh+d4QshnpURIgE+uuBwakEx
vpWwogn6wUa+pZUAQYbWhfcM4RPdkMpSgcQhj2Fxvbc8dhzYfHGeyBfy4AwCSVnX+oIq37NP1GFT
f15R5jIi52oErjgDl9gLm5gN6b5fZG+zJ3g9RMh/j1I68S9o+GOaKtgtVhJxYGmzN5Ooew6M2tEo
QoldF8Z3X6Vzw6OiNx9lF5DRdews1RK36wF2QiDFwqydmW5lgfVsGhB8pzzJsvq4n+066ONNAz6r
wGOoXXHVdiB/Q0OY+enXlcA/MjptxlbdYQsB2n+PjKJ1A2V1xjGYh/Xn1J/c7GCIBo9K8pbAhQEh
G3qKM0SWNPLJLkiMWQfSx1XH7NF3y+vYR81HDRvWsUbrk6xbmXPtEjrELvu/n3zEdwH/0jPNXoqL
OxHseq5U34URqyVzaxfL/0L8E72Xgpr3BbXzzVLOV1zHEHwcwDoOLaBL3OKOYzLiezHcrdPUdqYv
xmtedvPFzS2HnS5OM/JUZVTfQ1Q3uBrE4jufs3FOPKgUR+/0EAohKIPRGROTtMC+goxOaj4Pho0o
rWTVYNCiY2cwv4137s3pjW5cOmi+7FI89cVWVMRMJG0QMah6ZgzuPX0pk6ZPPDzgFFbEURWxTwHD
rsochpQUrpSZz2V6oI5OaE4ssefU4q4EeReZJV7llXvThVjtUsK79Tn9jbB9QfhnFDWrwiBE1H3u
Ao4YV9R/Ot+R4fZy2GTi8TKLjTaQSE45oOFaKOWjrbjAUSFdNRXvXsHE2M5/8j0Y5Z5OcqZgkNQX
cWMr5uL32G5te3KEv0mERTVsesoZYzpxSom6Ys42Eijkv5MMrAjOLYVvPfYIyRmo7Afec26wQeKP
H3oBnetgmi52lcggSkItYhI3oRqM1JGR7+4x0Fh+6WI0IVPGNmMT/SM6KFSBrsUXlJsN8XqNgpKm
f9RaFHqWe7ZD07auoSH4+vlb6eKo871JGm/Zw1EKDB+RtUucOQ7A1AZjKazcgEpAFLwhQuul8KYy
W08KjgB/FV3Hom7FazZpoJWpdfW1+22f5ocL4z+T0TGXtMnuGZI0kHFKO+/tmvrArWlsrRbWXg4Y
qhfgYsSgpTaTad/0y8LlKGxNslPYU6PYf1Nrmgen5KAvmzb/YcMnx+U8prUp1qoyT3sM19V+yuKJ
6t3uEvnyzTn4GD64NqjZFCAHVSLXtMRbbtVMsjdAdEmqJI1kepKN9TVzbW+c2Y77FlGCxSMhvD6v
KixW3EoRnGmWDJ57k0Yh63YbHlKvGZqPrdmkAEa3ZQ2+AIqEm2aFGw4dPGa2KTwZe+IPl2dOClOg
Tp+IcC7XD4HrFtB0zPpWVOyjVCETgKKJA3w7IOZmPP90Pcnitqhl5cKoMgWH6WhQYYsIK7U+3jPo
ZhKhYC9Rl93fa5l/GBWMJ+76SXGh2t2cMTX9Z+/l6Gyh6l0W+21J0Do85+uswbrIx2XPMHsPYVwJ
su6cqGVFwjeFHaBwKreIx78Ht/iQezRPeKAWluUGGfZZBT5fVcJnrekVv2J9sNKqI+d5QB9QYA6L
kCpI6J/AQD/bT53+rMjxSJLVB8mnKuw7JorvaGHP4Km+cE2l9NPXNUsJmStlKK3FW4YPzdshnCSC
aVEaZ/V4fOsVwUBOu59n4SdlBGO2bZMCKBkfmI/cDrR3rh1mWeolgpSPlFverL0R/MbkPvjdIIcc
18eNS2tG15Ik5mK5m5E/YwOub5+dmjSIzlTk+53kxkWhOfiegTDXdZMj3y3EE5NftHYK2r1V5o9Z
uWeD7vuOhM5Z3CykzjZpoPJBbBR1IuCT2PyVzf0cAw0eK6Jsn8guO6qhp6Mhtxf/frPA3iKFgJ5N
MuHAVT92ZZw3mickZc+QK/hOMHcfT29R3V0XsPxRPfdYQ4M16Q7zpsfAX5KjGuzAAa//gejx0rcZ
Izxh7U+phfvigBUj/VdopyWoleC4TotoyouvJ/YLgbeD3AVqeNbiIe84BOaMbN/iqohLs85sOITk
P7OQAJgpz/bIujRJeA4Cyv5CUFBD5AcdsFLigdkOdk0g+ugu9mz0/GEO/USRyBm1QELT65eESOhd
0Nj6OHW8S5MpLvOz1rQAw9mvIHh+lbnwqwxG0ZvLkwgyj/qg2+u58HQt9/qpFIQcQoT21q/bmTK8
7b3J9YY7G/FN7TU+jXoeC9plCiEvuTZU+vIrnQU2MF/Q0a8WJoGmiZlYaajtsPSA+nxmRnv2ZgbF
TgGkwJb6Ua//Y8zwHXokWRMG+AyBq3Bkv0+xofYfuDxcHGGJUmt4uMfiF2UE10bHsuIeWcBovM/h
tsbpQVrLZRV38MB5tG3cP6mOFzzlxVsU6mGhF0K1XA25TvKDdEDu+Yjbp4Mk5lUcSaBHeMF2kOhb
OFQWn+zc24alHduc8eC2XDROpMBFxMIsaq3/Vm5iZ89mq9oY6y2MftCEAQoNQO1P1KoGENr8tXk1
FzHCvl7r3dUWZXV+Py23MC/ZhiIOinNp0Nz1dTc5+4xUUWn8KGCjY+NOXi2N4ZIOqBu8gW0rOa2t
JUGGh2Hr4i0qT6NoOgv4uwC+JaBSo5yiA/4klk0QcIOhn6muF4tCLXeMgv2DLllYwYP7kdFWGIHF
jn4qrrucBwFIaFZtsm0o1xoLsYmpNDy2y+RDIQ1MvoUI8NGyves27nin+udbOPwV6Dp5Ijx2hBPH
jRgCxRFpA1oxHwXpwbcAHDWoHPTT+HSC2uKaZxyAprE/9nviJcSaDiU5QDV6vNYAhSGqTSEUFzOE
0J0zsoucMQdkCFR87ZPadea01bK0s5mq3BPDIxxvMtfqaVwF+Z2DVBKmQKxl4h3/WE8QEMqIOsAK
KHl85qU1XILcwW5goOcGBh96HQ5hx7/1gpw9LVRZJLdftSiUgyuiP0TUDctlV7Uwvn1jwbw8u/i2
1npbbNS3P4xLcIAGuQQibxMcGUIZsUUB0m2YDqsAQviDpvtf60wbegecCSO1NJXXFTHILMJO7tkY
ywpwm9l9LZXdT6rLFOQPjFRUYAR3r2BmI311mfg2r2MlBcMGPWtrZYQdwnyCObjjJ9tocSC9Vz40
yaPEsmtcPnp9hyDADh4GdERnRuQP9WGGQeV+S3OzbbU1KI0AmRGMOOhx7xDShoA5zziTicLZY2yI
lic2hW1ZK4l/Asr5W/cVOQX4BQnwU2L93j5kDDlDY9PJxn0z4X68WRPavXq6DWqmKpu+pACfg75O
/pofJQwYFNTNviqdL57Y/710By4NRlJcgTTVO9Izu/LI4KvYPqHbxCKa1IrmInwnisPCfKhL2d0d
xTmAxeSUpJ6qByuDKmFzgRhWBRszQGRjOfw/5A3vp4LE2i7cFKwWVur1lrtKk4HVY9Z680cwo94k
4OQjSFO6SeZsp5Ty75ICrb0K7AGfpfXfKGsBhUbqCDUt0YMnk6WcCzW3qcR6Kx0SBgzlQzaFd9d/
TqSf1054QIzVMk6yC0HYj1Q4OV9n1pbxhruNWxz63ysqFCqPUhnihwvo8LjJjGsRzMNpH5LdZJTT
g4QSYxwFd4GIDqM9R69wD5H0Vqc+7d7Vprx1dy9PoP5zwgC8F2FSS6s85d8n+Ei1oFLwEiXexARc
BqDB0LqtxG3FKWCNZEx7igTfGcGM3OTSWuGkE/2n+cBkkvk/9xDDiFEH5z1h/mvnmlseYdoLgbtJ
zGX4Dp6y5CKUA5izFfXqpzK58Ryxs1UFNrE3PJNadhtFPx/noDmNOBuApNJliidgLloq0Ryt1yv6
oHvOlJh9VET6wFslXLAJqMkzlH7YxHnJ3xkUQ+Q0laE6vAOrVFLFjSvEZcSMdnkvgRwdmJfp5DgG
J9GDFgzTXmVfZCPlPzndOq7zZP4Q/aqbwrxeWFPEgU0168txEcFxt+m69d+uhyjLWaXLCpphDcNW
eml8FQlxoWDX6HTgH0se8QHsef5qAMVQksI3DOxYkcsfXBy3tfm70gRcqcD+wo48FgcXTTvXziT3
OznYjSijr4cxzQgFKJzuSMg15lNWRm6nCiiDG666XfEktGx56sOZXPiEmnpLAPRrqJseXcY/r7HJ
anXUmUXcDrY8yTYfEMUsZTzyPHF+XkO4/x7oRdrzeFa1MQlQ29XJLkYIa9mHCO0n3qfvt5JgNEGb
xOtdA9ZiQN99itKW8UkwyGfJ1c0b4lBAhUCRKB0qn2i3jpRsbV6fI1DWjRKj+5I9Z3rM8QY+tF2+
ApzXX2mhDpKhH+cZfTaPGIED84I52c8ymsDVwk3DhoGVV9co4onHJTR0QnmPgSfCLzSekYcFhjzQ
eeCg/CvLxZJ3I8sEihP4oqPkMpPYjZOu96KJiNphB4R4jXlx9A8XQnuzd6ZSgRjXdPeOmIJ03lpJ
HU9VQucEjZaa/VIAB9y1+32WsXOVZW1bi0Kq+xiDimlorT15aVpdf02FfEQUL4s09EGOhwEadK2u
dna/yzrJqUDA6FpZtxLt5wQXmbwmzX3G2286y2KSVKsBsSbTJcfBBsJwd3AQr2xCm31JctIEK2zu
2FV09zQeCQPL4o4gkot5CNwI9Dh7Rd9E55cseOK3awVILx6EzQLIZDHMoeDfTjjHLuYH+uJe4dez
HOMsdDJa+dwLL9AtXl4lsvtqCtn5VubWjcASYU2i10boL9vexzYpQfTrIwMLikD0SAJTKIERchxg
4Sv335ul3ZEEjXZQYNupyAMR2r6zL7igBalfp+P21fNyWpqHMriCsG6KFduflJk/VfQQY3HOfXtO
s2U6uCDnHzaq6bnVbXUisWzFsYDcnMFW4AA448qgRKfGxeStG0n9Ti64tHYB6AseykQK4UbtQ7jx
wJy8huflSBmlzs+1YsdjxF8yFw+Hf6ZUWpVSYx8XDMmvsTWhUACzFtE4MxoxPzCjsAbV/DGCqvcm
RTBokHIuzsaHg8pnbiTIiK7B31ZG5lsm64V197Yo7gUXSf0/ankGMFoC45bB8lP82zi63AWUorO3
fpH6dkznwpIplI+zfgyUgZUmE26JeRbPtNIDi4Sw+TIns7ZrGj/R/15cyzZSKWEpW1MvKT6s8crm
zR9hAMnYpNkfr5SOunNwMTUfbsNS2fCatF4xkU6/64QVs6u7CH/MDhVgZNtoXdfM1ixjgZqgnUqd
FjmUxiQqjx3Wi+BJUA7G4OQmk+NVhy45GfPUTJzSPcUTu5H3YGcyLogBego4USnF4iOkcqsQ6s6u
FWzV/r+myl+1Edk0Y8YYfOUQG8f1r2dPwHprseAFSPdR0n6zFhL5tI33u8qlPnvEnahVCM3VXvM1
NVusinBoBHxCC55DrjcldzWhGlKb+W6j7e1EQbnYa43+TWiT+wYzu4bn557l5Ja4SH7WNARxPPgM
YjdjFWAztbtU0llsOyskWPByE5YpvO/zuNtnMUkSsZmN1Nd8w31qIhBt0fx+3ml80OSeCjZrH8aS
ggLj6WeLXS+WSPnjEzYUEA+zr2OmXRcksiFA4u+goPXmdhGXYci67X/03MQoK50W8aGLVsRILOwH
MQ3QpRe5V8hkDLDmWzLVTqelIyUYInXjyw+uibXZh0R02Y2FA82RdFUgiv736M16B4kcQ6KQAPk5
VjVzcXET8/y40DiZOHz0zyT/EH45YezQy1BTOu3o/ufyXUZNePv9lpkbYzdCq+gA1STImolGHQAl
7Yai3lWEXISGCRqllOsRer/Kd3Ehkkb45YyWmu+T8We3V62HUnLKmRWjGVHt5iUSzj3HTfF/+cBg
/5p+XVCl3mRc23gVBcM7GhuF6PRwpvg+wHeHKJ5/hrCpU6rzUQNHQf/Euhp4j6LXrjzii7GWJ5Z6
ja2dRaFy/qVjVcMXixIm99Tk6pkObZnttbo5zw5WmGNW5M3x1i6BjU8lq1LRNeIlUtpM0BlDccqp
fJlfLqQJnRo4oPkv2z2zDGUyatfo7YZue040o5K5KBKewRj59V+vucfHp0TuIHdJKZgosVhjLH8/
HtY6ymelrJSiMDHN5W/o9mVPv9Qu4Uf4T1qZHE/Cm/sK3U19h7IipTCoN4MBliO6hopzqJX2XD5A
69SuhZRSFRcnLtqhI1bEr0HKp+/z5Dvyqc74urFzvIHlqn8wLYT9PzuVwvi9cddcucDM9WJsE7HD
X8MqkSokzSF8yrlXVOI3wc7dgbHk+O+rYuHJGYrBv4q46POQ8d2QLFby8QR2FKfKMB66oyCLyzCm
T/bUmhGmewdKufQUIRAIm56PaK6FRVjErmCGhIlljHs/gni+4B1aUteLMSHuNvE8Yxg3F0dz1pRP
9RaVMOr7yTV3ywAJ5vUI5kzQq2k70Qz/if/NiUW5fTBJIQXrGgmHTPePkPXIEChgfY98I+EApzRT
kA7P2W7JtFJTPMjL2XtUBVG5s0q9kodx93Hj04m16xGePdl7EkPXTnF0eZ370/N55jOFnQRllkfb
UWcSWGZGms8CjpslUltxkJMFsDQPJrTBRaiT610BZ8Ntzh7hSmlIn3eR93G+fpUOErKYxbGj3ur8
yt9ti2v7bxASxcaEqDizPx68IG5VFPBnlIaZcf0I3tvjDoFNwFC65d7utBuPwpNh4x11QpD8vTM2
C8rpFeqlPlw4Gv4niDG1mVuzB6rMJwazM5bnMdDMZh/fR4bn5Jw6lzIUyZYrQh9Fssqgfv63eaHD
MSw0VL21NglGta0lvNxXZzYNJuBRkJVsHqqE++Bd07xFN5NyTPNbKicnH49aeXN/38dv4pgiXfoW
16rD0tIpM7nDtvY7hjvvXltdgBfDCRpMNKMJQeEZswrvj3CphXnkm4gqL8ow2l1VCD2gC0Qxke4q
vL4wtV2dOS7LYHT4P4M/AdnqpjANyVcaYgpkBWqmsxs5sW+/P+nxToJtTxvCuST+tYFiWo3ntMJi
Vp7nSAvorX4YWUc5MPvQIuFvx+B0PRrQ0Q6kZnLyaGsWvcNLWTui+Uo9vbQqxVtOjXNK3/oH/9Yq
FnLVjoFk0qw/BvkePRsKZ6dEJxO9h/9oBqkDF545IGkKtms4C7KUjw29F1CbklvuUCU/TF8XNnuD
GHQNbLVNusELbGSRL4fuUvnrm/pMks4OtUrHZDz9HKNrUNrnyoNnMnkdounSfUEc84WF2IE5NSek
CnRHtts7O4Y0zhvq4nahUdHq8cWrnNunru5DGjOo1/chdoKtC574of8cEu4+4k70AbiBVDraTBK9
1eeB2BqQVyrMwUx7YZzClbfBe9BAk8+Geq/S0emStHLsDjuNYiUp3uap8hjAq/GOzb06C0ombHdd
V2WQ3/6vYznIju42sTL/zFzunBqFRfO9cjbDm6Usq4j36IFlczhOHGiT/lJ4V5UwjejFbACDVTxO
sJ0jk8B+ukuYJV7840GSIXFUhIT/x3AfwO/gnftVApy/RWXLIjSGzdbwCYj9IWnRsXS9gEXZ1C1z
Xfxin/aRqbC8gZqGnLXFEnSZ6jOXnXjZ9OYENdAK8sgu5jvQXup+Al1zCBBzWzzCZEZ2+IcSG1B/
JFhXw3ZBV7Z3wzYRIXGObbCZwprUYhiHquN4NbqKQQl7TPL0zkuAUSnRCzeesqEX4Bj3xYaFld0a
F8vreARfAGaIU/tGWVwEuSWyzI1ixzgr5uDSFnnt2M4lpN/1h4WPgaZav+AwXsvm8i/3bzJHliME
/5AXeuaLp2nQtzBkhcjjbrkjkWy67YP8FsD8QA1/J6wZtcG4lrmGVbSY/NUhNlQZLXBcnDI8nrv0
fg3fTOV8Z8i3/qVTt4UrDHigoIowBxkaLa21JWBOAmilJ/GNsXzq/EGQ/won4QfEIIJFX0KU+0Ja
WwtTPzY0Y8cWCadS0VY30ESKi+ex0DCB2PdqjBQgUa1dDOhVyyTcGjKL84tGGGeqD9BnGsDYt6Jx
4Ic3sJNN2KP94NMX7JSZURklfbgsenIUj98NSuGGDobdDPPQ8h1xRwxScSTHBTPiK1ApWAnBAShe
xipTAcj3PJh15lwBjLZNcjXlQn7WwRg0dQlnDwefJPx8O0PeUgQUwjQgEYA9CEXUtHpNyNwBn+CB
NXX9NCN+LSKU8/MpIkGzocZlsRQSZTaLnkulfmq0V5jr9D76g3G9BW6SHiyxJ2nelXjR8E75K5y1
NNgcN2uG8r3JEqwCiRmqmuOqbniUuUmDB5F5kHNb2D4gOyXPiKvWzkVcZeaAtppWdDWZgDtLV438
ljCSABbkx6wFgYzPjQfTbzIZSezWJ7HAbQBa63sUXn2FS1Y60iFXXv+oBf2BJgyWkwGlBF5hJkYu
IYPMzkYqQ1hoFHNnyVkm/i2cNv4CkyRWZiuWqU0IUDj+HdK5K2VHWTyIa1eaUVpUnGQTvmFpbOLa
yOAYbLzgYNqP0ziXube3xH9koiFN/K3nvwwYHjRBPwb65+z0fw2av7vEJeZxSFd8n+BOSqGTsNXN
4m3aLSKP2mrL+I/GnImlGrBfKDRrTByjOKC+RNeuXBPOga2YfN0IytQs7gWumx8S7Fp/HOr58ecM
KW+H0zo45Lt5QLP4bzluO0lZM9wpt5fkCLk0/gQD60mra+4EqKvgGREd2yjJ/KRM8J4mpYdoAjTq
j6rH83GZp8R5GUHqSFrZaY8rU5E59LLJudcrbMs+VfUIxRnzNmlvCWC9KEBg3eMgjz5AQqIoYgWt
OIoCJygwwTYhPhspOupOobCm1Oefnolz+IKaiFIuGcJh8R34kv2IPfzY9xUFSRBu1zvLPN2Ur8DL
3eDnqZ0tcJJoEL8SioonC4s33ubjJUjleObp/GDrSwWLd03BQmL0Mmtl7wmso29bpV7ZfaKBQifB
B3jGniiOS9et+uVijy0oV7Ba0lxCCMVrBj6cRy5KfHwlsn3gPwymgufLbkQnp7QPOpvHEe4iJCNb
1Ov5sGjv6H1GZM+oMQ38JM8ObYYj/yCFtr11IH+RSpAsh2RHvEVteDrp9mMcdjlOQYr2J/LmSiaY
b064/KII1ZZXKhkV1pzw0cR85MqNhGG6pG18L4JPDSf21xioCx8Fwp0tqMfOcWK8KCrlTHk1GlM9
ILKf+//IHrApe7wl1zNTmVFfjXqZUvWcYKKoY0MffD33ihpNA38T9CzR+IryCL0mGKNqno6H/EWJ
6qKJjTBjbICDOd55dHD9YRcQa0hgFu+VByUkul+cEmXbOMosH1f/75ysGGLLMo7191AX6B4kduky
rgkL3NcJIxrHIPgrgTX/QGgkUQzu08PmuKmsJhauuzZlWo3AltmOrbOj4WTUhQThx9mWjmnrcA3M
xBwS1lWzokGULbA52xB10qQMP5shvhgjnI/ohDboBFGdyRn24PfG4YoqAw2ebFfy75IB+PxRkSKJ
OaEPdhfyVS6h1UwNoQGlwf7aDetCxjWs4M/s8vDrFIaFA7pc0JbFtmShIYBhwjucZ+2Ze7LiC2EB
n4Phor8aqlOutmLm8SYA/Qel/HGkaUOImEOWL9YBRsnseIWEAWK/ggBxAQJyJjwHPFTBxf9ATC2B
QW1HRnQvRIzrpbFv+SsQtVaMi07Ywtf+FXLF3vDpYIEiZ8+/nN6zXpxlUpdKVRoIg/2zQX7VNTyu
jVTFxtEb0AduWiLNK0M/cW5TC/5IrTl2iSwzRxcfvVqgTyLIzGc2IO6xTXvTrCZBloBQw8/v9YCS
Drywn1QFnOJPSJiNE32CjO6JXxrT7GCe5xgjmvu7uww6vh6CQX0CTGAyTyE4GKqh9gpopi3EtLab
5gSt9g6srwbQirC+4dqMi14EY0p1z9io8bNfF7WhUuEozteWWnbwvz8tLoZLHxcnMDt0DUu2Hb5A
dJ7Rl9zNBHDQJC9TgH/xMsSJs8muj9xSHSzPvxbUGaYrt7MlLcbfQnZY3ZQXVWXQss7yzMpsoRuc
aF89N5nKACfPQ9lfJrkjZl6M1F9J6lJacf7qLr0PdDVqONZutKfv12NWeGe7mXCuMMMJT1jZ0tUo
s2MTinRPbJevUpJG4u8xcDsryYUtEBADW67wYC95tBuUIme8ThrMyCyNYRNQgAbGyiBpsr2t/isA
zXLVE5QCKXbFp3MwRdXI+fiiW0R7zQ8NQg9HJRvfWjyg1OFW9zp5kxScvYdih6n58K7mJFhg2kNV
fOpMR8YjBnlAeA2TO+J08ht2uuoGaNBATNBmeB89jRUP+8wvnvdnbm/mNYl2LRpa5Wrw58zt9SZw
9gSqwDwp2Ib+iNSZRjw5at9JRAXVUBFOhAaXFgLAQ1USY2FQuMdMura6e1YQZ2xi/HrbXQbuz3AI
RzE35zUDhdvFBZWdHmxw4OwuZc6cqldPYpsdfcT5zytqIYpJ+osPXRISRbaWRAB3Rjynfvo6a3K6
8qDR1C2asKnG/fqEnk7bBdmg/cLG9YzVwT+vgbdpheuZoo5oG0VIsVsk3o4e7hN/h2AeauGB89pw
Lh7Sb8asdIM0Cm49fIIxNvC3Brc2UC/pZiG5DstDsbxWqA6a3awf/oqqjHYapYrZHPIYovskvjjU
H0ZwAjxfGGspSmVTwDld0P8BBll8bh2wYIMFdw4pdhhFK2ioX1ApajVMOFQQRqvQyuBHJ+6qWUUZ
9MrciJzKHTaE9rmBDp6/u/ou14WstbRNEFiNNgiaIqoIBJccEMKfk3KCDakOKUHmVW5MyWgTZJsS
3EvJV/nVdN2KXHcPeD57qLwEH5qMspd0GuOy4fMoBer8kR7jTImDTgQ+Du803RFEAQ2LY5VmVMuf
3g9uQ+on/qB0epZlq6BxZ1FcI1FV+3g/fA5qc78sUAGEoVNa4Y1yV2Bkb/56CvE2WY7ILuGyC3Na
94+zK1ubTQOyDI8SDzy8LmoyARLbB5+U7KUfQt/x4SbpKDN2mXkZ32ovZaLbeMw5kcRRa+3ybNtM
ax6CqO3Exf51fNqpKL7wLy6B0Qy5+x217pNaRpsVc957a8mqggHML7Fpz5i5IjqTzhf1bY7Rvpgh
UXvBqIQLW97BF35brbmQJkiZ3sD6KsN1yiLCywUvg1stVY+cwMbFMtN45LgeJyUMdBh+oYQ/6RxO
CrswlFsjmoyA8e3jCZmbpcc/bWClL9uj++UPWMHjpPM7xQf/CGW4gKL0rwm1eyUBXFFC9gxR7mxm
Z/INnDIpmm6I7L4j+pwgLoFXH3BKdX/ibsp6b6puc4cMBV3cgLMW2WkdG2sqzNPMf52NKboadeLI
W2z2+UdllneNXJs+AyeMK/IyaCxXsYOfcmTTTHDjvdV3B+P04OjWqJ5yuRboYCha1UwAVNsXuMUM
+TKV6KyMGLZ8/Xzj8LkheTkGLi2J3p0l8WIH1J7pdBNMWLIqsKP3Npnsz0+XDAjkbwc9NUkq4I6i
LCU1I7EJ+qG0WIaRdxXXjg3HQwkA52hrevLWCTdrfOW9VlYZNNmDqhywbQN8rQ5Akq6XZWfGi0rl
zKKc9FAOBnsSF75EeVq2CEC5z4EenugMOAFHKYICQCx52wGYr/gO6JxuTWo6djYXXkQGAstrND3e
sbIdsvwM3uAWGI0aCd+hqdIbYkJNtffokuE7FoAopfgeHlrMcEeoOmNmWPKzSr5PAL5R/GgNiEbl
LJo/5usNPgHu1My67IRkBoUHoTv6WC8UCnBfilzt4UbyE2iuixB071dGFA5gbtdvq+dOVrXKpS/Z
spSKdGIn8UQHOWBayrtGJrebG5qR6tPSvo6kL0ddyZxvPx3pkgxgy/A0t7kGszyGJL1RWwzQW8Wq
LVBBErCxkiWTJGZmFcLnjZjGSgqZuIESf3FVfH7/FCaqx8FTIGe2ZGvFoD+otjk+Dt6Bjp18X97y
2+MTm6yQmqmMxd0JZUsH7kzisCPM6quRmx6Z7qEZXcyrNDF0fxXoPmMfqn9doijTXmYmNNRXpPFR
PpzeYLNio9J3qby9cRLreur3RJkWdYwhmt6sNPPp4UBC5Qy/5Ur0a53+YniqUgwNPqhGpKYeyYT/
AjpLf/8GKZH4KG47YbbtQf8+C+1MOt3qY3j0DZJEDS4LNPiluTDJLKKV1n4nJytLdTumJ14HDUF+
6384gAKjuU3VSojDXair/75pxIRbqkMH2FKM4cuZqCmLSYoDGdkrzRRND9b/6lyka8+vwApvwimm
EkeEWImJNaWNpQ0Fd+qguVjMKS+Iuw+zGFu60h9CciPscxN1byq+K7eI/PB6vq97C27jmSBKTT0E
4jCEZG4VSd1zX5pG58Xa5fF2GmpFti4lpz1UT9uTcD6ah8B56A8HyKKQDb4+reuX0yQtZIEQXdN2
nI8Hex8wll9KE9G4mgo7bv4vpzY92x2D17wUkmSGY4pECVonwH/IDxZpf/oqFpzjTVnjyQncSBPT
hPxsCGxUbxkS1QJHcVI8aS1zZHv3ZcS8+mtVFMbLbo7LDklSbmNw3WVw9VkyeSVA0sj8zQ28cuVK
R7KeRbdJhmLV0RJK1oVuKTtNwjtOzQfGbUxxEzonPRhulLemmhFW8eij9y60RYbwUbmZvbgeQSBm
xABKTfGYQVvcH9bRDgnYnPiVP+nrP0fFWtXih5nMmkFCHnHWcB+bODtBu3ncoGDm4a/NeVfHQ2Hq
1V4tUX4UNvuA0AIXbXQA3IVna422y3jDq7k/qOuHUYj6/WgxN7KKyh2XrblH3SRgcDPLDh9ToDQ8
5UuTEEZEMsfQhxm2K8lMh54UL7+COZBghmjQYt1UnvuVVoi0aPT56dEgYw0ZRycYalzl1h854VtZ
dnGog5eZbXMma/j7pPyzfCxXjOAOkLW0D8ivaA6pK2W8LmmQatbFmhWnYfnzEUqCOMIbAkgv6LDk
KSw5p0GbLbVdR61ni8gJpUPbpc90GPubtrfZExQz2YVkFbtn2n5Z/79VAv4uVmZG1PIm9ar4et0n
7Y37ufu9FLt0iwliDRbhcMgHdz1l1SElzGfEmzXiX5FQDtJ+Gl8ArB8OM8WA2j9lJ2ayhCGGn2d6
nVuTL9td6TrdsCHFkNTQrb1X2Yv+PxydOuGVzCAiJ9vSLxfF1xs/BZVZOwSNuTvdSLfut09sernD
VUEthHXJnSIaR5wmGYCQOo2/8Ih9i9vq3s4RbiM5JgGr/TDA3iXQb7v8OPuEtLPynqqWWgod/Xhd
0h981/0gX5UUcPG5nliMaDLgEoBxooaEyLRw9rd6w9RT6Tri5Dx9HrI8g/FGR3S7GsEtEDICZ8sj
dx3N+cg61YTqIb2pZEn1qSA0tQOZWJ5Sv/iZDTxq++0qVdnxGiY6muZOp5puZCZSu6c4Recd5SmD
CrLjbDo1iC+BSJUQSRdFY+PkfP7JS6nW6yyCX031VJSbCe3l8xxcVZORsJ79BX3aoWq1PRrAQPOJ
AIDA2PkkQ6TmrtAp7cGKP3OGXgEaf0Zerk1zgblEvHF52OGoa/xD+7ECkHZPUYQTOnnI9FQSgjQE
QMRik4HvgO7pjynPxz7t6/hife/SgXqH86KO1qMH6vwvrufRtrjbXdCp510T4qS7GnpVxjwDkgXb
ey+5jWOC2aSPa1Zzm6L/XKSXdJWRqbwh2LmglrStLTaqgBJAtY5vAcC/G2LorZzSK1qTYaQuAcPH
32vLU/Axj0fCdGtDG2kpktHyi9tpkScNeS4Vyeftd/MtT/gmTonFOS+75V7iAlI6lSRwTu6umd7z
IYer+ZkQAF+wTHpgbUEb7t2RY92lg1ShN4i/DTRUXe76tXkSo1jR9L/TenQNwGkHUn1XbV4wIrkj
GxrV8zYfBSD1nXijzG5wxzUo/JXxJhoI4UwZj1kcy+iydipFxaQe8pAbMwXQrvTxGAsvAC40atJN
EBoEaiQOtfTg96LUwmbYRGH14TSYEvFtdla/wgTU5hi3p2OMu0OiC2/dDoAZXbPoCRKQgSsPfjDl
J7j0FqYGTi1qhKnbJQMXXxD3+DdvujTz0q3njdE77x80UJ9pcTUrp0ni0yIjjm/vQmVEaYkA/kHd
1pIOElTmZwOfYiEoPYv7HW9VLzaQQDcC+qdWUyn0/jFZhDJv/AiIiRuFVCPH0+8f8tZgY00m3qP5
KvdhShLgpJNJsY3Bug8AtG6Zlffejr+rr+eY7GI0ijv1t1s4LNtiOn5jJtjYE9EKWkEUho60Yb4h
rNiv3aKGrj1hxCzOcF0iMHkTXTjohj9ikf2tD2LKbzidnnzqtXPY0oHyBI1fz4xXHI79r+Eb9wIx
GOAlucHyK37x6SZ43vQZaFIhiD/HhEIgXvONRtmw4LIIBrGJzSD2RpqZfe/sSG9CZ/3N1USjG+MB
Tldw+Xqk3Bm4+K6ie2tDcmYK5erPd4BhjrLcPzSIU+hWyWmEGBwLZRMmoFOQCUwvJRO7pKURnUML
KL75oRXP8bdEM94Kz1eaDbBOiaTUTR3quNTwcdVzP5+2sKPtytT0BJYe4XT5cOqAAQMgPd5UNqWo
loQ2BuO34qXJy+QHOWLCeHNkVAwiduqdyeDr59FfJknardwj5wB8at7j0sEmQ8ImdGoxnoH8A6tO
NzGiAqDCrLsOja3mZVc9L0LMJxWR1OBJw6FDwVCERSbgQYasXasFwdhtbzksQ1lflC6JtCl9teGz
C01VaC2PDG0nI1Ml2VwXNB858Y0i1o5wKOUk6r1jBWIgTfT0//STprBVlLxdL3RfYT/OUlkFrTHJ
cH1z8SlvhH1D9e7hLfpqM0xBcOs6C9jvVp8RWwXPILfVMM3tCx5UeoZeACsg/uZTIQ+feVqIcHBv
/e0DC8Fr0Ax2WWrEe8ldfR3uL0kA458AMBtgg1lxMiuMI8QW2csyXBY4pzFAQ0kTKofk0f/sppn7
HeCYcMXM08wSX0xzbFqKKLACoiQserFPbW9HnyRbwGbGDVN0lNpO2uWWowZmIHJP1XsSWsa63fG0
nPeoP7nGLG+hs3X6BxTrDUtHegC7dVzJr3Jumg/ao9l6f3FdskmL7khlMslePSVNXQzbYmCjEExP
20J9hHJt7nd7jSRo4gIZH2UMtofoN956i/4Penr3pVaz5yJbops2Q28O41Fi+9Er8LlL8NyQ5s/Z
IYmtPHpxL4kqyyftSslihYC3EPaB4gQbH1phJYVzZTnQ+keo1+8ja8bMt5edgvtw+k5tiFlaDxdJ
1EjzxT05O9443H42R40YnMZ1GKSvUtkU2jSoLFVKXdVNQED0yJOKtxMVQ8o8wGbQTwTN5Lz/eVcN
JLD4O4p6GhDM3uF47PgI3ir25A4eh3ZZduzsr3wBsqb+Z+La2ejHepf6Uj5zsAVwmBz75gPV8fAo
ndzyixgbcTih0//G8D/8BF/E0Loa3I/hahHLxtnc4TscfJSzRtVaHPLxa3DWsiJBham/IN8T9AqJ
fhwMGfMsw2t1UFd4nqauUzfoJaiDO+w7fXXANuI71DZHRL7FlOX+IqeV7j0GcM8qaRbY3a0tt4/8
lkbUGtXMcZANwhv4Ausaf2OWQgiCGRxbv6zTM89eGSp/531HZyw7bh+US/uyMFwhN9UKI5dg6bb6
8/CNZZ6zYroRfZvsMyEFgku5LXtkw+Br68Q/ZhbbmoC+7mrOqoeXJPuIv9vc5VyXrZFF2Sp2m4H5
KbjVAvQz1Nk/ErbAHDWIKBhGsgBuMuciXDXnfG9Lzgthq1D7djIEIaqzV46z1veAP8Dsw7QM6EgZ
UTq+SmNECEx2y+QgUf75ilFTTS/HC21SNnp/F64ty09JCdJ7xu9Voo0TfYRCvHOItxFp4vZEdTad
mLKfpKz98Bm24Obys+yQOZqy8i/sfc2sEZJzDbYyXzq4uw48qMT0rsGGthkwQyKsX6Y7C5X0qoW3
eduU8wzuzzBWvWsZXBGmCBs0AHhTRCbF8yydgSZSLccyjhC8Ty3qP4mjXUaYpXZKvkAWjgFbMzJm
9iGrKHRmO7rDhFNnt0piBRntRIYtGcnLtLIpTPSO+5fwY4mFMppnct/c43OWyy9NBAqF4O0+loKb
eXHnRm/c8J96z1novBelG6eAU5p3we83MFJhhhhKrVI6omq40bk10MNEkxhfnFcFT9ReK7vXIg3j
vLPX3Pe79rCTfhJKmAHH2zUdWHepLdVE9UqjLV/oDweDJiZdPJslbBxs6A8Pd0w61kLSfU7aumqt
Dd/TJyJ6GGWxizLqdu+ltcO9Z/ptkyC8eug1jq70nmVR7ryAhhi6yzq0D7NEWdTzzEf4A6vc0Owg
bVb6mQ3VgNnR/gsHM65I1tiUyZacNlDnSBo32XudiYMfLhRWLVynz6osTq5CSd9QyXmMdcMNqa8r
NWsM6vRLIuNU1SqFFx3TJ9/iLHiMiCZmc/HFAOM+Ex5mtVahnY5IAz473Dw9+xf/aOojY3dGPbki
/uw2hP9m6QLIw4ob4S44L2wh9bCJ+asOFac6sGuGJl0KZ02sYYmgOBdOFlhZ0FsTSWfuBNWQ2tEU
OD5HqoJbP9e/5A4tx8U9PD+kB7pN28n6rPGz+uAAhtiavKftPzJuM6e11eb17zty1OxeHb2uMWYN
Sf2ODi1sWP1UmjCaO2KipMhnlc1JrCEoEl2kStQwzUYEh44uuNrHR9RVCDK45ZMpMUc/3yWWbae+
VAftVSSWoAa2tTsSPtZWOSrIMq9B48dXDeK/9TFUS6axMOaKvw0VovzkhRQNpunav7cV8WjHUeVV
yBbVBlqx3v2L+8zGv7nhC0EpT3zEQdb8gVWzUIbgp22abUiC8aAJJT+NFK+0gx5zBjzJWwxqzWCG
oqytYCtrP91EMo2+h7jFoDN5jaUd6oQeXJAmzuNU0S99Q2x8GwPTiFuzrAbK5UPfBpUdFh9vnLP8
nwwH1mn2UnjS0PdtUjmWc1ZaLgvSlzdBlga+DG53Xf1JuewhIstSQ9wfK1U+MPQXQkvxVpws3+E0
ALHWd0JLALalELj4gtn3nI2X2zXyBNe5EO6Z4bKoUEnEv1B9HeCLYMQtB4kh2aMQqpQHU9Vy6iU3
Vaz9J6Xxc1lMTX/0BZ0T668eXS1+gnZOl5jzSYiOC/n83oTPy08lygnVZ7pOR9W6MNnuYk4ZwVEK
MOexM5Go6p9ojnZTGokJ9H9BZcQVhFOyTxEd5YB7Ux6vxDwyd+kYh4/6F50sZRHH6yeIjPKqB2/z
O1/Fa+TEKJeyxC9bYb3ZxG17PAhdsXZvxkMFQhhth7UkfW+ItYCkJ6iW2N6s8zW2iEuozpSyETfD
PWYlKRweJPTV4A6qSI2NoTLjOsCU2fV0iXBl4rdIX6OB9j9CKCTcek3mt+mhHBL4TQzwMQiXpIVR
CIqtnMG0ftLgOrDDczxDDcYmlCbHveKSGSnFI9yauHdluHx/JWlEcgxIqDj1sboX9OBVB8KMsaKx
fUsW7m2jDsVqMs/JbP2GhH/N/IUvmO9w/YrhI7CG8T95citoTNp6YbJQMUm16V7vijWVpJwtFcI7
+S3bnHUzFzQbT7GAqPuYn6XWaRy+tpU7lQ/AB82jmZxrn9i8MX/RbT5iCkrzNrEWxDhJsQqSgolj
fVyfz5eTnAlT4VNB8mnrvzMpUeeDNSlrSF/2Sz3Dm/DSHVqgr679/PleXtpPM2EH34Qw3LXwCq5f
C/g1CSHeu4HV4MwF27baZvTF7cPbT+BhecH2m82t6Lk34hgotnh4Sl9CSIDSIHTDiPBU1R8y121V
oOMnS6Ut+AUJjkbMeLF8uuBvGdZ1Y0qPVP/PXBC1JlfHQTVBeBp392WZHSf1V0zBbSxXba9TD1Po
fPcwPzEsn3RtUezmIgrp9SAFqspAnmEzMs2B0iqusIu5E+0P5vKBTBF+WCgMRcYXLJP/NIOISwhe
denR3OlYa1IT/DbArwcWXODh61LcY2+rvyIx9JV4Vv0YtgOtBuEdAPUg+QBK0K/ldH5/LUPbs3Ay
mNWwal7lg0h9Cl+RYgWvlZ89kx17yeq8nxze8T2rUP9B7268iwX/2QV/ZT6I596Cj3lKnaedfGRm
3R3DDjche+eLp8AwhvTi7K32g1XJ6FUWNYcu4JDHRzl0WCtzXomiY4bqnDe0fNra2SkEaAmDt2Bg
uiJNH10ZEjPclSmpi372ol9p4MBIlrexG6StzGPdy4w7JG9DQwCwE3+K0bZXPDyooES1gIGuEDXy
/wZWdrjGZWbKjrtJByH9lkg7k0viznHBZPLIkWcrrEI5ZfYaf9FI3uj5y6zOW6zUzlc24hwgBSWc
O4IDA2R6Z2ZnGEkeinqZoJqMWu12ddgjFqEK43lVwb2yOys7XK+oFwAOoz7jk9DRvH1MDOIPZkDj
skAVPp/7cCkDk9hCb4nBxkDxLwOVLw49I0YOJybjKeqjru0pVCFsQOzG6tbW8vwea5sVjrYH0WnM
Vsk7q00AaQHuDOQsEA1KDpk94QX3T7b0Tc44F5gVzlRjwmLu0VqXeezolWLRtRJM0FTF9jQxAxG6
u45dcx1MCxd3sgmobYo+e/S6A0VhjPy9rRp4FJmNUMMBhof2xA7xd/3Q38k+AY8Lv53x/Zz93Rvy
HOFVoekqLqMpqclyrxoxXtLVd7p37q8pX/7XxIgiyaqBGRPkst+syU5k+zQeujdMXDN2pJNBwYaf
ylXBNZolXa4GcgsRzGWRyOf6vV5s14RuVhqG0PX4Q1BzD/azD7FJUEdN0uDymTVWqP4npme+b5z9
zKM6mC8g4ORh9zQwHndH09qIh60awrkbn1O8MvhvPyj7fld3Pqdfr99N6G3FlLlHFjSyaMGhAPLA
TjXQu8UCcQOyfNZE5q2Qj4WJ/Qd3P1I9j9FY3gD7cZ4N/RGM+38JkW59cijTSChk6THE4CIhfcR/
8yzoWtvyT0yiSr2UGXreyjDtm1lQ2O1lZr8Yd/UsUWFywM8ZoBQ2qB49czAbQ7NbQ+ZHIi2TgkWR
c/Q2tqiTvmi0sbyC7dWEHonUQg20laSVt2EHBeiEgIwJjtAZNdig4E4OG4hNidAw+FCmHUZvliV3
uVLSBAJ48nzl5MNyG59nWa+QBvxlgin+N/XqZoAnwTH+lq1G8kxMRJDnJqislpchgugghOiZnaqT
a1ctOdToEbS4xZlN9apSp4BG4uiZqNZ4UoMx4v1ud4+ZA+BQvjmf5U7r79Ddl7ZgN7319IQfkriF
RH6IW5E1J2hRtox8Zet/Llo89bmEXUSXu6ZcGSXTPUfrTKd+CG1BdFCUz6GtOJlZZNAjENU3Bgxu
UUdHblFjCeveQ2q2s+9JdKcS/zvmlb1sP8jISVf9CILQjsE3tz8BMTl9QX+qAv2eUfeiI1Tb4gEZ
nGLF5n576XqCIELIzWa4RCVKI/ooDUItMwOVEk+SYZssEE6FJPSrie8mpc1h0Kz/eBALOAH/5twZ
IQMwr1q1zbkdUZe1UHaG3jUPHrJG3bnPBPXENZ+ei2hET99t7NZV1FSace6sErWUKmTi9TQMRBxp
Ph/oXoLkuPEsoa4QY5FvUpUxZpfK8dbUUNVre+vqhLajKBvszk4KLikoiwH5tYUK8oLRjoCzFLNF
0v2aK+wabNi1Y84gmxvVzmDmwJUSkGTASWmY3Io3AAFfEFKW9/o9HQJQSxI7Tiku+0+4IC28oIXQ
QcKdrfP1Zkd925TlzH9zR+Ioc1vBleUv8I6RmjQc6IBj2qLdq9KI95dGKSuTnwrUIe/5+aHjDQu4
dmzvJzaMyNnXOQCbu0+kXZg1jAsmWqrcRBoJD9OBKnyqNO9s3Sxxd6SYMVkmtJCkbs1bMEnuFuOb
4saoVKCdR+oQhzw0Lxq1cEGhVUZUhqs0j8Kgk7e5QdsFk9BQXiyndw398ggTgN7gBxHV1hUWFaED
gT5YKZR/MCKn76aoQ3DhWfQOO6bm4NWH9nxmOWBp/WHjDvvYuMSuMxKLaYxopzzZbr7aR/ILldkk
ujyDw4Vv2D6wc3TbciOzhRGB4gFxRPdrCFHOmdrvbFchqNpUNWrD1C3JdYPBnUa/MksVJ1mp3ugg
WhPvX8k74bLVnABKK/rtXw96lWDgLsnWT48kd0xaZVyw38BDsSL26prcGjMJsYDoY2LzYALZV7Mp
JdOOdBSivVpWSXqNgtWAlUXB9f9JLab2MQeq2q2/1iYsHY3xVtBBVhfjmhe+L+b6uZoie2xlI5nl
HSPc8E4U987b2Om9or0/Qp3Y4m9LRftH+SER3mimtkfvnL+NWD4wPcKBySWM8TC1IrUv97P/aYz7
rsf6kEfAY/j8AUj01Wa/FTT0648yaDZRbTBe9zSqffyhJICwrdT6RKrq/KU1+OYdwKfFhRc9FJmM
CrGFNCaNkhiBk8YqljVtYmKIZ3mj1TY83WDvnioKJZzvY1xMHYlE78CPkiHGtvgzN4s2OQGt/HHM
RkgyvAe6b9N/EDtm4BlelryI8AUexQcvXAf0pa/OcAdkEv9H+eg6HSCTcRI31NoUq3o93WGB/sRh
vPGSomWFLHPY62fd04KJvgdF0/iewCLjgyfxvXut7nTuRVxR6UpxrWalJgGaE0qYa0l005k5l+qJ
47h/P1pCz6nOAtpR1XarBOpqm08RyTnA5wPRBDp0c3igA0rh5jVIWNIIZyWO5LLwQgHRn6vbg7b5
XsrGxgG8hP1I/HurKxHsk/wvqIHVgHxCGPdQKh5iwMisblLe8JTzVB9I/Ld5+po7/UiSthNGCcPg
7zFsEJ6KCyXicIefV+HxkRyS3cVm2aAtcIMGhyyEW/qPV3Z1GXX0VgE2J4fIXyEY0ZafMkIF3nIZ
7H3vyH/uCgvR0lh/ESkezWj5OLf2QvS+42vvHk5lPVJWSwVQp0d+vpElCnA932tf6nVHGgeQvPVB
byiTjj8d7ROxE7vHJ5OZOC2/e7lkaxAVaWWMFSiIRIWLXcxH4hR472q0rb9n6R6PJAthom9bsLXr
d+h83F6Tzl5fA9jFjgY7QthsJmHfbrch6On7KlLSWm/s371tv5w3piAsLJ/TAyKnuMHR2PCYVVc+
eF3iffpYXhRpVixIifwXIsNUm0WuNGIaIyhV97Rblhf1FqjZxlZLe3ywvkcEJmuouwClD7dZUQgm
etG+BpzDylhma73CNaoOepP1K+Xj/dXP8qxycxwBEC8YiHySTwY830nGigQn5NCbMZ7muBHvPhd6
LSdSwyJBE/lLkwEV2A/IqnTzgOXQnV/s6V69aY/tRjke/yWBr4Pr4eqrfQnWVHxmlmZj9qYQ1kQ2
gUXWnAdBrTsAjVyNE4BtxRguqRFRGFIovTBlAVPjrRwfUvBYSQqfJ07gVhxi7hF9aegGqwPPH9Gv
Tw7HwwsrRH0BWro188jL4CqneILIZ6cmKcNQ0JacyUSrbtMH5cVYvb6kBfrjg4ecwrcfhwfl7Bhc
V1ndpU1HE48P26GoiIP0t+1lisHJnWogwE7R+lhZKzX0kRsigBqhRVoGjqh/kKg9kxR5gU5PKCNW
4+uKaHNNtKD80hhhi3UIvbFHzTur2uERTjJlCJ3RdB8vSLJChIHdUYUDdug1ZEey8vE0BwZI6VUI
Fd3WAp+oyjIcwEZ6sMtmbj23NIkhuezZ0aHLBfoTjQtk7bM85k/KbUGWn3SRt34b3z86jmtZuZpY
wcUud4gNJiflOY6pvs+8VQcnByBnF0UuhGGh+cTxbNGthmT7zXH4UIML5KwOk6C1Okxgh74pAZXK
2P0Y5HMNl7EsYl8NPiaxpulP6MxF5+JZfw9slOEn+A6sTv4g9tJ4bx69ysBZ/nMPMDfedGSWcmSX
FhAi9aJ+cAX9x/BW6puvQ7exlknoelq0tnH+StYCffA/BSVx15Cd2RYzWvFw4Gc0SeHV/5Bx1ASg
8cgIHuioozhTsbkKluTWAujPb3e9x9buFoQTXCj6b6/KdHhKQkyRwcf0KfJ8N1WisMqWFQf98I+8
H2NODC8yOVbCeuofPtGHHJ4RSYltXYi+OuzekxZKbmSkqnr+Gse4NKdBYx5BJxxMiBBv5lOsOqT6
j0S9doMqXRCaOHkSD4CI6v1gGu5Cz9AqNICKgoxRKdeVL/ZEif83griFVqvj0tTpB/XkJVqT2buf
Jim1zUvH/NFE3sQ3G1nIhzvdfaISc4QCGnQXpVAFpPsk+JW3MWXswbHfotDfy0E6rzO05G2sWGDg
t7XsM071H30PiltC6A7x6q8/0vLu7u77SL/LBz3q+HTXMw8olmtjUsK6zMTq/UEwOpzwq6NQXlro
F//Hqdu5sS2ryy0+8ByW4LHvdYSSPfDZfjtZ4Vmi/if6cP2ukO09+Ws7sNIzK4c9FWFNh2PEoSqf
uSLvtoi9sW/FtI55rXKlWIxnGYfIv/FABMMqzqkaz4dp0B0jfp474IDUZhTBGB1b4BQtEEF1Rkuv
L/aIIe3E9zFPqUP6tNp+EaE7Ys3TwxQoSzRiXjYadz1BenzjFPnhq51XuMx5pTyXYpzO2zKreqnF
fpldFKAiK/PQzwkC7RHDauIFYWCzXJuY6EMxqpXw8XVPKwmqJMMgy1IKYnmY7HoEwtC/dBL0qyDC
ndM0ryEx1cKUs7+L8lQPlrwW1dVyVhEvYu21rQLEcVN7eVzRbsYaMVTiescCM+0KVs2lJbbMZHiJ
zAdN5ARlu7Ti5wJGtP5QzejECYoQqpUekOQ5vCrEVx7fsrUo1TpnDL9ToT1OOLz8/ntyrpPt2x0N
umTB2IWimLvvbN8ccuQrw+RIRpChZZLQ0eD+UWT3RNV/ztl+GuaCSS4bpGlzaZEnM+zirlYNlz17
g+pOT5/BfjqrY5UMDA4m0RBdX2hEdhZ6zfFCh9zo/q0nGb5zQU8JBXMg4avqGLM0NI4Udiyxq2z/
713vsdJAwywLMhS5/V1Ul/g6WXJQ2r0f2NSw4iJb2jMTLMfZEEHOi0QFi+WCr3p4ePAlaKAwx+Q2
aDBVXiydQRFBBTvi/ItIzDp9gnPwVLVJl5ROt5NZLcT+3K+ISk0/ODXLf87gUnRS6Qdjr22ronRC
+HffOu6vx6uY1wUtVwl0SP2eUDQkekfWcfUnFzNNMTg4u1K5vIkeOyThmfANyCNpiIEmkif0yAoZ
AZOMdxQ+fFDDg8qUpjiX2tPp3GxCNnrq3A2qkFOwWOZzxowINlUg4O7AfJec47WTo5Ic8ueND7Tl
45FXLqSJbKnqLO2JR9oTHIuv4mOPdPD4/FxqCwsEBNmAfjKSLksU5qvj334DJ/l8QXBrLEhHRfQa
0WQEMICb6Ht58wymRm6jvKJyptNoulRYQLfUVkQWzFQ/TJ+Cz7oMoFcIZ7BWKn6VyXsVnT8+vVew
FTTo9Psk58wrND27KJGpW/vQXRvV4LDe60xI7ZSGH9d+bpsA28P3wDnAIHm8z5Z8u7RPu7PLxz9K
THx7cvNG9X5LUcH8EpJn0hSneKNT0/5pZGzup+P2Iz9B/CiY/OlAHCG+PpgeNiTdIKQmYnPHatgF
/z0MEwiaxmZO11szqJK7u1YMqhQ2xGKpFG+Y1J1EFYLXfo+fKZtMDJnlPKsAORuvaN4atNg6L8Q1
U+f+VCvkWy56WXZkU+NQPl20J7SnI70WZGi8t1pwOFBkZN25tEb5JGsfvm7aALQxHTLIVAve5l5s
/4KGTMW9rUmmLefmYcscbhy1N4fk10a4wWLzQQ62KBPomiBSpQ1k0W/9/hJ8kjIijk2o2CdY0ll0
u8h9Me6MnUFz1+KxY8GvV3kdD+4IZjkJe0ysW3hH10uhYCqnwTKbtgSIMOvCrh304bwF27ECHFhn
sRIOwkhiNULsMrzyHuGgHZ3rfafjpG6fK3TIzTdRXZ5dGBJNUtgfxQHHEoZI4VX9plgbx6UIyE1m
zFY1B/o75C1jM5ucUZzTdDhBLzSDTVsD6jkzqwV49I8YYNFcLz/Z7sBN8k7AItIZMCciHDVCXSs6
PwTRLF3qDJANCF7ECP0/g3/slZvCF3Z02o3CSNob3gZ70YVbtIZQ6EvC3o5hLxMWm1Lfoj5AoNEo
qaqh31DjUcyiU8wHureKKkcJTjqcaZBmknk5KEg1BvHzGPpZ7tCeXH/+fBEqoqYvNPoqvE/AK4hO
pJ8ubLCuo8Wjze5EhGPs96jsZIgeZK1SED1oB8zVJRhVgYs0Hq6uGDsL+N/PykkXn8I0Wr5Al9dw
17gVH2Oks+6Wxxlxpvdw3EAq0V0uY6lv9soDukgCnnRp5clpAUPVGAjuwraNM5xri8hRXtENLbGV
qTfhhzN0RP1HgmfMwh5WKgJebMdypIeyfYPi5jWa5232/6CA1a5kJKBiHY5uiiQzj8+lXntnk80k
vuscyCwxlDByZx92phtfUCF6xdlP0P8xUs/8zSmv1PH2tySsBSVhJXh8fFOiP8NfJ5zpUKsGK2Z7
pLygcV6gayG4SQIAcI1np4XjS/15o7FCD+M8hjZg0f4f+Zs5qFZpu1TsmwFJv7MmzWZaQptvAJXj
JGMaYOOy8yA9XMdLOGbs3QkLaBWOmxyExoOc1Yn4ee/Nli9yZyiukozXfzTyzCmKDT4/c6N27UCq
GSROk9KyyemVsv9ADzkWnDgT03qOHwQZboWu5Qx5GbnsVp47Vo5c1aNPNMJ6PYUUI0cyaoANDNZ2
jdFjg7roVdaI651OSQ8s6yxcqX5fMIVBUOkBvv0b5RJHcMxOEHzM3zgg/l1L34Vo7dWBbOnXM1b4
CYi//IKd3Ms4fKZ5IooktjWYLCN6B8OYTxwuvaK14rFZfxgPM7PP6nRiVHLObCTe8yC+wFqRoKIJ
bl9amRi7zIxvv1/Ob5LiBYPvcQMTIa5yj4sAaLZCtc1BSMZ2/JvDKMqemHzOobKOUWhI5RMV5UwI
a6a4Lni8bkjf8ghg6cuYEsIUQhBoHLjEJ/8Jh5SRP1p9hEQJQ1kXzXdzvlw3lovc5O+kVB2hkRYD
IntQGZ/pwS28ffi4TassrFzUy3Eg7vb26ZnJLMvvct1ZhrBugjI8hs0UpzaPOwvKjdPrgNjKz66c
Oc6MeN/TkA/CI8ERb+c0A05dH4kdknyLp0YulxA4ibNMd8Vm4nXfhXWa7iSnkzorTjqlVVJSn5Em
QhdfWaDwdnnE/vxZW/AOr6lf3Z8hed0+DkyUFyGRMZ0sasiI9LaFeiCFbiDnWZaCqIoaLYFd117B
kZKXwLqwDS39cz+tUaKRS+mrZzg9iAHsr74UWg4S0OlEgFIwqea0dUZKd73oedBxhTQLpILD6wtm
KZagrHW3if5AeC29f6kN6em4UQdPbrgy/biq59fiTkY5/yzmicigUbzNbwta20fYu+y1v2usvsIG
nAP7LYz9+jozvl/NLTl6GROztGCH6NiOrePYSIlg6Kpd4T7+Rnw7ubvrdm4JnLG8ereSgXxCD6pN
4u4OrCKqsdk5KQBk4D7iIGmF66hxixqKeO4OebzSNlO5q3FLc407xHB2oODEczjNZ5F3lVTiV3Wb
CVqn7/rCo7MjObFzoGYm81h8/Md31W4maxWYy3BIcCTmHxzfPw4JMT9UMO5aFcyie/zmkAYrgET7
Z3DjYuQGS4y5kI14+eY2510CX6qYJKn1lv8vObiHbF9PDhya17XTCXH9CDCeBP/ZBFagybj3pcJ8
taTcvqsmOU0mDZmJysTSPj/zhFi3NnphPmE+Fwq7hZ4c5ORDxZt6lO/his4SrJV93Jg3brzHEvku
pXR5zkRuISHSLLezZakMueja1yEMIfHFjbzzmfLLQv+kcuctbCpnUEQKuTG/mKGz+8vvNkmfRH6l
ILUxFgpj8/6Tne+cvD0XFo1dJC7qqSbUncw2TIeoNr/BhcLk024k8k8qUBvTMwo0fm9BkhboB1Oo
KlooAes7ewWb9GOZ6+zIyzyV5yfZVKN/H++K7nXVx2O6c3w+/rfL0I4m8LZooiqP04c8COxihEl2
m1uDeER3TzHVnjS8jLb1cDurYW4q1HWw0HhoYj578s3KpwrVsf9zJutOmS1OAMCtpHPoAB1uo+n/
T6Qk4OtUKj7IJITsyr1ts2ArCtD5VhNYPlQjIlqt+npZG24vlwwePIjbf2Ck06iB1C7EC1D21bLN
KSnYVZSoViYh7BJ3tbhVsAVM1tkVE7vh3O5Z6VNev9pf1ilE+sxWVPIXhMzXCl1xPhB799f2qXql
5t4Xn5XLcnS48ldsXcqCaGN1DF9nRspHjL2/ymhQ+R1jQSIWHmbw9TG2xrd01xIKnuUgXOZKSj2V
anDANR5NAsV420fe+L1y5aSzPT589x9BrOdNcr09Nj5FdOXWtHK3GKHuRaCrGeap+JR98vrmRgqu
kqCc5/yBs01/a6arw9YH1LzKMymJJWjUsaBhq1vF0YkLsSMpSohaTSbXJegjLWxwIDaUlgmj4hxc
JmXiwFdHj4TTTSxLF5IT29Wu3kunVFukQwtfff7e0ZFkAw+Wtboxl8Fhv9T281I1jFrYeFvLGO3j
mT09a6NmJ2fsxbpWf2TuQV65d0dCqhdvKGRpVG0Lmp2r5BOLof0w2+DbV8husH8KDRMUKVU7WcaM
h6fSomLvNdvq2j8bD1vDj7ukCxzM1KeoHiX7Y4KiX5mis+nEEuflHM/W4cTACNwXXzy1Issyr5Q4
OGAII1Pqok8Lfx4aAc/3MmcXSgqip9GsQH7xMy+5YnEDHXe0Ij8sKKGmh0+vNskvkc1G+rveBnwx
9Cfs+Gr2keXVPCpoXre0nfrsvhWkC/8i6jxBcV/QNVtfHZKKLhIhFSElNdPi0EzG9p2Agsgjrokj
jaVybr8b7CRqZSKkQ8UG7tbwJ0+xjqat5KJ1aoZv7tzCrng1ecONiZphlyXlTIAfS9Vvcz1HJ29q
qe28SjCT5YzDFldqqsXUhJP/YmEVR5d+oPbCecuQVVW8Z+0ffWwS3bc12KBGhNz3fIwKuOxkBRZc
yLqvHNccWpbu9iDPyO3NQXnkfGAjUnomQOzlOoPdohjbnkr77TvJwMc0Z67xT6kMPjjEK9MCygEy
dnubH83bmQN2b30pSD2VmV/MyysCtAAnsFjLGfNgy6529ESp8zleKnO5/bbHbR/y+UKkxUaL5y36
XDxp83R/Dq7BksUVD0xawkNEJojiCo18Cei2rmA0z9jIgMXc2sk8NjmcuwPrFBioZG2oFdEy89tM
dP2WfmEHwQgCNvB+lmxDpUF7xewFBh6d0cN6uyyd9Wl7j8sYzoJ91GU4kcZw3Gci7pPGq0i9NGtl
dHjlCffiej40KGtWbXBhx1cGEANpw0eI33cMMEvN4BarAwL6Plm7YV9IvTXCB59QiRj4zXpVF2Jj
2dFaxVDXQnBQ9GPtfRGDfyWtxbxmeGqOzZT74BsjP4SX+EBddZRU8ReztK/Gb9owqZDCn6Yf8n3N
66sTlbVZtgluHFuY4wOCT58F0NKpEzW+NltnCQ5qrSw+1XcnY8UfvFtbf0GPguwnGfPJGSbg1upg
9D0ifsZzxHilt1ItAU++5YSEvDLgTnDN83NzQ3C1vuRyYfOe4ClSq4hWo80g0SS91swnyY5LFqqi
a6jgHUMwyrBbM5ZrEe57Cm/2atsJIth9u5esAeYyAhYge4q6PvMZwZaN6L6qLqcx12t639mIJN1G
F8jRcKqUzYpyB56TpyV3Mst81IrtjIQxvYpMaXT20bFd3DJQWKjVyjAm1G/HIY+kBaoe+BCUIfeN
7P02RiSs15Ye8Je4OsIRtktZda1zT/vGa6W943piJ7x3zePUxN7+g7TlDB7xHzXReKYyny5twMpm
WSQM19iJyK8H6xoFBO347/uQqJQp5CuZ35NypLik9+l3Eg5DF9gfZueyUyTQaYIzQek58G27+qV0
zWyHL8qifUkjGgTyOkIZ/xZ/ytt6lEk2YvD6lULMcPLGQJDSduTFyk/SBFYIuDAu19qN4WKC0WZq
EvDrCgZ3KaHQbwEKxiq0WPsqyzkuyzfveh7YQZF3vLnPgt/uXChWvKg98fUyxRhQ7+AfXRmZ8Niw
ZpBBrfFCFyzyelzI++oxl0VEpS5tA1V18qdy5uc+fs01c8TtWeyqCB4Y+eU2ogAg4rkpXejGjFlS
XMe1wDbGQ+i13+X2WIn3gVCuzcuHCeP66EUHy3unTEXJBncaVygLu0mejJlvTwuQbreL/XhwDOl2
8PfOne5FchmtPHaVqUAz0IbE1PqRCrZ863loUjXNAvI1zHPi9Cu3Lne3+wHTjeHxe2K01eVjl7uc
bc57IfNYsgU/YXmE64nPFDvjZ70J1EGxRyX4mB1P8xjVkWjZh25gbg1I1VQlCTxVTB+X0bE2CaKy
R2v9BQ72In6XckevI2kzpkzW3Ey07BwU+txxVQwURDQnlilOXNVzU94g/v/qfE1QNJxDCz53+6hN
UijZm3Wi7XHiCvX1+Wp3GDYTiVcP4Qppa5aCnrLn6nKwSt1E9IWxJsMdwoRwkPNrjgrajAK3uw/L
PjaIhGoMcqTTKmdOzXVLP7ljnnbD05++P7K0zt3TRdhVw1N8PcmsUy8NkKcTpcQgpfY2eKAvE16X
abCmhWR//yot2Xpk/N19WphEczTPZllrpehY9rWoS8+yUnoKrG/zCi4fvXwHOCxqsbNHXGyZBrWm
XnIripR0P0t4zTjgS7Rr4+K+gKKXWRAqRq3rIuo4FHGMi2YAoRLsicNYztAxt4tr/IVySiHO3IR8
/WHpf/CXmq6wSREmEhaVOG36SQSCH8uXuciXUhJWM5u5KrrwTO3CH3x9Fngegb38hyNdWm+Wi6ry
qvYsAub3WMzMbDTfq4y/uZy4pH9MsqyL20LP+MJx4/Z1xeEvI/ib25Jhobf6yZDXQ8YutYuXz9GJ
JMGDOYk0LembxLP46LcV46q9S4LY/F6gjh2l0Dbwm2kQpVVbZbObbbVDjwAucLB3fGXJVrpywZfh
vIwWXnk1kSRKWYrH/yhccByXoJXnEqX+YzmWXgtbEOLcuuA+QcIIoTcsef208hIUetEtSE31/pOj
Pl71jEC57+qd4Kn/fOrMioLKMYYKxiHZJlGVD/MXQAx0MLjYewfytRImFNa5TUqCS0cFaeNZfatH
lQy9vNr8i+JE9zgxmTehTEAjdxzVy4EDF8MC0YV7XrNfnJ5WaoddgfRfJ6b7njMq7caiUpg91XHf
5UrC/SSBA0e13/bHAl3FhktDAIC322rSXV0yFkWag8FQjnktechq6rXpkiwTR3X8h88Qd63DXftH
e2IHXc7UEeCsdiUmxBVdhPzt1eTNfj5aA8i2vfJ23taVxppINpk83wMTHYTt0RPF55W/yTPbNsM/
BLyamGcVQRdgTJZu9zF/s3SEm7DNS7TZPtrfg2gg74fQED2lUleDj3StzvMK9Tmk/tOe9VViD3Zz
+jUbnULSTcdfeNuNBoL5cL59na91VAqhJ0tYPAgSkmce7FYreeYJp94cKrKa/tVPW+nuNWRLoTpo
KX+WxOTpJkJHsV+PFbmlZj5bzryWPS7HsmX7keVd156Nzqb77JfxsLNf2I44H421/EtkDWoiwlFU
TwMAhMCHw/cHbv6//1sYcangOpwDRkYACE4P/FXixzm0Qcq3UAuz2mW0dAiRPpVfBtfrdZM/QGQ7
GKkAEHDZJmWkCPF/UWahmUh7m9IoeoP7f+t+0VgtNFClslZ+IN2kY+H8X41WOjcJuS3qcfmBqLfz
APOhkMBC8WZ/RdMQ5uqKMKcoWHGxReUOa52N/j4gJajarZlQLVq2mQjSk/XKN8BOxc/5iqVQQWdL
jjq/8/TpYa4Dy9+ebdpDQzEPDYh8wC2BVHgFDbEHEEcoAyczDLU3Ag00kKja7HZEc3meYeAn85yG
bE0NeiL8IyzviD0qFY2Bb59UCxBvxNiH8DV77tBVlukBGOX/N3Oyt3qZfttiApLCUxXyIGE5Wnmn
s+NtnriGhNPN/8Oc4UnROX3TrtaC62fQF1K/pJnMoEETIURMUYrFj5soOQq4AWISyBsW9Rz8AOtZ
oOLnEcCUO2bDamb/pabjHxxfP2NWx/QWzJCoOLeYpKoCgl8vFerFLeeCNteIlHm8qIG5okC4vPR5
JSSYoJKHgROI5PdcZxYxpf4Iw8khvgdlJi5ngsA/4zAbC+BT3I6Us52uEIrQDB8gKhiACbr0I9Jy
hoXWwu7mcIPLJpuqW7daKIoydBOVQFOb5XDOgIgtsjTswWtuXShO7jXwceFmlogGe8HSpJMBdsRJ
dubG9+q7c1AwGGOgWR42X5r8jPvD2ess/ibnV3GSD8GOSuQgIBrUjoFiGzj3vXMnbxDgV6lJ2JFJ
Gi9SE/NXhP555Z+b2upHdv3ylTSqtnrKnS31p8843eRAy2uweSImeDMbnLyGFjujeU5WNwZgYXtn
yackr0ZxpUnJ2/VJWppvPWGGV+aJ0vjeLm2dBEKNVrlXUGTmwMVHb7uKNC0744WIuqtC4/a0FWWs
1AeP3gI2V9KtAPYoXEF9UINma3YHAfU8M5ki4/sp3LJ6GQ0oAH7cAMr260LNI3KOks6i/gS0L0VQ
PRuqb7ufnLtbC9JyV8IZY4nP6CnJ2NlhmjQUAeRoImsnzPqydgIrxU44wSGjffffHi56tKdGNhNh
vklOQoB+aBx6O2eb3vJ39KU9x75/eETOSeXb85gmlZxB3e2OCrCZthEsBIbFMp+QgwJ4aByZS21p
GqCdaoS/BtJ1oimDpVgw4/dAswQBs9ddMZ8M65X+G4F5tSX11ruBDvNN1w/VXRCgz6dzVCRq9q3F
rQUvE3h9+xNKrxsMrnsyiwBKnJz9G7kdHAB74Xr5Vj2wsHlPMcZkGQNq9fhfoobE/i7kRZSd8+TJ
4i+0sThN7A/jHVUqwI7iCoeLuT2ksrWlmqUJsDYjaEE9BGKgSNw/ZZ6yRSQPijp/SqgdT9V7cusV
Q23uDSjYabxGLPGvhyQ+1g8fTokATKabeZ6kJVUNheIWWnsaNn6k0menxltKGvbb95nhpOv++sTr
G8Mv4pbyglhUVH81tsplnH/nUrha0XWH1tdk8r9/e6clvtIpLcZx9neRVe2jHB2KTa4QCFr4Hsg6
QzHQkOmgbj802dKDHz6bDCGd3xLjXz9fDYVSpghqmFkR3gh0llPY1pybJb9MP+FITxfFKhzb+2LP
EBPGfatqO6KFkPAm2ITVeiPCx73oE8HTL2JZ4IgQ8qE+CY/oGn2ts6TSCOed70IuyEyu2hp5bDCi
8nwkuIKyexQOIJr7p1dz42B1q5nAhvhQ9va/jAjiloBOScos3rYDU7BimNOzq93j/NRR9EJZnhOg
6E+VLBJ1CqYWTRkWhURLubYONdjeROwE2rpVyTxJXOegrE2xAHRN+ZXTN9GRBUJMSmVJiRnie5DM
2WdRsmBonjWrSu0JwHPJX2DbhnfK8ev2lONmVEd9dSujoLRckHQ0exLpxx98uPtEyQWZyIhb5tYq
ut2+r7PgEQhJK5ADTMw5Zhaj6T4TAprlLRsCqEp7GWPegRMV8l5kBpggbhrL8+xW6K8U+y3ULMrF
+w3eh6LxlfPg2Xxmmz8rtnosQkrWUor4Zo6c+3uUF5QZCGudI9QUa4H0ZPQbZL7LDLtZWvMtf3uj
oMmH+o8kRzEADGTT5xQXNx7GpXltcIizFTEGUY9nqn/7lDfBfE/zakcplQu/epWm5dMxqZ8Mljj+
e173B577IGe1vzKezmK8KcTPdKQi7kAA1NnB01bKWVtbjPwVR54OB9FpwluU83rKdE5XCtu8isoP
6yYwhna4mt0BBH+RMqDcRYmEg/cYnIhPXulrfJyiJ7l7Dkg+5zN11E2pBB2jwVdOJUjuwYtUYL6Q
SBxvxAhQTohddAQBrb75/j9Asm2yPdx6JglNQPgEI+ra5oclZNw705z/mnohwNSE14lr2eDQqL6O
EQjlO+lSyxu7KyCNf0O+9lu1tA/6/fgOvNpZGRzUd9v6TySurN1CzO41Y9lJzUOlTSt13RHskfDk
45BTTw3WJae7+xRuG9EI9VvUK6/XSqEZQqVJ6VhNC61U7mSQIRbDtNzFwTaptXR0fm9e62kzowvo
iIyDWztAaMNGtAomp3QGPB/huM3Yp1NLLyWVopoV2Jza/cVNiwqPHLbHuqnfCEnwDPQiRBS5YXkQ
QdIjlfPWwdcDll+JEBWcf93Hif7cRwQvkydE2P2VPpzRsHNUsxlxRl3dpkoBTUoyGzasWSTALrSN
+nq/c6BypyPqHf8wHjPq9A09fbGGVjliE2kH+hZa+V6ntMcLrtFuxPUXy5M/gOvIB9fqDQ6G7i3M
2aLLl4KVPIHOMdyKJYpIPJ4mU1YM3/b30puIJu6pt0SsES977TlglwwrBMlZh0XnUEAblq2fVLer
1/+Qpcd8wTaRx6xp/eZ8sz/LhyzXZbFkYSWQz//XHUxXv5Z8qE1ktjaG2bia6y3KMl+Eim/pylEv
41ukPF5h50JOyuqjMHbAJel/H9mNT0TdHicw/WVKNOSbJs72Ps+uiIAJyeCbJHbBM5A12Y38/CWE
w/KjeZ4bSOPhK2YpRSr9Par03LzwG1/XFQwFDOFn0Ka0eQrwo8z2z0tbgV3Va3m6IyhrgJnB5Dbw
uf0KtJ35Pa3DKm2AkvmY8YS66pRKZ591rkqOWz9iNxmwr4FOBGCsARmr4PcVj0sqJmt84KPMHgm5
14PXDrlIH9N8WUJ4RWtZz1YbcCOEbDgbzffv4UNIZuQUkwFL5uywY+cvwA9t/BSeDj5VeFDOduYo
/DuGFgN6OlbPC+iXWlJIDRbzZuO1wLaUyMsk+lU9PsWHp+xPMGCq4PGA2Az+Oee1N5VfpqQ2iIY/
v1Ruo8B1qshcsYXVtnv1QcqqhYxiqPpNSVao45SaFnSxzZF5cH983YNv6ZhdxgCaIsUFZbouLclo
Q54f/ICc5VnJ/kxOgRzjF2IqoWj9bWoxbYEJLmYyeMrSoO9rdU7OdxHuzcqLCZ2Szq9tk9eH7ZFC
qLscAPO/iig9O5E55aI45K5EWZodrLg915egR6EWzdeX6zJ+i9OHKKWSaAiksleO7xA6FJmNz+8F
xrkAVo9ubwL6UOYj6agTJdL3LHT6HxDwPKvsOQU6alSU9WjC4FlaGLqYOp8HW0Syn3MyFlA6mjVs
h4gTD9dmCrYvwL1XxDVilKb0i0czRpgWPOpsW3ULMhqtGqpFFWhOY20ruynIc60IFR1E/Jru85Oq
01wko1ViaoPog9Zn2IWasJFNIXj37L7U6tyIEH0doVt6zS+AtrjCHhIa8190FHlOQOWa3Qdsz3rx
ZAIvZZRehX4Cx5ZnfNkVIqterrcNw8t9xhjC1lwKOOyUEX+OzZv3ruiaTwe3Ht2GovwFE2CHU5PF
K0QNbaGHnLqeHNRoeCpBZhWXkDw2OtM0uErcymy4tY7xBANJetYN8Thrw4FnZYj0bVoqp51BlcTd
6hFyAcclFfW6Y82ZFcYyesGUJUkWXIv+KtyYBBvIxWSY4KfRocrhibZEyz6wKI3UdkaAKDI60KwN
tJrYSHaniN/U3K22hPDNjFwG0aWNdKyiTjVXLpsEcA1W7xkDkeSY8MrzLjuFlO7xxXPwedxO28Vr
uGf2LU/UwbwlvSfN9TF8o8eT9gXcoBSIEqvxvOsfS5NcbdPfEAUNTodWh88lWJUk2XIbXJEfBN3j
0jUvzP+ce3mSA8PJHM5ICpJSvzGo9V7grdRYa1O3kfNXt2sezOhNfzHuXCOCEPDsqfGZBPtuyigs
LJCHavvWq46Suku1c/F8Czy9fCv2sJtrrBtTUcI9uD4yYMn2nb8Ttg8DToX+ivy9sYa8kYrTFVKs
FsDylijNRTpTI5iOzh99Q3HAPb5w8Z+IEl/88T2IuSG6+jwCmj3HwTPI77/IdD7gmSQoDCxawyLM
n8stSCqLaDgjBf9ew4KS/+hQEE/Md4HkBMcyhvM9MnqNVWEa9qJAYUOeq5zagYWv3Fme3GUZflPj
3zMa3AnIKh0wRUkY5qLr6h8z5hIU2cH4cBOXRSSOyemlgTKWejGbplTgVkMRwqwaUoBAObomPJlh
VwhghsSqj+tH/CLDtRJMUpPWuizuDX0AV40MDXFo3l8QvSUKrsQYoLphEpa5mNoj9XG5b3NMgyti
C6VEtDBYX/eHv/KUiZOXdGOCh1MuQ2Fv/rmobf2Bfc7TGJlOjRf9YsQtCWTe/YDdVTpD99akg5Ik
pmDyLrPZWiqlQFRCSLL8QewMqt9wV9iCGJRo42SkrMqvc1fqzJP/7ZYYywik1KZWBK02hgc7kBD4
3BglLK2Qe7CgA2RR4ksXx1Eq88FXgQ11xkj9NVq0nzJYotMY/FmoBt6AxuEcyq7s+RrAABvtqQhd
qKP8Nvl1jvTn3NygWfGp5otNhI5Mji618qSYoKKr7RWavmEKqjOFkmNkoRU5dQw5u1nYOVGjt6mS
1gR3BYQ2mkTfSzQ9h6TEyRo0BqUjSs2N2SnBiDMOmEx4GHIydhHl95nGAbLqTalWsb/lNX0fsMRe
BBo1v5QPRTMCYp4o+zcjwJzqm1MuAUsAGoMCT+h8iYIiUZ6010T9JzkhlcCsidT+tF7Uaytbx+AU
PjB4DDV/S81e+uGi4XKNPKmWxhqgYEq9iEOAFf0Q+kf/EWOgSz3rkOuJJXRgfoM+hJ8R8+PM6UZ1
Q7+rwe+xxVibfeEeB3jhDXjAWO2VaEgsQCJ1fpF1o3T9nHorcv4Yp/XrTCeCnDkYXZIvxxM0wLx9
eWeEhcwB7g6QsdD+fXn6oHIM9ZCGf+zWZJEudOODFv+cxNikduvUxzI6tBql3TM326Z61njRfkQn
65W8MChULY5VwNKrGCjmgrjE5KhHpzO45/yUa5aufSg5M8m1GxWxTYoURMr1Zl6x+DRhkH+XQN00
cgtztd8pmVFbRKHc0OeFpOTgmzKxAoCrZWvrm4ODwMwSPTph3ZgaJgf8+vbLMXtgtFzyttsKR4p4
B/Dc7g1EeOn/DcAghUSAh0A6zYcaWM6w6ZpuQMzuM7pGqQOvl6c9tSS9TmM1IVfsY7T6S5fgLrAp
pYObn/zII1nfWfKJvfVcj2jBsvWpB0E7ldUQTyPjQqrcEeNdoEe2JJdeoRzRmTpzdQQVMqgvwHrh
qVnIY5kwxbN7/8jSP6zikXryeLEnLNHBoaG+QF7p9drg2bEL2Bxh7h6KCpuvEzmRr7nrWE3Tow3m
aHToKcSk7OWdeOA79XnzmMw6N5wn7uD1SExByMdiRShLUG7H1EhtvZDZECHUoUJeRMGar2+0rdO5
W5qONayN0zoSZ3VUluaxaZpcEddFgbcfO51gn4Zr3F4KtOXUyizbl51wPpcX7SGV/OW8MBvpiHWi
zR+Xg5nzX6zL/xf401nIMvzr7wonbzURnjLeL24ATXpKMcsZTGEr0YtQpzpq2wuty9SwKsBx0XdD
hZ149bLU+P1jnlJPvQj9Y2Lqo2Mf/HqaIKWXRrmeYfGOt5skYIVbJ2thuH3YruRXB/emYVLftcw2
Uotvt5VmsmK4vtf1X+ulsMsYORxO/LZuoG6BgZvGFWi9GPsfzNYr4y7XOnuSQxuQmk/+K23V1mOO
L5Uyi1FsSJUGxo0Um0w0I/pu3Urb69jUcbnS6DwlpP+085QJRD0xwyEl5vPXIuHIJWKvtTgihJy8
dQ65sp9Jwp41Kj0AJL/dOUdAC/iXIFO5QqioD0yP1ftT78Ar0gjpNs30pwDsIbeevHArOeTutbp9
4IKqrwd5VM/WncEjZdm9jKf8VnH2rI4Wd5tpvkZzmuFTHJP80ipgRV8miqSYGJYEIbpNd1xgLzDq
rMHhzBLnGVf2Y5VPrbxLxvTMCH7g6Lh9t+dLLLvVNjWpQO+lHSrtTYVxn1dvsfS8MJz8wEroN1L5
n1bhLDWMk2ET2wHCcXLgtPwDuJve/6YuBMzh7Injs5YMBGePj+1WkC/6qOQJyt0n9EwheaFWxYu/
OLRYtI5F8aLwYAglauVE7F2hffJy9A7Yu1CmPp2lqKD0aZPcd7ij16Ihhlti5vYHmcyq6iqUsTzW
5RTNQc9ikhXi2Lftq3gUgTlRHBjNF+NsPd5Fpqx0B7YJ455lehog27HTW6qgUiR/NZBJ6MTToEgt
Y+ROUQ/VuiabYMIi9bhPNpTxKj39KXiueZNsvFV5VyOfmmSfup0jIzPQnG1ZM8/n0PdrQ6EG/V99
31HlT16/aL+gojWGi+Gg1qeQAqj/1z1n5Kw9KMtWZQenqaQLyjdv1nWaxwHseTSLIi1bHoahGYPS
nKikfU6FCHXWtjJa7WWFL2ABDqzMhIjZNSInJLxxYgbWhfM5f2Wlt32bqY/qzTBO5kmU3cltHIe/
1yriA99Nqsu9yICBpuuORHcKV+2KFj/bzeWH0CtVhF5f6j6WYwtNJzFrsXLzaQpIfVP3ZSkY3w/f
FaDZ/AEKupfR5jEQO72AE2MZHNoRjqE5wYh6iuq/26Gh5RXsfWVcFQBGJAozFZeo+UzM1PrfIQuz
fFr6Fmb5CMariz/WMnNhfcoG04ijjuVDvT6Lj0Nkh4Z6c3Mgc9NVcJORtq0dDrJv5iQAsFkQd0j/
F+CcmW2B1+BY2Xz2HY/BzFcpe/F6q0JuBjm1D6oVM/bsRLhvKxklOFlZTgRbsiQ7NBc+h7mcTY+M
evdzyf07io/Sye1HQ4uj+vSBr5Ko8DGS2DmYq2ZmYRmLZLmtVxu9g7g3hjbqjYxN1zom1dRpLmxL
1yPuuQe78M39QtUjDYOyuBZ8AslvlIwHe21RUppXEn1V+IQ7AIQdRDVNDECaMOjvpFIW7t16XHxf
QoEcBKFACDjX/EWsA5nt5zgBD4AS1BglYucsV+zp2xNDH3FLleF4dzR7wJYG2OFg9K0EmSmn/T5Y
zo2+HmgkdQtUH/sVbY5c1BEEyZvXU7Uag3Z4lw3Ay1En8pFiSphjYMIY6dfx+g8/k5JhZlfOse2z
0D6UGMI9QROljZUaGKFj7UvkyCQmKNfC6vlN68KAwP0ZyT8VJT6c0ZD/LHmahy6eHF5KI06DFe4a
Y46YbIgN7Z2bbNoHSvt/JHxKhaXgeVX1TjcfC6ol8kb0EHB2gbKEQtC33UmnawrtydpekGzsBDer
bjvIIThT7xKBFXl8dOV1qZJMqYp35ka69WldOLPrE0igvow7tOheyHVN8j3YVs88PYwdvpHzJBYu
LYn7IjhSDO5uI+yjQz+xA6+mbu5JciWdVmUmifr925mtou8CSHKS6eLqtfkKmx7kAHeNglWhpkpz
Y0ljKaGi667zfznMmaUd+Or130fnZhuKd+jFVOJEYyyXVqTyUbWK6sTppYxJA5OrZc8Ul1na2L3I
zDS4J1UuUlEPOgjbWIY0AszRUW3sTARHP5zPhMWs36RQlVYtjgQCFqmNrPVL14BUUEeSA4CluHei
QUhtXFtnGiAr7eTo1ecy2djAc38W4j1UPKX+aHT3wT+l8w9ubj2nSKv6cwZ+S4At268lWgh+U4HI
69PGIrmG69TFQvY0A/RIJJSEDbXsgJK9W2crOgnPUUnk0i/YVW54DxP2Jxxv3ve3Kd+M9dLzeCtR
GsIIoL3V2AbMwS1Ar5sdUelQAB6ff4KoS2Udu9rjgVPQToB0agMEwhPmwN0IBm0TAAy3VOAIGmJ2
kl9Vrt3pIuBhlOobRnqpfLpvOCqSTC0XMm1+c+PbxFtC3GvfM/zGYHKr+7k2aalyyeIhg9oeUIhr
eDZ1VhqqSKtYE6hpqP1jYyoHreYnSxXZhHNjUJYMnK/eCDHpcK5Uf3D6MGXDi50EOCuPM7gPjmE4
ppntqvunKzIpfzQfoR5cICJMfstnpKEre6MhMdnN426sfEg91Q6MygsKZyg3YO09M7qDE8lsLfgU
Y35/EgywSxYwfn8CgUI/ctFwtCBH8KJTuHwhx3HPeR0Z+S3YsiO+F7gTUJDCOxMGPNPSCNxRqeZc
GMSc4Ijbcoe1robVFh+PNf1jB6qbDUs38Yk6a26WUyuRja2dK+lKpM/wIAOsMnTmETntke5I+5pz
SUq/7y+VWtsgVi8GIvvRTVN/NCeVLLS8ixenB+I/1SxWAEGxZQ+w3QiCmvIWwX9OV1J7PEAtF/lM
dtaHM/wLRLxwgtKQb+HimClr1wNeOE/tzsd+yq2i11HcK0P5SdNNVsuRrKkkx7YrcMw9QPCr97x3
oGRt5OXyfy71QanQQaMuomVV2El+NuJkkDbIiQzmsD8kmkaEgy8g7ajV6PdY9v/wDum6fwPcUvT0
k3HlzAtLhHJdWUDyrpy5xzskgV7SLPO5dRmyECPRhey6/1Ur7GcRgUX3tqkH3AZ3EVH3OT76+JWw
iTx9MnKbYrpIna+vfPxxXN9phowAHSsLI8UcKqgt2pTOPKse4wrgZKd/IXdEZJlloc81i7cnT+BM
Z+r1KOo06ZwjQtj3j4fWmzzoNt3BKxJ5tf+1mAt3nCc2RhGy2bH7yjF+Lx7VZwTI/MJg6R7o3+P2
yFUDq73ENr9u6qQ6HoIxdLz416eMzxmXAsclsnMlDy1sH+GDfyF6mF2VxiHDwYJUi/Ad2zAJbtLh
zaIseSfyMXFYNyWbEBpi2NqWYV0wdjQrnpgneGkL+wafFSANeoz5Hxu9pyS3R09QAa+nac0900hQ
/HH35RTwefQHq57nH+ffDUxZHuVKNljzczqxg94iUTQdbA+O4iQo3Tn7D25b2JYL7o3bk/zjlci+
jRI8J61lqZh6pVMSOEQmCLyzQ4uMiPT9m0nlH8lFTDe5047tz9m4DNb7vwgfHsQ7f5wOuPDKn/mk
Aznxqu/p2OC63FJVnhSUb62SKPzTR59QFWIWcSiDYQ731PdZMB8O0Imv7LXXZVh7PA+CvoAH+BrG
6K9DKP/A606IZJ7Ncgs6VBg+maRIDRnKaucgHoyQzLhexRcexzJbt0uThCljKrVdY7uQe0oijv1g
glyIUQs9K87BXr0ku9CJJRByXwU8MSC9LvZkB6e7eigfeIQKINHG5+ObDNN7CN6dSQrDm0ffeMex
Ou1s5TZTP74axf6YIWOh2moqKwvCkGOwF/WgVI/eFZoD31FvpEg5WPWPJocUlxRtBsNsWApUYwdR
BBzy4CY6OJOg2jHSYBl+cHLWvGSBz4BjZd66fimjMzvQOOCaTP4WK9EWv+zY+DbYzbOPnGg6Xr/o
/hgEKnIk1HL7cYRQOm/o+H5hBzvMKzZio4eFz5sldyBOz2LiR7gEO6jpiP/tdv20MnG8LYJASMAg
g4QAp+uc6BQ3PIykchPWNhZaEd8mULF2uhDoCKMYcOhDNMS/qE+9Df1y+GcY86EVJCH6TacvPMml
LLlTQZ6GdG5rx4755B1bt7EXnOWMtTtqQX6vkkozb5tgcYYkm09m9Kmlj5SgT7ce3TiC07dL/1Mx
u6iv+LSspTJ8sxpxV9mXuvDwclt3mgPHCJCq+lc9/BJl6FxJL3z5wZKLOs2YgwIk52RpEIPnv23C
+4i+ec4txGRQVqvoWrO69mJX9gCi0p83J5d0Xp+tRH0tnGv1+btLnTunTODjT5hFvUcTdRQVA1z+
vzXU7uSt9H2blqy6uneUcSPz1fW4OYOFiRXffna4qcZLxIpomNgIL2dtgzRho6/K/jNwpZbffOMY
YZQditRrTvfBXMeYxqx42UE2VQ5KmM8rqYf2EMq/k+wFi4vuVyhDORmcbM1hj/6eD4pTDtmU3AAd
3djnImvGF5FOfFCp5PkfbPXXbijyybaKmT29Kbp5ACmu9l7nqaFN4IfjqMLewzIVMlFU/WKlHez7
3VAa/BupJjk+oMCDEWUdd0N/4reI1uzKymAB4o2u1H4hZ37IsjmSb9ivskbXmxOnBz+QtAAbpS7f
qMAE42FiVXwK4KT6F4HajMnKVs1vM4lbxmGmVJ4lVwFOyi/mR4fm2ypv4M6XhhKv45k/6re4IczE
wt1x5CuoSVOLX8ufZvpstfJa540TOi4w6T+HQZTmr8n3jEctTH4LzY2sKNI3K7IBANCK6A2FJzuN
30xRuFy8swXyz/s0h++YcaLHQSZzemA4foXjyScuZEsZApmlKQa8XDIQ1C4ITd5fh4oq4B9t+8z/
735M7KxX4TG2Zmd/mTve8x2zo6BOqi6tqgNX599abEWSfoH3YulhNa8T+FKu5cFz0F4Y5/6I2BUv
uSQNgn+mTcjTcROxNbhG5/s6aOQ9TaDNdb+zfueO3AKuzVRcYiSC40nZDXsR0Rv1hzxXO90nI38B
EoTckt42J/J184j11OGJsDOEvINzZDXHE5Xv6yJYvCu+GKiY4agxnhD0EjBUMXV3ieRyMXVylD1R
DSbCEtldh7oiM65JkKovMj3bvSfWsCDvHHTAI/cE1NnE5BBJjgtcTKPtdloJuSX8rh8rqeKvi6zA
IljRqwFHkRcBWdyPjaosfbfa0i4/OOQuPNHX/yi44mf03B37+mLLPFKdXBC3bTBaqru/d+1hgVXh
eGunL9Cy/C0ucsStpfaunuueUjmPRGtoBZ9iWjsoIRiq80n5jnHq/94gFQupZnLCKjTm6YPPRYS8
JunH4Pl37LjOrdpGLzllbVx1RtrcIR2L38bdLAAaSgh00sWwNEssDjUmTO2GtPN8Ou8N1ced7kye
SCM+DRyq+Bu8Zrft6vkjSLQPecC+6WeJwxaqMMoWREqGfVuFFypjdqLl4EbGqfDUBtxN20y9X3N6
oRrn7wJTLV1ERt1kRyKzvRGvSF3yusJ+hZ4UrpMzIhwYGIfU/bpvKLfFGxCdGULQzZ44jMjb6cbI
sNhJDoXhnpThs8V0mRk0GcWNOrK+c6+aHBG5OfJrwstlKNco7IobX9/PEFqT/BqbRmgDQhYY62wm
lZh7PL5Py+3Dm4j5q0WvHY9NBsvPRT/N6820oGLq4D/cKpDRK51HRM2mKrHV3nU6unOg1gE3x7uJ
N2bIg8foZ5OduJLBFbBQ3rJVlfjlQisfCBPuq2DmGq5HUZxzSQHBRdSazyQp9aPGDk5EXtbcvfPn
XJ2bWDMawwqXuEX58PnLMuwRXJlE8IjCkxKoXKDzPGDw+T7B9W5uBO1ZR3Jr7IKJuNkK1vTKp7Zq
RFockIo1ADWeFDuCrgCHYcsa507DB7A9zYy1Bafk1vsEEHauQp49iQ0Wy7vseaHhiO4oSZBXqzwW
OjWNMUuMEhafvHRQWKfJFjfahIUiSlYFiASwsC+Qpuu1CaXnm+2MK2LAiK1gArI9xpandLRebnaU
6RyywFBsjExSsubJ+RJEDAGoBrb8UQphJF/HCVDqfHhbSErUqJdS/aEq99DrWnS9RMa9eORv5o0s
I4NOVIiBLZc3Kgz3Su9wWufHhqC7ZYcwsUUhjwj907d8tiBmXNuxr6pINjIZW2kUi9on/nuyofGh
P04sgSJbrSKmXJPosgVSy0JfNd4o4a0QOe4n0+ns8GHHYIf9KJbxFK1WCNrydCe5UM7HcvvwJxuf
HH/ltGE0KHRsRLAdqQgbhRakSQp/VvfQQViS9Zpu/PeRYoIczaypbHZXErHXOXUdiUx6L2568fWd
BEbHa+tgQTkL3qRdYCm0wlUEuqLHyHVOcswKK3pTkeccXNb1oytLPtL6XKNoeYRCIEvP4dkn+R1V
xxr7Ry57RG/N6QjnrjoRFgsLfvC6wxTgpZ4lGedXmM27cQFZ8Jf//5rNJGW8Qa0vEWMXku0qGynM
kiMo3wTRlzqTC+8b36kasiM6rv/xEqn1PSf6kvHlzyNu+oKbr7bq/We4xSEL1rLMXX5IJQu44stU
VRus8Tkd4dQQtjfYoasAhDmj580jieYlfuL6KpTnD+W3AYkO53inrS6P3/5VzcOwNYGgY/+DIuOL
mTCeLxw06eG6llX6wZ2Aj99n4Pm+xcfAwYEWy/hwubpxO/crRQiOyuEf8uGPsaksDLUc7GapRs8B
ESzxUPkW4cH4wXoj63ukGaHhyqykDyKq2nKIFNjrKggMZgM9QFXKOIV2V11rNSWfg3kJYZ4cmHkz
WtxBcby7vh82QSHpEIatFThRTJEQB0yOBNg5NF9xE4L3/mRxWbo/SUaAm4SgWW8GOn0NYyX5a7/6
5z9qfKUt5q+xXGuP2/yNkh+GCmDE3AUX0AM4BSCzXRkOaslsWyaE/ToJd4a3blC80upujM0pSv6c
CUiAZa9dKEPiKJAR6VhoKfbVv52DIGUiprylkb59aLJ8mhGj/+JQuYQgpNu9jWjKG8Broy/GMoCO
VwYv+N4mNCtsXpT7L2O5HdJVSTTmQ+DwWPwI3cIWytODUjviKM5E1kGvJKok5rG4iTfYN9owWzWG
JfHp4qoBnQ89PSVMAMQQtmZGiYHPs2NF79jn09u1HJAbEW6uaId0HRDPqyOVVap9q+OCwxLZK5qL
rW2C4DW+iqFw6pJrKIOVjpcnSlIvOTkJVxYQ1abSu7RxWZLlySvWs4uvJVPi04crzyVB9sbRPoTM
mcxIrKdCNWnViCdHa7/lvSTOx+YuRrqMk9D6YP9SwCMWdQd2Ew8fC2PvV0x9fVL7iNFhaR3zq5Y3
VGq84Q+qrgTVxL9pc48MqFfDeca2I+1H0J4KnSUZc84LUSpJ8WlmGbvBHqgWBBNG0tQqfbZsQE1q
dW396RpUKrdDkS9Pjhv0+/p2b333h+YQgtDoaXjflJdVnZRsOOJVVV6eP/7lXIKLMBOgdgsm7lOO
ZCdnl5JSlKmGnSxV1HspQ0c3GWdc+aq8dD1WWiorpIyofSUfWwyUgfdKJMrsX9bPqCIeD/Fp3F3y
GGihO5TFPEYnUlgRUElXxpH9U5st9KMnnCBbgavSvD67KAzFq7zFU+cPZ+V2Xmmp6FqdxwQqGKXz
T9Qbcf9+pNJC3U8WZVkxCJbK2n8HU7c+mZOIE/76mV8/dxMakqkHFcnB9o4aYpOfQb0cZ7iM1RzO
XGNoLY+cHA8TtKh2q1q/jyBl5NusPdx2SGmSBvBf7RJ8JG41a+NqqH/DbtnkWxtCVKe+scZMHRDh
xAZCsjrIK9S2sQZwMXR0zTt2UGQrV0FavwZNt0/g6HoSqy9CXGDjUb7UIZfGXM+aiuMEgni7ra9X
iBvWgr/hpseu8h8NnAsPlwoEGnxYdJ5rpgqaiG6hCt4uUaA9J1utwvI9FYULfVZAxRsHAjxeFErx
POLHW3HgeCHNuzII5kd5xYgDcZpnRbJJvpnUHT/pOfFZ2Lf0N7qePYJh6EV8WBKRrpYy2Bjz4yGm
dSYry/AP2fb9wIVsBWrBe9t1t/8ccgbT2TdJo66B35EnXMeg8c50PTYi6k+yJpSOrC4KDkmUyfow
3aW4dtMkjlCJcvuUybJdhwN8GnGJ8FQ76GNcLgoSBSHgop4530BYAmO8xMgRkYN+ETHhYlMCGtWw
BG2kU6nvQuRNgKUNUq4+szCOR0ydL4Yw+h5t8G0uDZAm8b58CyQPaAb+3FGk/Ct/t/u3vNUNKH93
U3/FLC3oPcExmsHpXZcBTeRSiQcftuhPKCcLq4KXvOa2qp44U5J7wiapO+2s2ILbnnUuIRjLmDLi
FHx5b97JTcbcfUs4peaYoBtxpVx//0ai+AmtaeH8lZ6FxyK6ksPhpP+J42Mhht9IT3xelLOxGNIP
M5EWHpSYprhR8nMoaYnh+0do3nJXcb9344GvmF3uXVlzsUiNslK1KBG7cRNv/mnUX9Pvdj17IhxM
NvoQ14buhW1Do+q7Slol4aBOAUucmUXKh1KbqXvN2KVoglKeEbI9SP+YLmwURaT3XxWgaU/NTdx9
Ccy9UhWAyVgTwNPW8In8TdvECmcMoT0V+iNFCY9+7KD2ut/uYvhzn/ypYTXUI3/5cgpQmGR6Nyyp
ENI5+81wlR3JWf4zS4OZPulk9EGZ34YiJznHrSf/a+EqH3PfkGnNObaayC9dPHrvAafvOWV+b95h
O9ElkYCBiXtIZj/MD/BRJR3G7oWvoRIfyhgEqlgnMfIo1yiP2z3VXB4ND+8Qi/I8GJOhBkN7Nqh+
nQFTsOYqjOpH0VO3Md+u7iAUjChtFVIELI8OcSFWTkpj6H5bY0sviVybBDMK13OEaPRdMo+0lF1T
QCUEwhvP9YPRsGr+dg1/bd+tAsfZKhnOPAyfhDAWlqn9Lu/0UlMWMD36C2+8E0tWL6Ry4W0/Xp4S
lTWM5bLVjNXNzGKuUqUwkOMlwfFIUoR5kKCtDj37+oeOcQ7JJ9TIzGj0Y0KTvnkKdFKIend6h9fW
DNEWpPJfmtCnTvxVRhQJtvdmwXgLP5vCbck/+Y3C01O+qPSFPNgVSRs/bk/rfTY6CqSfQVq02GKy
sK3URiUzmdqwFs4Q2CfAyNd4HQQqIZ/WvygpAbtO4s6bZqb4/QY9B1nNoxIN/PVsNRVZn9HjWLk+
i/VcT504uanOkLf+J3sbmBG6btbaF7YZHvcalZPLrQMcnDfQKFXm4+RfhSILe6GEQO79TCw1G8d6
2NaC7hVE/DkChFt0pjztcE1qp/ejqM7POJAHu3S2P7sV4Ira3UjDwKkCAWbPOmo5A+i1nolSxCT3
/I5GITrxcepR7cDwMFRqpbB3e5MHFx5yzY8UilKcRU96cNGlaA7ODwTbo1zCX9FgYuoMPxvki60F
wRnMw7gYsIXgdC6EToGUY/EGemHcHv6dghwLzjLe55ENfybi9JOwbSiwJsSTUuJCjSclivaQqdOH
2omTIwhTYvzPHdidH3IK14J0TJaRlUiEtw6FAOP0E/uaRf90ykJ+Uwt+TjSCwvkc8r6rx9EA3957
4EBtIf6LeC897myZ1tKsG0Nzb10ndeTMQ5OwU8mv8B6jRNoAT7emXdaKuBGwUr1BB0lpLEK3heKT
HieGMN8MeVbgrh94NRegJZHqItRXXDUqSUUQ2E9BUzGDliWnArlISvTRjTtselAChrfEA0ckcRbi
q0DKiJUZDmNHlmSTnFlpVyCKIqauxBWWWHEEhWbVEFPWLRtqrKtxVF7El4XlreKctF/FdurUkpr2
11J6pUFDCtP8bATAavWalDwlkl7RoNgqf8izuXhcTK/z9iqI8idA++J+UO6Q44EnbSJ92P2iOkKg
HiGJRoAxRPQdFrBZqJ6oUQ84Vw1gKDYzEm9i2gVdOCU7fDjy56lx7CQljcpWoR1E91Svn75xqeL8
69Tqc3qtVJGfF5W9ua8McQ8nFtyDpavt8RZ01nskhpThv5+DTZK/KriPLmkVNDkf4sQu05mLvlG0
ewViVVqZShn7ZW1vb5gFOxs4Gu9oUZSORvcintiisH9em468AAMthGqHS/Alkc/kpdXRwsiDds5q
BfOuvf7aVMMeYMHaCAWkvYVSyNDBOHS0MOfZIb+cnK5greBUSICTne7laFjbOCnSpIPQItGTsrS+
TMPP3RcF0Dm/oFKdYANQv/1zWogSSHKL0SlctkU8SMtG989adizi4f06S0lf7V9xjO29fLMjCDwx
jd9Zryci9vGFnlDkiH1nKklkNg9NPEF2scTBK3SsHFSwmGSSTEmMwvF4GbMfyHIoJwBg9BrwwL9/
MrhNdANVFmq1JnSqii/kS6PxRbuvYgbMKdznjM/uxVULvdJ8FBsp8GlLeRZrEZrODmczcRKfLc19
oAcLmeo0lG9C3ZXI6hUs8ukjifygQCeUAnn2nIRKwB7LPcVMaxg2jXOAgnfQGO03bEHREgLbHutg
cacZjrBI9d5eTWMgH7sHTbyVrJvGMFlM0+05/fdTAzCQgE265ZU4FgIENLBOG0Y6XoOVEY3sf8ZA
NvVuvGcNNLzW9o4AdkaLHKz1XfXgtGlirZ6txNb33bPsx34rm6DVfso6oP9iVc3EXvdbUBr7aYIU
uOcM24wXDehnDBNfmQuL9OZf0OhTlHmCbIFlDuAhIc8iXSubeYdBQGqN21xmjjQlD8xdFWrhsETo
2Bm7REaR2xaAG/1aliF9Xmmea6gQEu8nvPW+XAPnBPmiYcQUMXAGnil4h1v+Li9RR/h5q9KjwJ+S
sPDL1EDC3QRVFUlleLk7IyjkKaLnanKzJeQeLXVk5i6/9MKju/7nzEka2BQ2lZkRQ34bP38hbu2U
HoSTnO1hzP0j0xS8H7Mm4tGn2ETvwAj1OGqbTXqnfi/5BVj6rIwBsHKh8YvCGOjr/4ct3PNNubM4
zo2f4him+VA+RsL2ksCHjTHWmQMqDh3AuKmd9DMXW0q3pKgww6gL4+MntpSHCB6YR4lSsrbn7UHr
iHR1Um9k7yLKyYlPwLkOfWqaeSOfjC9obqtmrBwtgU6T0YT/rENqXNaK/l9YnMCwDqTKL2SxARxI
0CzQ31sdaYRfqagOxDrJACdG8UfuWRkgte6EmP1EGYfSaLJOHGyijlqVp7yEfO/+EOp1X9mGBhpR
L2m3mHfPc33aeQgJHohe5y/JkH1MyGo2qZTnmUEgyXDjAtra58yMXfp+lOxA1WbLd1vKPX9nWtZg
8wzzi2fvPCNTY6ZTwgljNqJv7Jj+h7zARfEPcHx9P3oS4OYAscOqlOLfkL6nE1qxosUW4AkNWrmb
loMfRJp85dXatLbM402umsTY3FevhigP7eyz6ujXYz/EZnwR7CNQ/g6gR9xqQhPKkb/0N66JLcfY
OipZURx9j9ccN6q5M53GgQBlZIrmhA2f6hTYTTEzz3sjBN1H7zQPT9913lXSLkOCbSzD1TZvNwRK
MapqcleQvLd3o5uYlwdTZpvBcmo8RNBNOO0PDiTttBUhYzRfBmGBSd+IqmTL6LBqhBwdyix18AbF
smTXKKbxzjpJ+nv21hu1/M8IlMn5Xin2pLzNp+iNMOSjH2pAbJJF90X3MOLFeMMOCRzL70rk7OdN
LtVMkrWF26gCUhk80O+AszIUAKlZNPxDM3js0lYPcCpnYM11xMU/+Fx40BpeNVUAZLMIOHNC2Yff
Dyk9z0hUr2HDVRW6arGIQxzfWXHBIFA1N/C4wVQcNaYu8opyc63aC/fHmojjZMyYOBdda0yLPKim
WrSnF6RLHUrbVVb+9KM9Agqq3gfn+KBxdGvc3Ao+yRk/JrBcdG5Ks6Sdw9z6xO3ZpyPkVK50yT3V
jPMcY3w89p3srwLRyYA4vx4f/NDB668d68Ga3dn28qKuVbUB5lrvVW+Lmhr9M/vDqExY077R8BQl
Utr0hatZrvxnGHk+veZ7ZYImkzJjHWOUZVtxDUOK+QzUFcV57+f74cnYhYHuhN5NKZcP+Cj0ptG8
7uKXp3UrlMW806xbAuJ9PMAsX+aLnLk+ciVfyt7Ta+NLZnElg6o/v1Bydb6eGvmShcklDMl1/D5Y
Kju/6wNxRje3OeTxfet7UeQ8T7rjwTrqYcM5qGR0gaQ7UeTOburDYf10zkQpXPJ6jkeToeGuUO/y
4JIpZKv2kWtk1Lo9nArJTrmNBQ3XjZQMPTfzSdU9I9QIuXpMHhbkxv5X3TSW2NgdUuutbQ/X8rZR
yLoliS0VOOhvGbqCcXuKsh92Xf7RWKiqM2zIcZhWAbbLPIHhLG73AzbQUUMXAnY/F3L6fJ9L6UKE
Wgn45Q2MGPH+JjFdW5NhTHSWfhO3Bjd94bjG+DvXZbW3YefEoncoPH5uTQyaCbg93PW52pT+kucH
QJaDzmw5acQlg8+qFT/50m5wbS68aC1/YIpOjpBuAxtFDRVWi2AcadJgOW/NDwovSFeB7dZ9GW3+
v50fjvc35b0GVS1hH7+3L1urjCrB9YxL1NXBOasBEtwou7/yOchvyUD1lltYjxb4N+c/GCwebz+q
FmhNUTfEPKWZCcG9WiK5JJ2hmVderwW+Ua7uY9a5t0LqRYpEAU0b6iB3Gt8RaL7r2JnZWYEJABiV
4d2jJJ8OXlsfjyqE6sybFriHHYBq3Omtq6bi4TXGWLqmqMxTgnqNpgML4/dCNA2oaqs7AHFAnPmj
jq4i7SbGCsqLptyBouNBWtzUy5YtcpO8ec81xcgKPGCOozmTOC53s2plEz/45WGgiPwio8bxEEUR
QnPJHEZ67IaoiE9YoIhoFdLwha/83mG2K2Mia2zR0zQytD/1I7hFbnMRSWqsawn5VoNXVKrUDXDN
47YxVkgXtlm4Do5pg5PQojkNBFMcutBalyYxQFpQGA1dpIwOlO+nJpjEv7kJthOgXK/AsKniUssd
m2ppAdUlp4Q9rtlCjQ9UAx/UuJkyRtfdK06jDVSmkmocXXQV0gTWPY6KxJI9Ele92UYZ1AhHBc+4
dMzrJv4wnFkUOpLXdW36go92MhtzLmIUbtkssS+tU/ooj7VQ35GZULtSly0XLfKl0Be+3H5SWUvv
GUyh6GAhREw3/YP2++HQE7BTe2UOQ6vMQRv/T7SB82k8W/vv1hv8i4numUPLsMdIL7QROqXlHVgn
ewqonr0Q3/ANKw++MgLwXzaR+CdCSKstKDjL19kHVCOiMCAm6PrvCpMlTBQ0RNAoJ5sxF479FI9a
L8NL9lxfiA0ubTelyQYU8NQv0X6rcszd3RVCOhIs26NLbJnShLby7WzSfDcK6/9CkQ71AQyIg5kc
Eb5xk7xl8nH3pdiBq8PGcxfN4LXsu8rIJmmsRdeGLlVXfeS8xu55SP1D3+3/ws9DPeDOCu6Xtf8Q
dVzXklEPQOVx4HmiruYwNe9+nfrDk9kN4Tl+hXjYp7lWBT0M1s4Dkue3ReKL2WFyJYhs/3MrUBcj
Kf8Y7Rrm3jbJf6PZd94s40p9uGICaG9LxenSltwDiVg1bEgV5VQGQm4yzAD2Srx2zWCQCQV/vD1U
ya2xldwuCsSMxv0LBQ6CGJGbCAbajQ+CWvOmT3H3WgrNuXbaUkpA4zvRYrL1P0rH+6Juf1wtk+d4
vFQXn84BugUbIF2jhhktdQD0zUFR9//5nzBKpMyjp86Of7tg6id6kia3mvt48vrH4ECMDlce5I6Z
NUaXptmfKb9zFLeG9jw03KmAbJjY3zQAlnI+hfCjqmyPJ+2MwyzEYS4wQLy55bLiEkQR/fZ6GMId
2+QSFVjSoBl6rkqYVyx2qRegkUZIJcfqE2PuE/y++GnCRqfifERj9sbFgdX6xh/d7k97mHtn/unw
t/wi2C8jMYBG1dSQCgsge2sFFz1mJjjOzIRaYLnGKZf5vrou040aXdkNzN3+cfvLSdAGnKBcjVlL
TJRQoYAuXjvY/6gsrOj/hxPyEABxRT3NBYCSSx7SPZoKhZRAvtMEFuC2l6yUPnMUqpOC505ymTs7
g6KcoIyksV2Kn+DoaXW2lFy25h28cKhPCojzLRlL+bFNTnLoyDxxwzu4qlVV8qdN8mYFJgWChHVx
j1m7/LI0eMvDvXji5c6TOmZWAb4rk/OzYwWJlS8EcLNklLrHHeHb+L+URDSDBBN0tgYUdenhs73+
KhqSnVzXPT2zUkM92ZmnjYKTdN7AjOR/ghs0EoKSu0mJ8quA7xEHxjlMUDEB5sVnLXHrLwfIvyAV
D0pnKhjw+fG5pmmx9m3xce2/CB0OHRCJd5p9nXLazmQA/gtneHQEsTQ9cRYqcXRuEcw4VuiMDjGZ
BEpuoH1jgKcD0tK8TbIRq+2XJYAYPzAIdPLcQH9Ij1zpz7U2/1wJGPrQGZd2b7aXtQTGD1xRdumR
/6HtRtWb9hjjMyMbWpoAIahvW8nFnqGVsNBYltJRo3prwz2kCt86EljWrXJYHzQCgA5A2SHZSdvv
AL0W/K9nHKvQhkNspt7wyzJl4nteg2FzELGBPzDKIDIb8/dVHoxWVjFQINCXufXo8bPI+wrfwYt9
CU57BbqCL5v8OddFNFcI3mChRsmDWSV8vedkcfxYrdWRLj5sP7yByKg4/AYkFtSSb/62xUV7N2o3
YsafVypIc/LYXAceTAbd1u1u5hRP+6Wjq1VxUtVidSYMr2tK49RuazqPswW+/nktr/dkbssncFCG
lljttXkwTUQ2i47FwjQu9pLf6PynPBea6980in5o8R8rMQtLmV0FcaVr2cJNKhiueTXNPER1C8bm
fIDTRp/sK9M7R0TfdrCv4dcd81EMQPvRKIAJsaQiKE9UcaTi5B3qL87bRkuYFsk1dnpOTG4qEkH8
Ny9pq8zv/wBXC5DPWcRKdmzu6aV4RtAg3OlO/wWh4J0+fEAmXeZPgvhl+y1ycrw3uWRQjIEsR+uv
rnUEXc8e/nkQ9Pv8JbFt4MiJqG1+a5CqbJPhqQWLB9KYiw29trU+khilbactpCMoTEJkcikGz5QW
i3KLB2EJRqiM4PKOI/TKj8PWISkvZdHkg1WBHIPBAVDs0rahNqhIpaOuLyVcXbvfx+ttZLYsbm3h
g4jgYPI44BCMnKMd4VXvx/nxGDxcnjH5L3Axw6CDcE+ZWSRjymoUgT99JQt4MA2bbVmnZ3trHVtt
lUGem0b5zVrxzr2Zkhliixn8/cXGZ8XkhY/4H/qguul/sLOqCTxHsW7HyIwNjIWfAitAGidtgFvD
K96V8pzVkg5XBaOOI/wPlALLWPpFT7g7/XnM2BhcPANDCYOcX3Oqnl3BhB+Ya3MJS+xvg2XdgAgC
3js6G0hzeA6Ot92ZiuOyqRgIiVrSfWa+bZxwwJMBOf14TFPmtDTVr9+qaBam8kzbk5nRw6fsgUjd
GZwtaeEsNabLSTGz3u4g9nxA27iBtm9xkQPFC0ln3R+RiEg50kfz/AraZaXshxb7tpeR9MHE0WZX
ScB/BqbfDSiLsw7zrZ+vrnkSq3jcxu0KP5S7cw3IeO8BwjAS2cJZSRcuAcmS5pqr7D1/mI+53Nq8
puSHBGMsqGCH43f7kaW1rDnUkeGfkQNk79d8XYrlxid6Mc2IRG0lUYFMKtR481oTtV/0ZT5/gYOb
y7SrcgS4NhXYGMFRSuQ73hT3yXNjpidMb6NJ4CN/P/uVsCPcBCaSQmfAILNTwsF12zeG+Luf4uBL
r9fTELkwjnffM5xki1UROJLinwsFF9haMMHoPRzjH8oomu/5Nu5EkgJn6Q6UXffKdhu3gE36YJXv
uLmeBb5Q+/f5zS51nwZww0kJn12GkDC1GLiFYq6JqVUIaEUoflBp2QQMNHoyrsBIXigtnsdmUSUY
m3i471Ko0AFe4ou5mOJ2uDoReK2RyLyU+uLdf9Xd0Vs8Aj1fHlN1HrsPqj1q9+nk60c+M/PbVXbZ
VQO1roiIoYh/Y8VooWUd0/eD4y+Ojlni8uHiA+FpTVPQCxvuIWqBUsWcoGJIOmZdagq3ZBBlcHyr
I8D9o5Zn5cTBK1QJMTteVzHHAyfemf6GYVV2O6v6QRKaK4IJMDi0MEP+2wqfvFY6gPUrFOAedPui
EpbyF4QLsfGGObDIcMJl6Ra2V3JD2fIwKL25LhdQJAFAQjEYHsX/CWl/BH6nW+OoZbggVAKxqa4A
sMBkpMF5eb5NFEksBL8fUfYkt1hifzXhYR3AgdfbZRM5fQ+WHSue8AiBhUYBw26ySUFwA+xCt594
vQOeFxlyJ9/7VBVF9vB3TZIo/W4uoRL6ziFbM2IqdjQBWmjzkXmH2cHTHLtWjtET3rzH1ZPym/7L
/14DpyBMStRp3hphaQ4qWClfEn26IskkotbsC+de+GxBYfCBtfEW7w74W1ZlVLI68wDGGqUu2v/S
0/IrMD7fAvpzXAJPSDFwFwg8VWlgZSJxb5hk4nwA/nIhH1GP3aJjFHvg3rVuOWbeS9UAQC3otgbi
ZC3b0W67OsLAQ053+eR6gTbHSp/4sAyeVbxt2tyWuPdE0N2Njks+MCOGc8nMtHCJvTzUesHYWStU
XPWjZcf4ybU7mVQIxjgjDLF8PcGlKhme93KlPdRf3s3s/JKf2coWIGCjAkCgrqLbDpgpyYE5voFo
L+EzA6tWOmLikqKxW22U/0ePlpiQhu13Sw+ouiq/4TGROPtINJgndqhslEduECXMQ0pA+YqaRmEK
Hitg2q9ZdZrV0a0cadJ7HyCps300PIInv9MelzP94Pt7k2GeJNJ2DGbhSVknrHuPfNOvaMD9fGUF
XUg+HYAhzhrOscfhU5Yx9tizn9Rf6kDM3Ko01YFb2M2e8lXomn5Y01dYXfIyu6OBJ9ALIHL2e8VP
+IyI7Sg0j7pJcllilxUk+x+SpqlgdvVLeEUujudgodalty/8JOAs2OCdS4aa0GhYwFg4pjVbVnG7
8MvRdkjaf4JvHJBzCz2lCkMeRy0jIkhVpD8u8Ahy5XqnAE1nmO57rjtmhKtfnfscVrvqMSytw+NR
CnnLti2gCaU5MlFbYUXaMUCHKvpiEw1iZYadBSwiq4udkxo9DnUmS1J7GIMcHvLptYhx+ZyFrf/P
N26ydzZfQkIDPPgPIPLoMs4g8Ey7UV5WjdZyfsTA3JzYfhxKbK2HTxCu378YtcXtOIfxfXBrJ2oq
lpgbbXkpNaQiV/ilnE8kCeqklPkufMYsWqHRK1Ik84hN4iKWADJ21JlU+oTO2ZqZMbSft1KFZYmP
U8hd26+oJLakE2QDG9H/IXqi08d+ZaSSuqB11e56xx40Q3Wmdsi/RSTG5JbMMWt7UgJ4Bv6GgnAq
6A4eKBEsqlqwV9Fgf/qjw1zRAl+iOWRfnbzqMuzz9E/Y/cpIRM8NxPi98FlcXrj0Tg3PQu1yqvSW
JNV0vFMnEPHj55hcZmqrUeqd/fZ4qF5V4OV6pExrje84MkyIO/+aqyaD8UsfHd2tj7JUW+RV6HGY
ktIWce0NYS/C8ozy1964Gj2TtZNQ4qJALbLrpcjOxslSj8qwC4nF2dPW++KzTDapbx98hehyCYtE
24DxFYOYy+JWdLtu6LN3Fj05h9JxMMvg/nZNL2Y551D+VQgd+UOd+GBZUNkKEn7snZN57T+mIKTm
V5gATOO5qIhfjChl3Bqt6lyBacSrNn5SS+B+Ng/7+Gp3Acq3VAfD4vKms3pkl7uxowKpM6eLBGyB
ySZLqzbihFFcP4Hr1VdZ7Nw3Q58n4shx/6xUeNWTkWIelKyuRxO58hmOUpFjc8+O1A/I5yInMl6a
qg0gxxYUcYU1eSxNOKLNtpd51yJbSHsN5f4vqzc2PWnyOUBWIs6SCOdUx7cAoPTpVwgw0APfD3Jc
vOoINpwkfNvgfJpULrQuqZMRtg+72rz9TVpA9l8eULcLznV6mUXlCxpEBoxBw8+JNwV1aPPjMgfN
QMS/3T4b8Q9LQmnrI7sSFciLHnKHp7D4V7TQx0qrBoikIfaGs19ueW54kjozcjBlK1lKyNOp1DUQ
qYPYvNyrJUExOuCJOfIDHvrYqBsj+qaf16O3EgeDDSv24PQDV2+gCEXuB4w8vn+AE2Gg8eUtrSDF
Nb7iu2ITNsoqwXUtXVj62KCwTPWD6uTQEItGoN7b1dq8nZTRe23JYF/kZyqrYGihD5BWtEolbrgv
iLJVmfSEIdPvFLuQBshTiZWvtMHdFgDXu2/uDzoB26Ml+p6ASzw2Zf72QxTlAy84EhXHDh1sy0vC
JxcCFLkUU1Jaz5dPypvsdvkzL6p8xfgFhEDV63PGS4ahDsYJHO5yDpI70U1q/+JF9Azts14nyXqN
0TvEmpzaTBmjjr1iQw/LYP2gPUOJO0Tt+KebS++fyOMckf+87yrI53yOVSlrnss3zId7VOY8oFeK
mhoplI8swE+ba4R+j/37QuLFzTSEVTSCe4H15MYBLVQn6vEMSbtovvoRBVfS8rqDSPNaR9AOCCGt
4n+yDj4oEsrTh8+DkerhcM1DjXkDJyhoW4oIoBnKDIn0mnvA1fps6FnjMrcvaWy30DvdtabSnV2/
73hRWvR50VaL3qZloUfDynL4uNf12+H950WJlMjc7pWHdc0KRsm3tYyqw7q0y4lXqNzpoCBU0LSi
YCioKDkQVSToqPtjlhzXgqlcsMp30uiOw2SfZcnqkPg3f+vwwbZAhtRuZOpyqrJpnP31rgZVqCmz
uWx0mDTMZE7UwbJ1+k27hDVR8RsN7SWm6t0JqmEhW35t1+fxdmza28o6vr/NbyJzOGq8QED66Fgs
yjRgWY/DcZ3aJNfyv0xMJgNeoEk9bOjBQh7A6QKFjvR29Z9OoA2AJ3Kf0DCf2t5Gd6d22QG2HoAd
unxyuDV0+5BgO02aMCx5+JMNY5Q3UlJdjPmz3Mf1CfBZBmlMKV56n9d7IR5td3bXLaOYI2L8f287
/cY9VqKiXya8FZ7dg3W/Fbcar/JbkbPAnI8EXtxkdhbDhJiSChDcQkjNTopgytEO1kV/7tfC2lLp
YU0MnDEi78RGnKHO+MlAj16VxTzJastX3rCgjYs0jJdpUsv2EZdrcQfCzx89HSivE874vzAxeuCn
er/F/oUY/pyrMuW9V9vapAN0t0vtE9qFnnymOLlOH6A+XS+jISwsFDbF7d2ggPba7XX1bzwVfGTu
VZ9I8puDdEwyUqf3X3TWQU9ojJxYgPmdzBUNsYw+3M/zBYmI77ptiBKyx3A39r/SVrY2teYwS38H
ss7hsP4se/mfVfvpAt3WoHyD+gTLEgxK4oopPDmPKzL1vQGWse/dS+3DW3FqEZ/a3wEvnmaJ7KPe
06ASMhxcdZM1gP6ECe2ma/2nED134bR6Udd+wPr/nmFlbNmARxV1tjmsPciGwqli34zWLKGwFXmM
uFzkWPTPfJ1hqQye4cicf9E41gOB6VIal3lcZhStYdzkPP3iWkLVvI0BiPPJzo6Te4MPJELdCcwy
rXCPifyxlYMKYIC1qlkC4WpeDV+11qu1DQoG8nGWGNCe9CFQHbcweaY4U/5BNNQRrs3UpXYzOqst
nXAbeBpbDM0YKv5PmjBSP17AJYtHdP4PQb0BdcG1q+Gi9qGnd1jbnGgfk88DxCr/K7+sFu5Hb2zw
nckICjtQ6wS2ajnAFTVlBlCP3S4EW7UquZ3ZMVj9IN2U3yCOuWmQ75Cs1bTDNBdSdFoF4dgYtPcH
uVjLluNtCp/fR8s2RDm1LT2gcQc2N4Yscr2ElHxQ3AaGjYwYTG7oL9jGNX+tQPowZwFmQFBAqnuf
e+FrWI7rOIQbgARoi8uqNe8HZAfOrUIUeX7sZoGGm9z5msVspMk6BLkftJefjGERoebZO+yquIZF
GayYU0NvZpL1ZXvX2uhIZhVvPtbjg2J9wCXiK78eexKLkfH3vB6O9udscFuz6+F4Hm6COADNfZoc
8Ghe+z/JXrXNvCB+d9c7sqxlXzl6okivo8EidyqxQVk76dmtdtyhgFgVKOlTkdA7/F9iRfSHPshU
IfyZ9A0s9DBccUvHOat4v/oRmv12Y5s/0+Gc3FR2rcuRBqOQ3WfOF6sHSlOjmUR4LrACs9AW8oqR
jl8S7DweQV0ZjaVU+S7RC4grT4ck+hdwx2hizhVe2UqYtiGxdUA7M2/BoOs2w6eEbUaxvfTiIfCO
AjFO3XQJqnbr4szVEySBK9vlwmXuizn51XBEPweku925E/VpOTVNVbgr875NiudI6GHGV/laxNMp
isrzTPAxAy5IN+refllfw6FS5E78SMI28VpFdTSG3V9aO243SbVXeRXBVEYg4mBBqMwyvQjjx3Vq
35IWpOEYcVG/LAKybsoAPMEMOG0HopczT9PmFdrSR/pFbH/i1nRY8OOdQNHC5b1+X9GN+WYUzZdj
RYdeQefdFqm43fLjDWHdZf+Rjw6sCxYwpdeiICxOXiVo6qzqz+OomA1AvhmO8Uu76oEdcTILDq55
p0g8l3Klzqrgik36SoZgiVUWCHkLtSNgXKlFjQc150ZVT707GlOpiGfE0cdaaY0UV40/kkbz48fO
EUd/b8AzhY60Yeaph/rnPqGarkIEHZwWL4B+7bRol7vEBLTulWS2+XJBOl3lz18Jh7/04yZ54gYJ
nFUC7z9VAX5LkvKSGJW4cFiLBLCzGpKKkY4OjrSb6BCgIsOzPrYz/rNDJmVbQMT0fpptF7iJ1+YO
yyMNHd8YYnkzI4jBwHXDsIGlze1AG/g7suEOT02wFgJ/HGzlRExQegkOKDRNGCa4UnZbAWPVJz4m
q9i4nc2TcrETZLCstLKCFYokCjQLpMKjrmTiJA/q49VNwlOUEMypz2ZzWLLlR9vbEJzn/cNcTn17
CBRLAyLE1CFKVZu7fMDtzKn2ZsIzN5KOvR5Ms9lTxGywIzsRU3iV1odAxQQ9Oy+dyJWlcf94Nhuk
yEPB0nbrhu612zweRV+Ojht9hC84SnrKkDu6OdJLxlrLXxKAWJSDRyu0aS27v7ysEBLV0w3PM7sg
gGMbkFZ7N96/qwG5lkl4FZseZBbMv5qnmM+U3PukxbOufjoQZ+ynwnXMig7EhvEOuI1nkWarbUGg
bkR7uxfXkvzQRqC2RcTvo/treDxPXIZTLGI36VgIBcIuwC7OFoSjMn45IZX3bKlApIjCub606/9p
SDT28NVy+PCTVYKUK37sgbocmtFnszGkZXuWv3YbJ+MQOreQXRIJGshn18ATR3mi4ovgE6amTj3m
8AyUnptJ4wFR+uGm5wPliQhfl/wk8A4Scgqu8XXMdn51r/xPOuwyyoDfNPpR5fL5f1FE/tQNcImY
OGzzqrbOJ6dn1tunlS52hW1+3WMz6+eHhK79Gt5dOU2wGiTPp7XlvzpsKnBZkwZJ33uC2lHkZLXe
/oYndcvDnN6gNwHDv6yFmbbSuuodYIjk/AAxoOu7YHCAx8TR+DcwaW1q/h+31i3PPDHc7lAK+9Iz
SoqTGO+4J9rWTX0iUYAxZovOGT2So1KwnXhqPPsokAhVO8mK6PgiR/Rywdy9u4DUKhNKAKwcPTS5
Uf3EnkALaXv7VQ5Se+KRLR+ASyf/8AAcbY1tXSNKUii2385UEO1Njq/bi3Tt/ZjwTHx+wfeHkV6S
I5H/bZLRaZ9VPoQY34a+pJZs2IRwg2fm7wb/PmZ6OwYO5xH5neSIILQGBWbCLwdGlT3Ab+kcWK5y
uAzroVtQngu4V+0BNASmi4cw/StTENuaGCdX/wwql/mCyPvlINaryw/tgcEgE8xujUPwYK8b6Fx8
W0L8uO1G0VjU5nGRXB3imDau6/IbzBWCH33HNq/UN2cL/1rEJKHFB/JoMbzCLY6vXjRLTNz2emZM
l/6Oaqao58fAol5fayLJMb2IVvWv61KBPlt2JxvuqRB+kw+SykegBrEWw4/Tfs3CqfJgE9YOTc18
lNyXNGVD/K2McEtxAAQLsv1FX5bQR4nAaIUinJCikx2owRHwnejA+ZNwGu6Xj1fRvL5aV/nz1CMh
Ksr8KlNZ5Wfqj3v5fyaLeel2ns51yBYFTXRQWWgX2eOUGwTXk8p3gUzT7Zi24xLO0TcCyUPAbdZy
j5WhsQv0BTwu/6+X1dhv6RMj2+se420RHbMG7deu7bFCvqrIQT1VAQugbk5xrxZ1h0ihZ9gpsxgT
P5iEOx2bUgPjkwwadNrHMSjCIu+JfEsZ1k9pVoOU6izGk9Zto+K75n4tzmGOwQzWE2YR50bfe+VA
xBqeQ7F/BQc3hkcxSRERZCYAKi8BFJl4Io4z4JhVVkjhU+PQ8MDYXBUzH0e+7YGpX9UIRfF2jGmL
2F9jkMyztyO8SFe575DgnONyLJGHWXVuAKXFPu2D+epyOIqsYXDh5Q3ByxW2ULWkuzkfoArUbJvw
IjUsTXpiAIeRoGTE1Nz/LE6+u22l7texxGgDGqi+tLPP+j053sMyJw/0ZrbARMvb2rNiEN/dYtVP
O5+ILtuZZS92raOd0V/0SbyAJxCowt8AUJKJluWJBilmrgzzroFX5vGoGUHgI7RSqg7QIpo/F6B0
9+5Kl6cGtZOdI27QXiXZPxiISIh/Oxa1wo7GAT9nVAL/gsv8OgQuWKI7pXqi0jgYlDngM0whUlNH
snacsTdY9Jg4MEOY9jIDc6kFOsoI3PHHod0QAagEfBjR2K6D7/ur6kDU1enISgrjFGFwC+UvX0Bo
dC+S4Eold8jnZtO70atvsxjAIW7/Hd3nd530YiQw+xgfEiw+ia0MufJj9tDXf3zkdvDWDqOJZiUD
Cp77KMYeQ8pxyTckwFMyarlc/3oP4lSToGWBWMf1oraQKtSuuPxvuywVP6XmS0TMqY3LpvQxsKry
EIBx1XoLWqbgcfL2yooq9YEVnubrRTtGlj6rvvE5T+X9n9fCb4iwntCo4wv/bhk3wnm6F/s9Idie
SzvceAqyWahiMGFIkCGITTQL7cL0ORLOHGEaOI+i9ixHeOqm6JprQNCoefa7LsG9JP/GQdYz0QSO
b1QHHOJ0kYTb5D2GZskzQoFKU2aknzlSyxPb9faU5Bwo/k0i2xHF+rqfjKPyiEDe82WIcbQSYJVD
C1XdJPEYVX8QLi7LMzVMbORHJsZ70kbD2LUgNYcMdDLD3unJwa+DZCDjF1inb1RSbIhs4sqzq3oR
T7eFt3k84Vs6yqvVjvBheH0VQ/Y9GFna+1hSjdQ1vj/xX17Y3qblTdL2Fo9SjaHt9br/fCNOvHDB
n1n/lB+UD59KMKomYaCG/GVSFWkaPFphqUawhbrkrDbk8nuPkXaKVR5BoPv/LMUgOjhPwuM5jMAA
MeRr2nrRwpyi+FppS28ZtTfBeM05wnMNXuSiia/CR7pkL1DUlQ2XNk52g4ahk7uCHSYVxJFoSp5h
ODGlDbOQbEYz/RrDjztX0YPXKBJN5HY/kbyXbntVKLDrLK7ZNrGB3GuB9QI7rixkKDpDRDE8xLDH
gLRJOyXXrPXRHpABVMJLfmK60lfzUGtFxenaccp4ghcd9qWy0zuTxcpI0CnU8aMkYduKdpqb57ri
D5krir41F0t7ND0oZyOJbKgGeef/loqm7jRr/bfSGUcxCtwL/dxufrrTbJxrPasXaeo0ZdR8nvFJ
vXva/JQPAmm+bfHZH7Ps8Ctp08obEi9HCqaQUPWPD+e1NvGQD3p+xjqBRHK35Q4WpLEif6lhz+7K
FThu/CRLwcFPvDNH0NDvKWz4mRv7tG6R1iofkAAv0kPQxtIsEa9SCsocja3Keh1YWKaLyJA+fE8k
fyl+X4bYS07SgpTjDj/x/egUz0YzhcVpbPLukpyrag4iQpnurSs2ZpRMwEBqelNLL3KoDNSqm0as
3dTJzPkNvB5Iyf4LsMCgMSny+iR/ODxMdevUXyfKbr5EFYq7oxU5jCjokOM1QK/3THoVIbrsElye
qQ1MuFqC3dRbS0+IO61a44hTuvEM5qLevChHQareOZV0pOw3J0iFmyg9/POGVGk2Y9TdxB11EJSG
pJ6cH3QnoBH4hTa+QlwiHpq8mfPfJP5LWddKRZKZq+PJInU4NxnfxcBUBPVZrriVkorHKc9f5xVn
oEZYJRbbq3XCFqGPJvTvSJotn8UeBkjN8eyYepGFuwZswtXtJYniB7pG6chi8/lzfOMnDXkiBLQd
LzmEBT7+eRvC393dy0Ksel7CV66RFVWOsS8ARfuosgHEbQz448QDiFUT/1JJmYzhSNUqMvkDgqO+
oO83s3C6jjccuZpVtdTv5ZWytM49RazvMAJOWLEDENbzVTLkwEQuHProcX/mIHX8JEENoqe8Wjv6
Yfu7+ozu6v/E+1rq30yhKJEhAJaAq863MVdDI4xB+uyI5NdwVKQtUhf5Wel1QIcjbe0X9cb1o0Aq
CxTnyZFh+zngUxQXLwTWtAnwsuGQEToG0jlMakRQ+XEoKEJ6EXRrlLNaURfkQ4VMdSjhf1Ydv/mU
el09D64W0qNdZe1x6EX96HIMzEOKFsJIJFaAki43mkxUKYLGuVb++0sIBeIFkz8mdCralEn5IHnq
3KMDTz17gWqAneMylc2JXByQcWMbGLXYiFmw0KWysrAMNt5pJJGBmNO2J61vY/qj9MfrUdpYHMp4
iShba7jLL7vZ5G7kz4IhfqvD5AzSb4YZpovpKN2JNRr8Ex771DqO+H1IoYDxuMmtj5swBxv9QFKu
8h/0/E9LjV5uNU/+7nUoVxOgIbio6OQhIMCi9kVmljQEdW0UhdNO5xBaTLZbICzQ+l/MyuLitj1U
alFRM5gSn0Dg7MkOx1lahYX0MDaiWrkGFvjDe0RhoLLGwnBb7KezYAgTOckLnIhqqroRGwqnWiWl
CTAB4bvJXPvoXccVIoG4Lsk/hbYfJK7t68niqqh0TsNal5twxE2C1p+aIorfPCoB0VZdVqTB/faK
hN9KSfe9T2c4A7XzQhNAYVKnsrXB5m5RzL3U/5VT7CZ/CAzzWBTwG9TTjcPVCE3Mh6PadGDjRxMJ
bG49PffALQQFmzhNfK9/QOL9sgEsFrcwiTj1nCvafuG7odvPzLB9OsS8KTg9YEWrybTVewPtrJvZ
WwfMAeYyRpczHaYb6i2Kftbycb+NLJkca3XAuJke+/u2NGqh6+gqpmTMZRiOkQSXWjCF5YuffI1U
F6kctk0hcFATXTeHzwJ7lNKSn8ZNz5X/T7TStYJANgM7/j8C2pc8NnZ+yyq0NSu+qTOJltZgpd4N
srzD9xBgt2LXGdbEJiLExpYkUhwdIwSDIxBRU9G6i9uiGw3+tv8crFpTzDz6Otc6fpPfppRntvHN
vL/hwVFcWOAAimr9kuB7T12f85vPlYcqYpK9s9DDLdRvVEHkLH8cxstWmhNiNIQy7bxw5r0GTmIN
7+0RWyn/o94yAP3OIyUf3xRvFwchO+1DQAG8aLlPNw0bmnliL8tFlo9f1FNnzVOFY6GzjGQc6/iL
XnXsPGynaYqoi2iWl1vEPVtQ5A/Q3VN4tgwO2yJn5at3t0F0KzlLiiwB08jT4JVbjfejgR819j6O
d14Y3a23kjRezbf9letUf1028x7xzul7/hvBC4jHqaMe5IlIwjKCjqXM6mPGM3ncEOBEJM79p3N/
6VTgvecSAOm7DznKVFLKGfskYiX/3EO77PotyHH7EPP8FTtaM8qTijFBM/kZfh6yYLc4CzPZ3Tsd
VAKqrpw8JBAJP3KsifwuaGw3REBjnn2R2pXNqPeSilGTZtqZjBoWPqUuvcvjq79CmfD6w+MJd1rD
ptzOcD0hAXEQZtfx6c4R1yMdAQP1jWKdW3/gusjVYV/+EOc0o8fHVeKCk929GPci7jOTAe9B2md1
mvieo+glEeZPbLIamKebuux2czc8tgX53We86uIsykrCcbG621sDaWM4EHyaOJ86e0VAYbUF+3Bm
ncoM4CqMYsNdJdVczsT9RchsmgiKLEam+0Bt5nayDtoaZpllZ9P49/dtCWrB63OFAA2qBAz3nxyw
jlmM7k0XfKIGANVK4bUoHl4xBIpZUMPztte3cbHevfPv2yXGvIoH9cUTMq0IQqYg26EmWDY9YuAU
fUnzdoJHg6fKxNsyklkUUqMo2CKhduuCamR5tbrFTkQhC2lrmPVj9Ptc3M6fhomx+AriPJbuB051
x18RRMJiG4UZcfZwgBMNhxhW2q1ePdtb2H0rxSI4ZmEfBxh+X3rx/54iAPtTkHmj8idfTia+ql77
iLnsY/WY4S5nSV+NgcycHmfU0v6PBzmNI+I3S4DsPAjf6DZCd3Jn2ZSWiny/HjqYKilZ98NfYwgy
wrcic9wx7kMcRxRk46Ir9M+iSeH5szkh3kSkraM1qd3WSMMmr+2ozZKrXD/Vk3bTN/S2MFOVzOGM
0D+ZZW9iXOAkN6mfvIt+ExWcoRU2/AcV38SZLJNVqSfgEZVKsWBxnVF/YhWd4iFpxa8V9pn/J0Ar
u7dd3t4p2bywqq13qXtzr6+GHgqyUuvvRX7MmnvCQVkOLS33mnhySt+yBY8A1CLz1ls1CJRfm7Bs
HjKidd4sEF7Te2IifcGqr2sudf8v2BxxFxnrs0s9pcbpYiUMJPuKJiCcqT0A5ibJ7yJQ2EATDEbX
7cYP/Vmwa673Euf2qdmRHdC/hpaawhUqK+bsxGvVccnpe/6fHSPQj5lg60fnfJVFtCcG/jT7ChfR
jPF6TNTRZOQrpVWZQKZSwPSrRjGYYOxxP8qXtWzfiv0LstdftbT6tO5JkcTMI/AiOx9Z4Fa72nG3
Dheqfj6f1YzjqE4oCRdJQaBx7y5Twgn/zvhxQoHV5FpbRoVgjqmgsFul4C7+naQzDZzuU6oLwIyu
cy51eib5FC5AO37wkOdqxSLX/6A/mJ0Bb8GUFvWr7zShX1aYtTSexCJI2B4zdU/mpDHexg7U7x3o
LFHDJcndWQem8aJPL58eG/x5TYiXJ5CNNHJf4jMMH1bpOQyBDMpQyj+kffwU6SuHHoe9Mglk7MyF
IKq2pT8Tx0Np6VKoWsHI505kQp6xfFwdweMYJ42VPWJxjhTHzOyXfbm4IKXgpRTFDssL+h7taLhz
negBFwpYBXH4D6J4XdCZ9YyQyfIwIvmSSoKOhiN+iBEUK1Nsrj+izwRYu6fMrDB4Old1CJlYeRbO
bfixe923McYsb0QKlFW4WRfGQqqnynf2sVhIItgDe7vRJ/3HfRmcF1nPnDTYSLeSx8hX+4puQ93p
vZGwc1T/5cUYxaceX+RV6fPUoeW7yvuKjv8I2mBvmLV3ktrpr1oYcBXEZEMVDzSsRNaT7lROWYT4
PJQtW5Ra9xSKRcs+FEMvCbQGbg4uiX9xKU1EHJJH9QroVoggmHIFbASm/Vb0Wm3yIhEfr3kGsD2g
2w6tq29pQMlwDd0ikUShifJI0z/7GjEEVucSPLWNH1dbn1Dih0pC5OTTof7CbUXD04jqtmLR4Uj+
uaLZdMPKOdjhzvUR+LC8HVNzPFNOj1JWZWy7kX1iUqtPh8SqE6Lf5farjVvf89IFdaT0xyRumFdG
EE2wx5/jXoIWTINVsfbTX0rYZjsb15jW+GtJpLWBQXtqt4NuvCqMxAHt545+qv4vK65fjfMY4K/u
i8XqZ1fMcf1BFzTJL37T0gaTQLZCxmz+DqcyGHhdg7JVF5k6/mAozKSZ4qIBw/8q3w3pMKlMXpVN
RnqV7Q34O0vivSz+HcbYxIAB6NcJ+UhAccpEJ016d3sxjMML4fZqXLt/fQL/Swfe775C/twcleZp
liJnLtMsQqtN/wwxN8GDvYIXecSjHiO33Eqerz2kQxqwze/otFnNLPb6uu0h8CnO2ybcKqEO+0Ns
7HHtc2sSvGMVBbnMroJCGfttjPDy5aL5BRk0uoE4WDhuG3/vcnxHImiNiNk25T/bqviPd5dLnbry
Rp7EpgTcDO4Z5LGmaNUwHBEUhFU9CAu56dTgQURI9rJHaEMMgE6l2fwhazaois5BWs9ZabLSfzaZ
XkqLLpsKLzTUWUyvEaqLInWUoUlwIbV1/u7soE2bbxxBK2xHzy2WoNeT+3/4P3cI8LByZiI2fGgE
/liPNeC0P/bKqM/VccFB3dtnb15Fslzatk0OjE3+ew/tNB4u7uDJza/tFZfR/fi6qtklpB300dEZ
2TjgeAK79300lRWnqms3R00v2ZZthuINsP0ojHL336isjc2s4YmRtukxwsmUBG+5f0LspFmfdM5f
kGHqIudgK9tc2A7sL/Y/ND8yJhLv9xzZ7C4fZ3ruO7ZAVcbCzZPRoZR8oRjYshSYWngYbfvXDxPQ
An/pwEXZLI/95M5AkYqI60DbF58bLzo7lJ4UxklzwhAG2ucxSo5iFtwKMYnF29FclE/XIcRqW16D
nzuDJDiSMw+L5BR7GFBSndnQ+1NTVbIYkZ5eAu6OgSFFjsRt7f7CcFV9UZj+0go0YiQk9te02AfI
BPTuylrkUWTY0Ec37Jao3oAeFXPO5eupkAM12nLAGNQtNCO7yVJU2uOeZ+6Vp9SgyqGCa/Ss4csT
WxA57ABUiuhTfNiidLwrQ24DvI2N9eTbLUfZoC9PEBZFw0BTs6ckZi51/CKtbsUZFtgCjH8YOKld
htv/ytrQngCJM6ivSDT3aOBU3k/0vb1jIfCjbQez1/98fp/UNMc3eXsTkWt3LcCB6VfVDs4gL+fG
qc+VjseRbOw24uvOqZaGKX10JArjtiXSC+KbqZ2xFq/oaFzlxONHq286eQMfclxwxLbJslfCruU1
LmLBSK7Efxwm+/cS9DaefNSGrp9yT52W3fJBig8wmuY9FZMr9i74JqhadBnPEtS1QxKKuUmpyHTL
9ddUB5IHqH+ORm5VLyPQNeWuQKr/oppDpQVDjxQaVT6HP7LeKy6XK1BRRgwVdOQv6z43NZKbCzsi
BUL9udpO0f6iWGtj1iGovp5ESEzcwgVH5J6ZMs9WUa1dPzjF3CHLZ3rw2v+FT5LUrO6O3fKCAVYH
m0XoZdd5VnbLCk7mEY/Y9tbWAOe7inZKbmE7UkxdCd8fqJcSTpgmhQCes4av9mVaS5mysbcqSI35
i++yLi2D0tFfbGzeTTUhzgH/Y47HpWWXmcqMgb/wT+pxcUBxh554uTVVNFKhAsd/uHx+2kvYYhxp
npn9ikoLr3tPDDi38lm55xbGwNG2omX5iy2VIuyoXMCssMVHwerJG/5R1BeQBgsSb6M6ykFbayvv
+wa2Btg60Eejwfpl+o909iuONewTl5vYou1ZNbv74ABdYb1AssySk+93asSFcgMFyd7joEjTEAFe
2ivisO7o7JX8cDbZvujpIP80mJ6fW/qLkf2XtpjhPJwjGOEXufyvluXE/TAZSwbGiQ98K2xYr/UX
e44GOntMwkbpTotxHAMs57uZxuo70AZmi7fkveNJri1HW/BIn6ke0WIRNudhXH/Jg9uHc9P9tB7k
LmvQkyEHIe4tNsVBEUsbF3i1wRbSINTTR9x8/do14xDYnyvesbQ9o77D1QUYhIqStp7erMgSnpGz
Zccv7o8HxpVFOR2aK61Ux0AOHNC6A0YX3gK+idwiWh9fgXkiBpwbc/3I30/PZa8VAkko6VrpIf9A
qYkpvBaUs7KJfeWXLp6AJ5MK4eeXELBJPyUcxyHjKDYrpL41CGSJHGceroJZscKo9F1y+xmIetHJ
m15puN/RrZvpqFyu4m45d1Sw8xg60RJ7TKP6A//NffeyOVeymQXUREKdX+/GA7xdggvNYdYIJW6k
X432ekxF8qNv9njN82K/CDJa9qfII4qCi9CVkasVYFTxSBr3CPJVrVsCd6TinoYWe4FO4sC7TwAM
hDzNiOF+mGQmE/oUmeje7Rtxdk+bigbC7T1JV+aQvDtUUPQeqGuS5LI8L4kdN7GMje5EoUGhFqWU
2mepW1iDvtG0oC0ILh48ph7nZWcTYhC8w5s3IE+lLe5QpHBaJWGeBNjfgywx8dKt4mYBQ5yn5GrS
kg4k/DYRlEq8BdxWksP3eCZ1stchJ3uj5S0yV7eAE3gEW9VoxHJSduoQoORaREDKzkh/3PEbdKUu
r7OsJMovePI76/EUTNj3Bv0Rxi7mHnNvaW5RUxyRy1Kbe5Q11u2cjGDEd+DOJ2JomIytMq+3IBjL
SuAMjg+hwStDj7fDAXcr/dgB+q6sV5bpq8YO09gHMQTzBOGQoOGg928eGtFHRd1ohWpJb1DJC+Ht
AkSUMNkIkTt9kCDKsMSb9JgnHjCcKIUgXBEBm1wCCulSsZazDQkOM2G1ar4uzW0P6qX7oTe0apaJ
GghlH10Ugf0cVQK36cdqrDK5EZ2lWshfc/LZqVT5GbUTTRpZWauaSyjrVXfQ8YX9RJM6j4uMyIUv
rtaPxlIb8uM2M3tAt714Xpluztdyao55W8HhV+h3Gqb7on6d0L7m0RJlGBbKmxw/g5bz9Mx7IQxu
0mAa2WyJ2NRirjOaZUTzLJY4YECXry9u1abfMUusyhigMOkmrVEa3Y82wcYc5BYA8pNIw++eijJ6
S/1y8PDlwjmNW1twiEL7rfmQChVDPJ9X306eucChvdtfmqCBq9hpraRCFHL2Wy8WCO9FC2QxAyfc
fG0AIf0+HA0Lcn3nRZPQ73vhgndrb+0Vj6MwV1+ybHCPn9E705OXsOsL9505ZAskkO5qzQP+u96c
CxDAkDsU+mHbOoDkYtKADhHMdsvsl3dB9D/cAkk8QZBxvBsq2KktVOXbzlXBSVviEF7g6w8KQfKl
mTaQZe2NpNHQYwBRpNEv4oH3iJdeyYSDTq2v2xy8bNgjW0mmP+rbj/5uCkf1lxt2FYCF5vw3cKPF
8SyTYwVHCyGMAZnZ/NQvTiBYC5TwF4V1hnlRM5ujFMm3diJ5uw6Efd1k94DTwvoO6hpDqNdN/fsa
U+RDBeT7nZnxTyi86CB0+CY01RfQWxF5kv++K9PZ+6vwL2v9pZqoEWAhetGoWRwg+TqtzBTqIW/s
BZAneosB6OOPtg45rYW+Z3nQVuYsRgsPjiFs38qtGkh7MHkZXT756Ds3dcsYdGkEGVUNWQIjl/Vh
Khooqz0QTK3npfHC6yoy0fK5QQSJH7DL6BMxupC0KU+BNG2vooUR3/oZgpdgJ2bKE3f8fJNGe2bM
aJ1sj8rM7YNpzylnCGkP/KkOnuPN/tQ8JtdCZcQ2jP/CTsYgTONRw5+5Eq5I70G0iB3QCokWwidw
iQf5Fe9TFW1V6xispypzDzw7eHMLTW8GPgDTgGtL7ht/dPwu5JbhoBZ2owlxncQ5THf4GHP5ivhd
eu5+Pupb0ZapBbhg6EVHHuJktJWSNiQbdRJ5zh30Qah0mLQI+uN12WUfPV1KwgrqP7Py2TRL0uGU
OgOQNFWPMW7guDHxvdRB60Y4Qi/881arI7KOdo1uWUkVBUwGv3TmYHBoavwzfTjJuLfhZMO5nGcu
PH3ck3Q1Ft1OnNTjCqVprcNQacgxOZdLwSTxdrEx3mdwjhGLBp7qvnofNbqTZ61c0nfB9f4diO9D
Ua1rlObidnUUYZTI3TBKeYpIg89dUSR4YeYIWmVA6nFZ0cAKH04M8mbxc4v5Oc9dg0+F/Sf9q9Uz
GqpH5Hv2RFw24UUbXZL6LiZuGI364tJJDm8TNpyc2uiEz66FhuYRBXtvID7v2qQyfN2VrZHwhTMj
fltJRpGZTer1hdb7w5ZtiKAxI5Wlh+hVIYS9jrIP7CJ8odUG51O/0PDTOKPWesUOSg8BImlyMZ7d
gacmGOlxVsCS5mmmBOBmAzydVMrGnVs1lPa/JWGa//9AtViHk2w3Z1205t8W346vA5QXKNNxGuEq
yMvsdoS7fDnmG1J3uZ50KUq0t9G0cSEFKaCsp1heMYDohCaIJGKUhXcbyahdnG6E6qVlm5bmHgpf
tUgbPBeTtQ9m5Wx/HF9xlYG02a+ai9UFcu2A/44e2oqsRfg2ingRUxsFWwdsKhwdiEVlVPj/hRuC
Rcn7GKWuEcuvH5kh1Z5DgCASzlqhARH5JETyZO6B8JN+0f2XUU3dcrUXvmcHlU8UcSGyCu3ulZeo
Q9w+lPX7EL7w5iBtQVhGuN5goSwHLJFa7wrd97rvcJt7L3y6XiJ92/hzRQqANw8UG5BDZbiVv90x
r43ckjnEnq3YQqtVKNjQHawF8z22Ak3Qp0bvPEu8i889ZrUDDZq8Y3gO0Qa/iu84uVxuhFbptquR
h+V6lH/B1Z0VruDgritH2132lsfBs5NXo1i5DL5W5UGD3LsVW6ko6dgiiHaaK2XsTxSN0S1nsAQ3
z2gM9+bhjQQ1woI65h6yv9Z03UNfcqNmGdGhnpw/wa4aKWv2H6mELC6h3vXKdA6vn0cA0jHk4K30
5quKJRR2NXSuginztOk0odWpvfGbngpM/aZdKzn/gQmq+XA3hlIg8KqPEUQd+DkvqQ4GiolX13p7
xwnD4UlH0dRlCPaNG8LqrOz45WHkRNfN3KuGeWildZW5Ygkw9GR/00oQ4LeQNtbIzVSvIed6ZFNT
hVkE+CcYP+JrujQb5QbXCxCK3rmWYTfZ1gcVuFbow0ITzcQ8tPLW+nsMTgW0EkjGuj5Suwreyw5Q
vI3B+RgGCf98io/F1hAH9uogKD7l8NZnonpzrXbhsUl29L4w2pR9iiYZPXXfxA0cPJJB+IUwc9yf
40Y5L2UJWheeROBIR1EG68OWe0s8mLXmqouUwodkMKQakxgPrBEcItJ2c54txI0AUvXGT2d2WAr5
KA9zYgC5HuB2lhRwXi3Y0w0+4+5ZGfUv85LUkjuMf4Wk33EIZW8zhI2qW4OLuMJebDc0JiVGQlMP
c7RUwzTokaEKrdDChAowLIl4EoRE72OHIb1z23IKvSt9hY9I2uE2o7AwJ81Jyv9bon5Y4nHyuRPx
Py6t4zQp+eIz6VqDyigTzsfCQ/SYp3cbdJyZHbnG4hzTt7nE748md7YRsYKjSG3B6pF/synln7Zr
PS7/qBpEX0RXB3czQxoZ5bqT6aNDfDJAf7VcF+h4hqC/Sy20qGH0V7wMuKLeFVim8bDS/qcyxyta
F61s7Wnz5WY7xMzAB6caBd3j6lf35PdtrwMgGbD+v2yg5t1tzg6z8DjRsYgvYhE4OrUnA3BdRF85
7KC4nU8ybUcvFqq3DyVtU2l2welE4CT7yq8PR628UHKxBkgjzkJH3FEmgh8cfIhSkeG/Y6LcOlPs
VUBzeUmGsk49mohwCCSJjAYVl4wKKX1B5sW/WFs/FWmNP64soicHl+EhXE4O9S/pVyaHDNulKXk4
/bQsN24RgTXZnbrRwbMnZvBOEIA+lDONbJxToPNzsiXUKaRdncjoegAcw0Fh0g2DQ1cClo+r5PZ5
Un4JBcvPrLYQIzy/rFvEelgP9TZroPAwxv4h3cD+pKQYbUTP1MNhTKyEFRRwGdQlWQAWE3N4SA4k
JqzCK3uFYrsZfOpEylyc5fREUaVb/NRRQjyEoGpEnv34Uk74WWp/Siqr31QxmBFOfEflzCBL9pWu
3juYWsQyHsP/BPXySlpPu8Wtvz2MvGs6lqAD9iBMGLNQQKYvt7W/PcQJNl0s9RSuWO7xlu0MUQDU
NW9JqyYMY6QVxaptVdHo1cwCBmi2jh7+fJI+57PYvV/Yf10H/8so/3ZailmUPMYgbtjPsE22zk7G
TH5YEhb063QoHbjNfh+PTy1W8zbeJQ0BE5afI/GzfolLChGMhby7QD+xfpyOVi6mz3oJj5vd5Zcn
E7fMrXkdg0WpenZeZFcQxUbzYRWRmH50MjQPesXdiFvjlbEhA9O9RnZuYfjNb7uXUe7AV1L6xPDR
otZsQEIQ6x/gZeqlzCfBf4Qs5cQwCv/d/i63eysRwJZS6sxypAN7fhp/T7JGTRDcHF2awADM7F79
3OKV2ZDvRbJIf57dhhcOocFIFJ65NOTuyj4zGwAyi5yIsR4thVDLRv+nxvORqcQZIyMGD26rmCcv
TkGjsb7K3xk8aBtlHr1xXQvTvRtWgaRfgtbwG5iFJcN64MaUT7HnkcMEQFlBdPpy2O7XOSVuVi3g
inA0C515JHSlssxKoN4A5bGL5hfc7aQYLBfO/ahfdVZ4IqPJdhUrIWLhhzVuGOHR9yTUuhir2Z72
+l+e8gHTKFgfFhA2ZfRm8aEkBKfU5VW67U771jDJUVAWsPOqOcnD+zQb6EBNjYYWMzrU9/choj+1
KpB82FFrKqTAQr5vwUS50tXJjBUUVw3HNLtwy52Ar3UkUOc60rx/JwN5EvcG3wByJt34pre3+zlS
fEsxHy+8qRxIxT/6wfDlzHPWM6QesHbbDb7pRxR5N1x8cvp6JpveW366DAUBKl2idDuQOIsl5VDM
gHnyID+OV2bEKgXUX5HmRPj+x9l5abMHvC9oN92o6+QlbBTuCDWDuvlG700rUADVKvH/QE6vwY7S
88h3ctsf76C1s+samKXOXvVZ2m/6P7JCQ+yhVGZLrLD8H/2zUNyQw+KImY3RLEhu5qF2V0s89PmQ
abT1AQMk/GOzNmS8S6CdKbc0VWq906JnHTtVjz58Soq94xcWTHXpwzw46UiliizRzb8VnmM6rWxR
9HU+cpSCvYhsxszZ8DMVL+2d2Ah33vRXh4k/WaeSGza3l/NuCHobhrCRNsOvOtBM1mMy7RYzivMh
XyKnoOyK6vnPaqaWZOZ4zl5oZtDl9IseYHdejkycpwnOwF0yvNobUEyFN6SOMKPjUhqlAlYlFLS/
J42qrvBeN5aoDpXQfd1ceG1ctjsG+s6sKaEWdI6LxTgsxzxSBAaLQ2F7h6NiGgI38JkTTGQ3FHHN
tT+ZE1W/gK8PvaQkHQXEcRrF2HCSV9gPmE+NK+qU62Qg84eqhwKkamWovlKg3q4AChQqg2bdneSm
adJBAOFm8wj2JL+GW5UKBzld5ukf1rjeP91K6GO8y871YHg5hpQnuU4oHVUmZvfPHLDZRCA4eHWk
tWwJF++Alf0dEwPVIAT/91KVLbdZhNafhzhUczm0E7EDbocbjDVp2Ms9o80O2ZNsLZiN1nAPl/mO
WIXexXRHbbRYVkyGIR71g/htMEkbp4K0wLoPAVqoMhy+h4pfneuxoFwBwQWIFt/FpAiQWYnAiAx8
eqT0C6zQRsa9+/VazcfWxtaVQ5/BWzNAaleEGHEHQhj+mJmzmYf2ouK1IHVernejoeMNvc8h4l6r
xxdlDJO4ktcYr2JiWQQGKuKM/NfTI/R+FZqYTHKkn4tQH7XfWZ/BvaAZ2XRMkbUkOT80vNVEcLY7
5KMtIQaXETc1J0lx1RfP3dFvupx22TT+ac47mDvQwPXn7t0EceBfgZAaGamu/SUqH2Qla1IAduvq
UqW3bW3Q6Xbya/MEeSe9K5oDb97ODAvnaHel/lYRpzuanglKoPV6wK36PyM6T8urDXGDyAJVf2yS
D+GyhJGEsMzY1R4/H04Ka+imlUrMOoSf4Ur78ZDTNovCvSOXEzvQ6avVhVRJ1S8h+iuBJcmXWA9H
RjykEymHQwu2jNHp9LzjW9yy7QKLO/Ym3qOP2Xit0sdhiguHsEMOIj/0Qt/S7Pwbgq5sABrRyasO
jd8QX2vxvk3XV0ixAxmTvYj0mrTYEyUdUnBbzDNUWMAr0ZMo4oNfxE0PFLaJfmqfuLhktv6oG2C1
OCCn7E0gQMx5L/7UIpvLjSB8milxu00WZcZCgjjI6xvmHKfvsnT+xdFyDDt04Du9lBewtYciUNTj
3I/B7cu5TnYxfZ+OevpJS1UAo/9NEuxFEYBxZAxGigv7yWdN7DXseTcM7T/WrGUfrwM2D99gUIHE
6xHT1es1sHn/qMjyrWFPDUWxE+tdUiG1p2cF4lL/NNWyAEjtpaqtnlUmTNfuc7dDW48fNrQGOw3V
l8WL3wNYDOpyAaidbmKSxustYZNy3+XVDk+2WHxT4dGcznJ/Ag8LELYlh01kFV4NjoP21YyB4u+t
e6jwD19QUvaMPsY1rEh+3vlUdiXAV6ZV5IES2b/I07M6PmmdnOvyoSWiBrPPSc+QUGuPhxuvvTnZ
/pEtuspSjd3CZnYuYbJSzcf7aM7ziY+8oVS2OaVQz3xth2SptEEt7P1kpTZnMrYdK1IgUNp49KVV
4xOttXIfN17BF1+Sv6r1iGovRDSqW0fns38PGMDECK/0FqTyEFaKaYiZcTzzEzgo5BmhVVz8kIUh
EXA1Dkp+sHC/Mc9HYRq4gVU6C1KhM+GvzXaqn5jQcrMWaLOO9ROTZp+YpIpgykhMsNwVAGITgBEh
NfwrwMrtDZBWPaF9E+Nx0P/IIHYv29254GVxc/dJ1NWL+GwtgawO1i4Y1cg4KjdDFtM+jo8ShO4Q
A5lIS1Q5ucBIjWqEMQIq5jRMmERrs8khAIyd4HbYdf+XVSjSvMHFS+6Y2siHV/fXwU1hfKeRFmV0
yV3K5/spC3JWEST7T/nw+U8W/QZOw75Pdvmt+jVDKMfjkCUi3io9b5zZwF+vyL4KnfYILUZW8JTA
7oKj88FnCLwR6fTSKecRMHLVZ7uV3dHW2+IBthk2Vt+XJQpPj60F6Nr+Yl41gEUQ+eZ4LPBTcebW
llgE8qPuYKNqb7tcJCOZi8zvsqlnUFaz4viHFlGgAUk7UflJveUJgP9j6s3sOSQhaa2nusHFJd+6
SdVVXxvp7wUfJk5AtexT5AC5FAVlVxs6wM4y1X6QBhsf80EvnENoIplzuMXFnxfoTkBrJ+J5zGD8
Egx1HtO7OO5VKWk1ypgYKx8XnogrC6ymcYWRygXC/xvd6jzc2CMnr8ZgjzpejbngUeHqytDqTEb7
Os9fESe2kutYp1pWl9Qb9fEEM8N4MFhJoFP/wvm0wrxhbO+g5039GAKWvlEx6P6hDzJmJDl+qi+s
UyzuJqZ1P4bMu0YdzLt3Di5BnkojqQuUadXGeWr9SuepL5CvlHFPt9qEgti9M8u3utigoeZy9Mxu
Vk6+nvjDz1O5gTFHFWLk349BUtKsgfZFJE7hXWjpIyF1BSe9sStxk1HEJTMLTR5oxRfxDox8LqvD
yotET283iV9SzlRe2JxnrTnPvOAFg13VLGyCgvo0DCPUUNicCdnZ4SoPsK3U0SpfrCxIuWrgYoH5
Vt35qkCAuKNakpSGmByQ1bPqjPVWsgHv7jkzCHLEXEwzV1PluEaWN5V3K9zhYNPpWu1+wbN68BBB
TWWA72DsUXrbOtfQyLJftf8Inf3Gz3c5Bu4R7i7bosh+YLrVgwo5LkB2LQdnY5N4u53eHx9l5THs
eh8XzP5nGj0WBYPkrDyTXfJVZjnfNbCk/BVlLcnkSFaCELpY2UiIq7AidgRMeyDy0i3UmY2AwJzf
wcvxPHp0eYW9yLvDuoMGZOSDXOPIaKrFRfuPGg5XB2bNRyD6dha478ik/ZQKlg0MRYOswWz6BonS
R3pCRf9LoMcmxyvX6d2sQxbLXstOTy8Yro7hsOGY4j55f5YcE/9W8euGrNL6qjlhgWpTkLC7Iulp
zfVL5UjGLE38YjA7T8x5eZFI2Xfh9fDWYzufxSPLKnymRKtYFzV23dQkXM5B6JU4daDGjul7upk1
pUxX6NlURTiRlkKNU+5QMl50EDZEok9T1IrboOp6W1sFQtBWPNOuIjtds1ZWd8/xbKr6eIy0cXgM
IIIqZiNva7CleY5uPhk1TY9/X0dZq4oOWmgYLSeuCUaJD4Yq/1SMN2GT7sFpSDn2m2Gli8niwg8L
Kgk1EdLJ3/8ArBOCPozs/GtyfynfhF6chTs/u9MHLftO6bapXAeGojMKybidUQtjzgqfbccmx7+u
Y9s4JdWn9hc1Sox+amV/mGQ+SmeZS5pnYke5+mDm2DjTHK3hucCWErb6R06Qr3Ds/kska/vRcsfF
wYhZ/Kabvwk4EFmkeCppshsGGtdfPAowfWowJyyCoOsgm4Gg2KJ3tukVDmU0bYbDJhbAgNjL1ETI
gD5hx84ZJe3QQH3yRPou6bWEEeRq3NrPPwwWFFD6aZ5fRU1YXpdTVuVpa9mlp1RWNzItL81Ze6Vo
Z0SD4kkMDMOB1u5Q5fnuL+tRCWAmMQwU7VsVcu6lnSUidxjrr7keOaI/bsWcr5G7QwydMs3yIjM6
KY4w6vuDyX75bp4x5NJQcqyFJ4ANRA17itgqFQ90HKH9Br9J3gttxqA0FEuSFGX+IeMFufKLbjU8
+N7BC7mmXJHeqJ+m7Z/pqTOpOaM5JR2Q686bWGcBDIimb7jTDco+9P/5PQ22i+g/HZYT3lswBpaA
ok9NCU6CwRp2/V1sr1/tQacpf2BjfNi6fUNL+dlQq2a6uI7GurdkrBzExKk3JPgPuSbT+FKAiVcS
d0nGCBpcv61QkiCzWeX64IXxFUfY/qY11j6RPL8/u4FTdEAcLLuxNuUQvPnFNvuxC9ShzWolk+t9
s5Te19iOVgrHkfzxZmn+kNirus/fQOjwAWDMua5IiIEuSxEWeeTwjpfbWoMRZkoXFhMrVSeA25/S
xYAQB4sAMcyCSOUcdLBexQ/u+rjvD+NVzCaPOC9Rrdm4CZSlXLLbjUZfl4nfLgQsrbKfJi5RcZRs
KnLwJSf68H6Uz4SC8knbBISvxGb0igS162ykHNv0YpCwKhOo2scvGntiw9Br405VqVbCub22g1K7
21hmDcFY9b/Xg6gFCktsa8lEY/jnsGj6YSi2NTdtNKXfSSYvzr6phgkW+AasX+URG7n7iJw+s8pF
JZ1r0Pp25jQ0aH2B7I/osVfFlzzGnvHmXtlzHf0r4ucqAY4Tq2FFnfO2w9G+V+4+lK+mFZmTi6Ty
sbR8EGuiXbNBh5x1mJ23ZbtuozrcIDGcKpM+24r2Pe7Ih8T+wNtP1pdpkOREY7Xov9+9goPVRT3O
h3EE0s6WOJRS3EJd2Xg6ulVy3q3phOll/Je0aSYuY5iSM7iUJ/Dq+E/dADxpaLmsQv/mo5fad16W
kvnmuqG1f4MvKvglTr8LUz0OE0tEZalxj1ufRdhVfvgN+zkGaPblGcaK1pX+kRSl0J0/Bp8ENaN4
jNupSct1fAaV3pZUkD/LiOYRf2QMDoTApjbRDGydFbbnTXZzECHYLGnPpNYKllbToKz14Fy24WF3
AmoA7KE1k5GdTnogYPjIvqUhbCyh1NdDZWPSZIM7NXw7ToogyDsCbcWl3EujOOe831Ts+qtAizjg
SuXu9y8E+m7BqnnnqDQdKV9lb9ud1xNW9Ae6shoWXY/WlIH3EAmfh3JtmGEXydWdclle0UKE22Tl
2M9fCCP/poKxTBQV+Tf2r6Zmx6xww6KEgsGiI42Zb0sA4PNSBQ796Mnz2OL9PTfBb8OaP3eyLsYs
9o8IXw9KHe04kWu8Wk3E0CUE2Mi5N/jncyYRPtZKRHLuf0tE86TgeCeDSBDBZGKAvY8nJeIVxOmy
CYEnG1tc0DO2mU8BuZ0JIQ0YyZoFYxeWO3B3OG9sZMt0Y0Ss2k6aWPjP/UtuKquBR8rYB+3FvUx0
cLHyGEvoJTZ8wpWScZ/IJ17XArQrW1UYN3yzj5iGyXqmLnIgZirfqIJ2DggEjsWE3Fc9zc9ogXIG
ZJ2UpVjbqkQxdKz5uslx6hB1vwIbQp9ZwpbmEEmwMQ4lAsj5G9bYl1h5ROjoe2FIYB6nHmloXAm/
FDhIvDv/z7l9cmQjdaPdY+13VpsiJt+BY9lDj6Fqq7CYr6ojKpMxDVAmsKQ+MzMaiuwxeHLBQJ1z
M4XMT0kWu0J3NfqwE++NKMKqIBbo3KWjVnCKkNWB42HVjYgykPYNtikl8U408l0M0skKBP3eTPIs
PygI8srYqERHhAVLZUkQx1CvbV/wFUijg08UMpJi3W3DeG6xHqmh6on8IonV7e4iCuBdY7A0ytpV
KLIORlFvLrI3vGZyDsjMyKAOrCf+DPk52qZFg6h3pbujZDOiVFEwHQYzDdBK3iXjGjVtdH1ragjr
VsU9x2n4keNa7fSMuHq+QuJBkbRIDoGW2vxLlBh2c/nUxU7nY7CoaIpybZhduwG8OFmoUK9CK7q3
HIyFkDUR/piEJl1lhsgKD2cjHmQ+sGWxxZxWgk8fDiz1qT9mUlKViDDxW7yOkWzsR1+ztOpV6ZM3
nq3HYRZlB6JtGboBXUcjnhwbOjvnlND/KltNUIBPOaRSKd42xyiItU4MzoNrNEUcwNXHPU2wSvO4
DYyxWac/xojc2TFf0bc6+nVOl/QSfvKGzZ+kR9zJ7lkcmH/8YcC/q1ooaniUpdo1LLLijr+I5j4Q
9kvAeN4l1vfUQlmvLv3wYG6PcwULRRJFjQbnEMfNX9t/MAUybchSP6mFrZSZmaTPYjtxHJsg2zan
JtCVkdOG0g8my5lTTHf+Smm+llYVbDS0CTJIpmj7I9d3uqCSqB35M+tfH0UfL6gtzZ80ZTsTPE98
ojDch6T4kbtOpOqTowjDmEwNdLIlqKfAptYogkX6BUctLGYgKMDhT2v0opD2mxjqWSXqm1RCabWH
J9VjKHHCLJdBulAolU4ydxoniX+cT2mbZlBQMIqqke+NC84lQfqzLIV7kC5DUQdSA3Xy5J8YPIDB
qnLyY/TGGRmsmQT7dPoN12nJKq1DET0ajXHZCOEM5PEdsxzfS18NkQf2lpFiXyMUEf3jaoctlgzd
F/t4e/Pc7VGDyDJrGDkgoGPN3XBo7KuqWcJR8WIFg2ONniVeBvg6lYSAGADbgopQ1/DD4fuiBs7z
hCe4ZDTKt1jbg0AHbTiVDmNbpQGPZuXH14BZDqODzd1Jib2QZibJAvXSupwJIbK1fKfLWWv4cogP
44hPxby/1XXyPprrijYRp4V9GMI4fLZFsJQiFvU9nkwEQZoDZdQPxam1g/XmU9rICktz+do/1i6j
TG6OD3MR5ASP+KOKsR63wq+4DqnMJ5kPnsJkeImsZe4R/XHS1VDFLbQCWe04HLjwaMSLMphL0WCK
oLFGYmpeIcLe/P8z4L80ZCducViiPIwWoiVxoZZKv9D2ND1bDEcdE9Ezw7WsA8BH0Ao3zu/bEjJ4
udYusjw/W2vc14wmHa+N+IIeHuD3gCPYvk66F22xFmFIDg82TmNwNKSznVifeIC23v9Nk4VH8wkF
FZi9tZjR4oRxiL4s3wF4XCk5xduaAXjAcJ3jOFyVsdafzptGYATyeDLezY/hj9fAoT8V5aSkeEGR
NOz+IsOnB2PD5/vbaAzWF5KznOQ14dU11LGIiYXteXaJklKFPKjNfdlWfnGNrj9Pzh2Dw4vODc7G
jRNPgZcZxtgp/XRudgDoKN54cK9bQiwNx4ltH2HRTir8PTHOe+knCm5ofRb9tFTWq9CLbIpsxoeN
4c/LAcuOycZl+LEiIjLe3IpSmPOY50AKox5J0AaF5nFmibV/4fQliZnlG3/gGmJaVNQAmzUcLVQJ
jq/Kab5abY0Y6Yr8nXaERhuYeVIUxpkmnlIf8MpwUkV95euSFrL2DJ5MK3AkZlNl+mMnzhw9KoW9
4ZZkxpWYtCO1BkIA4c4w04KmczVlM5d4uweFy5UBA22F9NyYqJM0GK5PeW3nWiEVy2rKkDmwueXW
QWC6AyGYDDdckXEPWwr0anYu++9MDwr6MzS7ycEJJ/zQ/qBr+rw1A3Gdf6jWo8eCznViwla3sOHC
09VxQYRRwt6OAdzbvTyShtj8wDuF5YACD2110/Pe9OPIOeL0r35yIc9wuf0LbNTp1cw0wwqrCvVK
7wF8NO0vVinGKldG+dHMZktglCE83guTJN2d/O1H/YT79b2HLKaJFTNt2SGOcTC0UZkLU5wHU7Vv
1gb3L8nw3YoDMRwDZggJkwJ6ieB4nZ/Y/rCFMz+LHTpLpWe7W17HKeOXsIGrxRHXM1Lh4xNY7AVf
gLg2YuSkyjDTjeeCFSAWq+zwJ8cRZGdEP3KYLilGk6bc70L/oTVUa/WppdqwgLPd6hOzzvjjb0se
z1mX+mxwlRp0ZNH+2S1TZj+bRAIvB4OJF+7wAm8Cp8l2UvVIUE19hu0BKKhOG4rTdyrtMI8AWOhC
xKfHF8BK8aS4IXhzuPLDMaaM0lfWGeItnDSbC4xs28OihY1KigYc6gCRa1Klaj6GGx+WVo44YEoC
ezQWXwiCa5dpe0pWOc0umlodIWAEqg0aBssm+AKckm7DQjCiciDrq+sR6U9mIvTGRye1xa4KWEN6
YnMmvxgwswbrR5DlRH3BwOBCBmj50EQX3dV3qFHdWlVgrHSAI0UMU3r/hlbSp5Lht+nP8sRmhPYW
fjVNOwkl5mpe6swTXtYaDlyupRh177kROxoHwBIRpOFIgPFnJy6J5Mxi9ZfNIEWPozmgqmcyI7m7
uv3n3LXatWyjAUoYXfMkBdzs78IYtiin1tQ4M2pUUwTOe0zPtf2a2eqsyoZvBOoXCOvzZtrbwymZ
oyCD8+l25DgUtNCMVpnx3SgZ228v9eV5hPyQD5s8Y3XDlS5NsV/fxNRdxXcDHNv+JRv+IlPgVt8O
gGkgV3HMvYs04SuaaKEyAjmeeZ8b/E+6cJZmp3bICE/8heuuPy3CmgF3EarhxSbar/i2U/+YOC3m
6bLRwkZFTr/agrruydcPblrpkNdLCi0QsZbILRvTF7oNKZU7YDedSdz8Zvr5/z+YeTlhv6+1Pr1t
ZD/EU2RZtJuBNZ7PAm7WufK/HlhqyhcprdxYXEHG6V+7xo/djJGPxjhxY3BfXENM8nlhmbaRaaQy
mToW8+n0xbG5zgcaSpHYCzPs0O0e+G9XLgHx0S1wubKVSYH6APky2ws9niRKuECD/YawF26OUu93
ZvtMbgpZRlUTXmpgv4Uzk0OsbMCi2+A2zMr9ig324c/9ullBxV2zN7Skxavs5/pMmm9w225UHsDz
wefDEilJiukBYSsB36hC7S/JlIqEihEkqEhWCOX2kfncAZfs4iw+atPKVRmzI8VEs/XnkH6Gme38
7xICFZI5Fa1flsiPtQiztji66OAdzX8O3X5raGvZZzPJhauS3ItIa4jXsCroteiUWdJxVTIKRizh
zpNjidTpxIaHoMd1M4k1bmp6toCSbG2BniBGKO8ig+jj0hQtMdrN+McvjlAG9oloZE7zZm7d6xcv
EcrvhOv8Co7Lv1uOGHcU++56xFb5jNdbzg0vgXxb00LJOBxg51+S3GksgScjHUzlzhkOfdjHe4WA
iUV1BlBOE9C9FCti6+rdpf/4ODYAOkRl7hEhf8/6H/+sO5ys0HURa1WFnFggYPJYSpOJ7HkdpZQY
bkyk+1vWGcD3NxM8yB16ghe8z8lW9FT7lb2ENPGfvvmGZ43MNymqZijuEBNMU3IXF3HpbH5w4hba
sjJRH2ikLCpMiD4Z6Ad8M1s3XbPkm6MUXE0+o1JYFyGjX+iX13oTo80EYqH44TWMCi3bHbMxUtdp
MDrksLlKZgFnvOI841/JqQ6ajdVQXvkL6V8o7vxpeBR4mJVXoiyy/6PIdWgAlkgpfnL9+f66Umbv
ES60gI7rJS6CYB+F7silprczu9qJXeBMbDMb1cjQ5jbdQaDROAldZeVXKj14DYCLd1B8XbbCU9UL
f6ndYORofakn/UuZoM363mD9wBKg/kRZOu9ZO7Y0Ohl3VqdTM+UKdmOFGnEvBJ3W2WEWxO7P6Tyv
mwos3AfSUz1isTBMPYxcrhyd8yk6KqqBgaFXFtwuBP7QQIeAV4Efgds5XQEpOqaFX3XB/ZbYRWy8
UC/k1/5UcquA4kRrqsiQtpgLeh2RjGvyTjHLxW3n4R9KC6Uyg1uVVQjd0jQt6CDQPKJnBlgmSr1H
g9DEQzA21guWzgGKsxh6Y1R4kb7ITZGIaQWt8PuiPZhuqudQD7GUj46XKxHLv7hKpkIL1Q/P6OLG
uwKH4V5MvzEgmwBeJR9uiA4nxYJuPfS5zlFOJe9WpBaKIHDtVOWMCFVRb7JINcWmBAGg2lZT5CeY
Rn/k037HEWtiwiWXKN7ahELIF/xklBjA+Xd6qdUIfqAZUfKhbmMvQFjJngvbwRZpUhvVYksLk2DQ
N4JyZRhacrb6ggNMIVsExMj1ykdZX12wVmVm6MeUCn1XHdeVMaQSaVr/okjmQ7zZWmT5EYEknwX8
4dxXUvw06hPLKrBwi+y9fhg9zv1jQMgw2z34K7SUi7zU/7xQPAFkXg/iRB2Yci5r2nlqISVaQeJY
NkQEnFwB78U4BY/h2g29oGorqoo89DjNuuBVoOrcIl2ea9Krlp96I1xwp6sTdegkjJjNS19geh0L
uJn3tnubSfqFht8klFumwfZRhNiX09s6whF5wv5MrB+8COaZ73GKD8Mz9m242sAdxAmCAijX7NuS
oFNqhqoK2C82j45Rc7EjF1T98tgGS7EuIRYmqSYKDQ7i7VM0rWcuUyo3t3JeY4SQK1NU9JHMZNKd
mhJzd5/wEe/rNPQL+mZsq06nswwTMboPrRwCgfNm2+1BRLy2qDg11/hBLI1iGWiJi0WMNeP8FutN
RcDISlysW4fuFve0EMXFt+h8pNtNZBWMs6KVNebwZuehSpHvF7iognzMRfhy5jg1Pohq6G+XF8Ja
73mWgyvXq1WUg887PWSxn1vVUGg7ANt50DAEbYaWuLURghP+VFjKJD6dS5CI5e1eTmrwbySfOSjh
jYm3sSWNJSXcAnLD/abp0a9B6Np1awWGSeAPqNAyF/ciQEc1MlBvVu2Y9KZQ7unIqqYmA3Cfzrj/
0jgxzDv8/JJKAOUar2CVBRQHPhPkpPw6BoM19fl/6G/LPsUJWeiofkHXfRUbFNhYTd62l7YtNsZg
ilVbNfJ0vKD13bOk/LtthH5kJhnAS9djLp69XTjzuoF2quGOBZSzF/Dojyi9P+A3WIGcObW45Hy/
OwJ2bPaJYr/MDU61OtU3XURstxAIJdzms4NCI4h7vZ0OXynyd6wp/fdO5G5twI1HfAId+K2PPuDG
xYN9HFC/zSH1P9N+2X3fLhLzVdU2AVRUVuDzKOiiA2Itgk85dT6wXqGM6+23WhCM+/Hx/m7BjvM6
JM5/wsHcQqTwRmBNRZX5tvdQLb0Jt14ByaL5onImOAuqC50ZAnJE4WjC8Cay5XPbm06XhxpRykZA
ltpQ99seJ08x48KCSU2+fxvAKYbY75A4xZ1K1Ov/hN1GRlpBjoOqSpoRKQV2tb8chkPizDrKnZiN
j8o5H17nmZ0uknUhVkFet3VzapNfbAig6amaFAweb3JhbonHRVQxP0gW0s2FReZ54qAn0TbigqEp
LGuXaP2FQtREgJ72wQS54LQqOnSvPTAaTc72KdwAPcTuwTLiXPQ3EN8WK1UkcgbMUpdPVzzWIXcB
8zGZYvjIsi6BIdTplyrfzrRDt9KpBaPjE5zinvJMqOYZlbIXdOMeLDe8B7J1uPgoYPknEJaBSM2z
htlR6u2sepNNGWu5/BqR1rrs10I5ohZIEvorvtl8mhKHRg02TKQ1iUEUW4+q+2oOt05yt4qX3G/t
LMP165G5IVOOP/m5bTifbjJR/gIvKeAq3Ud3oqABossReuOBt9u7gCHyIBD24VRJK3jnjSE9pl2/
+r8YfobwJfivIbw2kFBhNZIKW1JngASrfnzP/Z1JQVYDkOVE6LbXnZyLOrDM9BaKUtNA4lNH/hik
cx50TJvTYzEHOPYugCIviZuGEz+jAnu5K8mifoqjD3zo+lBonLnOqZIcM8eSa98RMB2wbENHLb5N
a8JLPogYH/NXrfw4Ad0lGXY7S6s5ccnoPyjfNJJq/cA9hPTf2bfrh/der6W5TGCZF4SZZX/G1OQp
uzfgjtBaeDuP5jiRV+UvrQBYPvXy2yQH0NS27SQDV5/M9IocHBC2lUJfB1xMebL1fsu0Cej0Ou08
bVzwg1Oy21+3RwoUv/m/Pa+J25mJuNv6IEXosWjXUdae01e6YY3FX0Am2x9AmVPmSFPbpYsR7KV/
3N+EijjNlIyruX60P1fn7JyZEw9DoMVnv4ZqxzicMnuZWAvA5H8JSilVm2ein38tFimn4P8kz66e
+B2KEpjCdWS466tXz4uwF1PX6xWT7SxHHc3ouy+b3bJNxcqGYTLtn1tJKzEokbSPDsPe222xKx4d
ZDfRDDjQdjEyO58VNw3fbpq0TXLS8JrJjqphZIcHkhtvE0avO+31Z8IFlLvf1d/oc40oJlJ/CUR8
GkJTzA9X/Tlmq1vSvPRZUX2ds4FL4nXyUEjNhwEMexEQUFfCMJNyLRG4oQwEgOjZHNl2tHnYc8I1
sksOg2GMpXA7NS1cg9lp3CXcG3m2oYRMuvpN2Qq9D6wamJsOOEB54Wwpu1xEkMX1Sb/eBzWR8I8v
OtzjuB1BFxsR5DdhsSJMux8gBeJhvrtl1RNZ3hJF6/g3apGrVe8VLLbTJrK9d6PxOldSwH10G6NE
9YxgFz09BkerxoilMKYYa8tlCAExD1Zq9T2fHlJqHp1tLa7oMwFlwl8Q5RFIKWMJQb1FmlvNwaNI
sFTmUTnkHgwZ15ce0sjKKf3zFJWKQ6EGN7TdlrAu/kLyewNDOOXaM98HWAbtDyTod/oj6O6afzHr
ac6nGUij8Hne2zGO4KTyDICPWBQDr+x+PBCHY7ND5DhoftjcNphMCnzQhqNTWTp9USGpJIs/M+BD
WJdRtaujQ0N2Vy0cR5nmxjUv8Hv7Foqzd8IdI2kZlSE1ND/j+RyuzarD9trc63wxFYSek4XgGP9x
oX+/ZmzqTtsxkpVe0xRMxh5k/RE9zP5oWAK1rH8yr7nG3FbyB2x84+n9R5g302lKjIka0mgCnraP
/TQZA02Nze2tyVDKnh6UQHh5CXFfSSy7wFABamEoIPGwJ8TwUsP0s9vWYxaLNrNMZzA2hPwu4TEm
+9Np4Qik5LhL/k7xJS1duukqf3RprpRnKRxjMq2arI1bE+zJyvOipliUF1WEZSRDbg/jGgwLBPaw
41dsLbawpxDZ/C8D/2vE1sLFv1DfdNLJgxTAR4hym3mrpGAWDPpL5wNFwkHGmqwBr1RcDCZ/GoAJ
V4zNdJCNcpJbKL6tiXvc6a2Y6Jj+kBdKArh8gcmcSuEcQexSBFAoH5a75R3V29PbDYlz+EIVQYN7
BIhSqNX3ZklGxZ1UUShYQ5BjT4knK0RIK3NoJk4H7R4b2ITkgVsAOJLtEkqXYf7kXNbJkE9/Ec8C
jYjB/H0U9/4LRlevf6/+qWJDl7nR0tyFduAS4Povcbue2l94N0N0dA40v/JBfda5H/5uIYdILS6x
o65Btl2UE3Z2bnbhd0Gy7CXGHYCVwoSAkl25j3zU6cTFiBhAFP/OEZWEQlAOKHhkL9xs9KDPmhGH
71sd45Cgr0OTRYPcnv2+4LP6AjsONsVIIRUpLHW07nPs9s1wpdhSryDt3126fEd7rmPczzmxMv3R
dvc3a7UucvzFoxsTt3XcHEzlvDvOiu2mu9sWeqp8wKh1JhivJBQR2yo4A9yVYtdQXS50Rg7509gJ
Ky3pkDPvxbHLZBPjoa3pUMaYp5s7rmkjpz+GJk4jNBdTkMpjl1mxEjw4L65QzJ6hbVdjwntscoPR
95PI21hXtsJhUuPb9q8NPk+Yl/cxj9wrG9cMenXpBpzJQVoFTxEa/e0rH9cDf+0cxyqBIsBPEsMy
KjdxMvZGC3nsESSiTviWrYlKSlTJwEJowY0PLzdbLwczDorQRTVUAfzPW/ii2SYUozQ2nBg1bhSX
GEjT9IrXHBsODGpcSqYeUrLsMPeMG26ihHPjIVmklDpRshhcdIBUrxNxceUf2NHzTQ4ofNChQMm0
31tlVrmqGSs5Vqk5pCDbqANV71VJKFrtjWbNXHhIy8hBjVtDqcuh9O70rD2ureRDoQCTqGXkIH0H
vXX6vOpK2tQ41TtWNVBy6plgLNN1R1eE3DpnHOYTqIDgTHJTbEpRQ5LW10kPFAhqEYUnCT/TV8LP
AfXrNTGebsbGBcpjKbBgzWsTtRO9Srrdolbp/mWcKuSE0vg0JlRbmkA06NjmaZcRIqsD/PRdvlcZ
jDaQTXE0fhg2pO8MCBiC1kw8KMf38GlkfDxGk3qQaM/76F5fWYZOAQpL62lLSKiERrBqcFcwxXyN
kXGAuvjj8/i8Fk7zDgWvVlXod2jEeYPVzfD+IUnAmZ9pVLMlzKD69qoYDIb9UT5S/fTIJ1hUW6MU
YdpZAJmQQ9r4vXOvVHdHb8SO/kaMeKXYrgIl6LYWM6zbGVuivASMLc+jfJMjaK9XR+GsbPJJX8qX
uyjxE52FOWJl2rNeGSK1p3jAexuA4LkA8wWyUP9fxSbCTz+DM8q5F1jhy0Slol8WvHor/xkv7kvD
8HJZ/mt6hdy+1qBZMG7qrVqcvawRWywKXNUr0JYnlRZMjEQEaPi4l8eoMLh1q7X1x/D2ZWjTMVV6
oJQLSzDKDKDdcaan7230i/+wLHQ+DOuhjONoAbeLmIL98+1bGJw/n/69Qs0FJ18FIaEBxJer/JD5
cCCs9ESHmbZZZRcXzU8d18/7wbOyxEW+Ma5v0vy4ZvI4syhrpHuiUYOizB3Y3h2lj4Abe5gbXXkv
U3CDseSlWOn1oAdCS0Y70pZ2t7VqMjBFHdlwcP969JLoAs9gxocuhIda8v6uhpgGXVPLwDY4qXgN
D376xvrdiPDPRJ9uHy9XCK8DAqUb4qqmNlNJYL+lFfL90Au9hx1k1zOgaPrvfbg0I5ezAuc5fcCt
hlwSg750wt5Nr58M43alobq4WT8XbWiqPJe3EjEgXq9s7jtfvPfuUoB9uvrtmnqvxqgwzxacu+O+
6345McTzAxXq28B99zRGdLIjaYtyxs2Ee83zuim+HOLPqQD+W8u89CQmNYaV4bvja0HdmIxJDThb
QC5HK/deyrwEF1Rm4hpzHnfh9Y72uTW3rSNRN5diqCJZ5GA5SllzUBlNFhlw+NOejiXENaVUSThs
wTQj6zCHCkwupfwGipsKsk4aIKh9uOSMArLJOCcOo0BAi/7pJ0rRJ6PPuue7W7Z9lFNtvBVcuF9N
KpZ8QCTynYzCL9kc7e3J4tMpDdEEXRfyJ9wOVAOdkIYlBG8746Rl8x1auKW84dhmyU+oAKU3ix2s
LxAkV9zRxCTYqnvJCjczZ5JPwdETDwHvAAgZAHVk9Cx5NBoIQV7Nytz0g+w8u6HXDW8YuEU6Qy3v
0LBHLZRJGjiSCEPoOCAQycEeTFzFODgpEvmO3zO18Yca8hqaqygI1dfljsgGeyEMP6ILRZWNuh/Q
GEag7oNWKWoBn74yPLwxGUZ3oySaeqOL+03k7uFdXHjTbGkKlJXTAK/ZixLe9+pS9B9sVBc91AyP
auYhPvASpD8WDvHX/LbptQVbdeB/EghUCWgKQYC/AIF4yh7U4XeA+YWI5edm56osCmFmq3iWuvj9
WFnjy3VD47xP4H4GgF/mv/6Zhp+W0R2FC9op4lg6yD4TTmn2CCzXAJD5dAj1yLGqljfNgX44Doyv
2WnYui4NNQ4lLY55PwSzFMRb3XxCyrRRTevykSKiJoFV0MonMOW6NEpLJHaxhPD+ylQ9S8foiTVw
8oLDlQvPsvPo5Tu7GVtGRB3nod9ELa+8WWndaBnfNjmd2mOsf7+hwcXKPSYwXBFa56xaPlD81tQL
UF6tcmI6Eo749G9BhCd1lKuspWcBlMDhBVw97JAurcxUB68cZ1d2oo7UeJAS1HQJXhM+T1H4Luc3
3tBCW6WRjAPpAT8GrLPNppfA1ki8ytWHNdYCHmODazrrjzYypz4fHp7fEOYR875rFyO9Et1sWvVS
sCnCySudKnYUuAWNbyViaCLdPZ8AoSe5ISWpcMKv3DV1QCXAmZTB/ErNJsjcjVSn2FRmRgDywANe
pC4mnC3+sCKSTeXc1Bo0zCexXNJHQxq0KOtHkoBzgVOYlzevf0uQCUKpk81yqrxDnLV7rnHkLYvs
XbbXfuzYSRhMKuZtVD2ya/uszecNToNKXGN3RI9Yqj2zPpOP5mpkCNz54Tzd5dI4pcY97oxBoZCt
r0KNuW44eftoIoSlcftDn0vU+mrSBGsJqYTSR5FqJN2zeLhI/eNoU9WYs2uEly8n3/007ka9F1dr
yr2tTw85mGdZRXoi/Zo8mEc7c+8F3wjYN/3q8/0CFQXLsMFIihi4Ufx2XYKHNMxscCKMJtXr3FpS
Wmh2fwblilGGhlOVtTzXOSmNLtJCgczsjAPkX75VITyMWvOXV0Fvuaj0lxn0lIW1SLHQf2tCM/KF
QRV+9fMVh0CqJmK+S0X2FdT3oI25/o6CGHM/cgt1KcKj9NsXlPcE6nmGmtMqvuUvmbmprb6zmOrx
U2UTMEI3pdxHBXLoltJeWkdIjUKNiR9zyo3MT+WkY7mjHjf0Hl5t6cBPSyQAlR7dthbcHZk8GFjr
0vQP2KFPjQpbRzHDCgeJSWde+teRPKgRfc4x3qjubNkcn0sk894zi3V0JZsRf5Zn9cCOZpL67rIe
HkoiE7E1T9PseByB+VDpzS5EpU+ONtHtY9Wf4xYo4RG21yeSnUVzKStVj+W+0t9eTxWBg1WhYrGJ
22HLdXBJ0bk7+z55Z/g0zYDYdKrp91lhH++uY6m7Wlop+pF52+oSRic38HoUaIv6knS0L5d/8Nev
Pe3f6sVny+ZieQH7R88etUlFi/uyt8BM6F8f+YXUmqUaEk3EhMO1WcMqLL1tnv6rthEDcWLTnT+e
n1YDFYMqVwHQp3LLFBdYhZ2GSgxovVwvisGU5X5/h7Ua/uhCqrundg/IH7SqL0DzxoTD8Np4jH/S
+AAum991LqQtephb7cfLngg1XBvoXUtBruiz3zlPrAZxpuw1OdkAa5Xem4/cYsVCtyIoq0q649Xq
u/va8GaTXzdXyGHUvFI7jl4c+DDZXtjX9+Spw+5zbvawASKeMFMwHlCUenrHNxS7HlqGBcZN0YrP
kw2RJQpsFyIMm8FyxUhuY2rHxzTy8A4koNAv/a1Dc2cyTI/Fa89KCe16Rpe7D7I9mQmualgsjD/i
p9rmDfSpE/hKd8OK2kQ9gbMmbvlLXiA3lEaBEmkaJ7elLl+G+KnHycn2CSLa1NP/oiPkojgOmN4e
m0dKEIoVL95kfEoPxm6QB+6m/xOQzFXfZo3NbbH/lkA34alRvTbhCcAlK6EwpxmEcWB6OD3Hl6lx
H5wvHxS+KOZt0cpLizyUt4x8cc1EUFOIKsyI6HBDwwf5MNFiqyycImh4p3B0UFXiZuq9zuPjcI3G
UkDFaNfJPbP/SMmi2Lgn1oaFGQ/gH1negmy2cGCPcaWcO3qcS/Fy7B/wEWrJhdDB5pihSj4vIBLd
4Cevt7h8KvGL3dc++zo0b3KoDCD10fa0Lqe5jO9fIhTdISgYt5lzQDV7XNq8zCduAlx+C02cLMlr
evvhuYq6qx+aZUbD8Y0b14q8HJ5Btlyjbd19xIqxySsb2CqGBa03VhewAky6LBEHUxJU0cg9fQ7b
985K2zny95MzknRu/R6qTE1ry3KTdyV2Uo7GULPCv3WsxTTCwL3nv8XwkpM1HbRXFGs2Wt0rnRPU
TP8KybbC8wBFiw/amFBoBIdC7xe1pevMxBzb2nRx8UHD4Kyo4ebf7PHSFo3p54ArhDcMohVX+yHq
dsEBViLo6vubzQ4neaFF7vhMQg8Q4pyNveUOAHdEX7BE9BSOTVapy+ynVbwQUQ/Lhr4bRDnhIctt
QXmH5pbU7AGQ9prcfJvT45u3c7w+twtzG2bqqf+tXTgCqXKYzlk/e8+dQzvbn+F+4imQKXeyTR0J
gPWaRL3tNBi7Pf1fowSsUEeppbnYEHw4ga5eVkVWJAguDjrMI0X3PObgSvrTcrMG85FYDonQyaHX
9WoS5DYMYLMPNrFpT52qtq+fQoOi/yZirrTC8mLzz/4HuzAij9XL10qSPXhB05PQNJE41aUkT4Tw
8sSFICo2PMsAE85ICUHXYwtiqa5/Bwl93/zXCAAJfYsPACLLReTHkMAWN01A0NbkzpDDYLNftQ5M
nNMXfD/+/wwh29TzhwpuMAjbu11ZsJJeBKcWNIEXYiQJC3dVhwxZ4gCm6+4+hjAGEwNI1AMvivKe
0/EbyZj2UmTOZwSYbOkhsHxlvZEisvF8ueoykrU80r1mCLzZEvj8XVX+J1sLYlHXqLlmNSbkN6Ey
s5y4abwqaRjZPZudVXKPDFFRkSCZtOKE6OmGloSZXbJjm6glnQrspjvnUGbqOhuEst3UDTduXjHc
BnaBaVGYgSNEBEDPRdOB4irYlzLuM1MJ5+bAoiVsbXN0diDktkl8Z7Qub89CJ07L1WARScd/xvd3
odoXuR7xtA5gDbTkU68FqD3yr1NWYHsUT6VVM+pegoceft0PKxDXYcbIsltuay6z0qpiONmX16GB
VdhbopSqte8BjUz0XC8oiFX/LQsgucqNaIgUSLHaJAI4qmd0qZTRclLGU7A3sY2HSn01zIlXmAlT
lbCv7gPDP2sT2W9lHSG6TE2uhQb6LLr/ij51q60uaNUqj1/vRObHVTpO5DmuEO8LS9JTh2Umt+um
XrqS5pB0HRl+RPBxeIrbo0SXxMErH3s8ng0K4ytMcOvFP+2/R4Zif5TxnoDGLiDUCo/4wJuzQpKj
m106IAuRDSveUCvQlqkYJOs/tkyLnREKPqxkIgRs5gutuxHFZb9Ekgq3wqpOLcy0fVFPzz63c1rD
bvqImk4rtYVNw8cA6Qp+eg/ouvNQJsHz670ryhU8nLyiHU7GpJ+LcXzWsBfEs/W1UZ1+1/juIkBU
T0GDVSQuqKnYcPvFXnfLK0FDtgKEztwKbmOJhWQcm0ooWIJZhxSTX8kdHXMRiH59uIPqdNv+mhFx
4+JU24unz3nxP445vnu7jKBRFnW2LGSFocKhFt/3xtN8QJo4jM8BhXzW8+XmQSGVqluKfQ5V4sXO
gFqq5Ywaj2Q/G9jzTLhADuxVAeDy7sm5pcwkvNgG7j1qXkmi9YoQgt2mpZ3zOfYBPoXdvZhPGi9A
mzlL2TCyz556hgSWd9IBWe/Rhg3AtqAsVthk80ZRzTbZBchpYwEBRsn7jF3BZ3UnHSuitXndGkxJ
8d9t9BcRnAxCX3TMLyS7185BKaRYLx4fWqMhTBrQyAUeMmL+/ZT5K3fRefsH0LPREdfHLv8rnFsb
nXZWyG+a8RDioLTqRuY9bAlE55qi+3IMuKbAJiaDK0lGm/cWfiAkfnaW3ofbdJettMiOVm/klgPL
VGOcildpINWE8ChRmj7oZg7IsQllh3SfjK1K5FGjyBIsFXxGeJIg2eUl8rHevHwU0NSHUKPjCCRx
nmrG3dy+WikYjMS9fGPAmnyGYpPkJY8dtzXqwn9hXMptz1EY9vIh7wNjQvwxe6d/MS+CHXJzTQVd
B/XvpGdyvZ7L1iblckLXutLwJQjV7rVO+lu94hAs7iEkef/N0lswQuY0IX6xFsPcqe/NX9jM27uB
JkhaxmpUei0nlkQ3oy37HAM5NnbuXZmTm4m/Gx3TPSAto3EdqDob0Nermh1crZEefjiZK2Exr38Q
CAYgV9oIt6/F9z1Zc0Um/NoGma4TqhvXRwmv34SyM8tn4w7ZkA5dpVUYJ+bsoVLsCEhmHHkiPGJ2
3lItB+n65qIA4NKz+20kgcJlVySe1Ou/4TBrwZbqJa4BGxcPJOSsnVhHTVfn8u+5FSbf2mG4Nroh
aoIFEzHkCLhNAksZixwFx3EpQisczKxAgBLWmhyg2nZSysPKzZl/IuAlToF4NYhVpuEbJyiRWMbm
l3tp4DoOR4DeF//jhhyOH7+hwT34yAMWK3WMzZemgVfq0/hI29u8XLzx7ymV2Mgt22E6xXR7CBfY
+IqybwyJDEs61ZmSD3MGTO35IQJ4Gg0jRt+TafzvNOwr3GnDqCtvYucFbREmLIxhRqxs6HENxtbD
NpnweRDvP8Yk8xQ5stJBmUFi6kquClO/VewkwxPmNofC1OOEE4RCmnH5PAlQWqt+gux/XhSEjUgL
/x3REuZ4BUgRe2SLcq3DlDzadzG7XZzuB7VOiKpwue+RlPdP5FHlFyyXYKbE1c3ucXJ0bywxT7ZF
SaLLjEU67g4lmLx5KKegj0KaSJo270LV5bIe/PmUJY9/3l6RnWfGwj9M1vuHj3Q2sA1e5mNv0awh
U1ThkJK5BaUVhM4uQqeanCL8RfVsKlCMYAhDk2/lBRBmSuyq6NST6/RhYjUS/ajJEs7575ckZbui
/sCMmgz4ellTF/gFf0nyLWWkKb1PCRyGr2QEX0MbCg7GLBP35AD/x9KBA3mVEFBTEk79mvfeF0l+
qZHZmuA3ozVni8LSWFc02SkCJwlMza/Qb1+9hmBUooApKFs38D+pe+SnQ3rgWijSWogmL7rR7ofh
Di4xctCZ4I/x/UP1LLeVi7BNuLJXJfN9G/dVAVk1DOJx+msYVca2KT4E9ifFOcvgaUCe1y0W++Xx
J9LQv1AFApzy4dCZk+02O657oan1FF7utQWPVbF8QXRyyDRE7JEQWiNNn6tq8koHjZ73aQN+dS3P
+vIzgijyOeWkuJRKBSmgsV3ZynyVXxqfzLfobeW81axRVXwdxOzp/KXl8iTf/3apzNT4tMFmi+sA
hdV5F2BIS+zp/fh+g4o64EaouxkVMZad+DOwZbxGxudLAyUShM5cIXCOACo/nfMTVbwCsQxVNObD
lAAv4k3WJgfih9hQr8thas5tZH5aEvFPsxWqytoQXx2SoZaJaT2awDT5CinCUzGat9t2yklNogeX
rbDaJ9GVRcIXUbxXexzxyogtVfdkIX+ox7DuXS8lBf3gg98NANrBWsAQI+Litw3ZkHVCNQ0t7ZQv
wImYeKqTuRTmBWRCivNlMwzl8nZbssQIicWemhPgagb0PBYYEPOS/5Zc5X1dYBjKYV3z7gwn31jR
Dn6j8DlyE8e6hufw2kdoXWz2x3eF8We0m10Q8e49SUUaB+UMqRXp68Mm4j21nLNf7am8WwfoYga9
MSlOWI0/GBPK74Uau3lQcsSPJ21CdAN/6nKoAMV6yLeNkehgZv+TjrZ/1HfP+i6MOmZ5h3xchkcb
ARddH1aKOqo3GXXbroZtuMC489ZzMmsXX5NgfdgWviRY/vs2ZojYenLD0J/dgJptyZpHrxqVcQPC
TwmKzqK9Ce6lDlZoL65nxSvw5WeJrgWB4spicKOJjdxm7ADCbYasWTY3ukHvDDHQtLfqwOIUTuFD
Zkcbczdcq0VX+FwiImzH96RQWtXOduiJCWX+BaXPpdj+WCsBmEU6/ET4EWtNozDyi62wnLXpzury
F/FBAqNhKgHa824SR319GI3egabOjl325nnyuhXDbNQhhMzjVYM2VcqhcA2hQN6F8yyvkaq8oIhT
pPjS1mfyQOcNonQVAYgLDGR0d53gf1e3xy7aOof8sxsQ2uW0rKkzFupa7Mpf47hTwebCNQj760/B
VzuOBoGYIdL+0VTTDsqBUkF6gr3k6jRTY7R3hS24AMw9dVGZnLw0zxvFzIczxgzkBuksgk5bLDi6
cNlewmRHwUTvibwaEvBNxUGHammHODnNG9pL5sJf3ipvkFa/YZwY3fgnhtg5+kyrfJMLhowQn960
xXsQl8nfvIsP8v0jJT3eoWezuasv4QxP7kdmQekY4iy22hlgT+4A/2NrZpBgkzMIH13SRNNvPxKc
+yl57BlvvcvL+sr3F4lTo0m8yD3Zog6lZ4WXOFoLnN1ycq/vnI+gOd5aPlC07WMNher1liQHk7Uk
AEuW7OIhEx5YQHr/A793qWv+JINuliRI2IJv5mo10YWfykYVXg1sh4KSiS438tQVSsppygbBbyjn
CSZZuBwY34DRMm8c6Gs7LnxxdiIWtagWnK2/wrmr2wjJpY8B34s+a4VhOEAo+ljuG+W1lpBThQw+
x5aruq+rErpb1lQGW76H8nX3HQN7zcHER0QF0kgSDrWZxKGnLraFpUU3v9cGmdXUaoozmJZU/+bZ
dhT/MwuHI+r/rb8ms7tyNl+I3LKgry9bMSQJnRHtVhm7wOWwDWsZZ49TTGr04Ok8ZaRwzQnyQ1sK
OKT5v/OB0r3+aOdBlNYwGTI3LW515f4ke4kv55qfhaolPN8atQqBMzWJx5Y80ktw7ZdsxVwl0xB8
QVP6voSdqZY6E/frpOORyi0ONVCK024RmPc23N6ZxbT2VOST0h58Cb2LsjB9rVFcTDmxYc13i/tf
HaPF2Jwdk9jHooXrByOlr7Zcxfdbch49jfX3R7OSid/PIb+uyvJK2YDKYVvAZgEj9Q+AmNUC6Cv7
hlj1SeO9h0LzIpVQ4oymHGbwX9kMDR3NO8FWVXOSWxnj6dl8oCFmbt709M986lMMa59wDPScX+qP
0v4XM+peqQLomBZFN5Kd0nLp5F4ESPYt9YVEq6gOizGK8LVpJ5tY+isLjVZi2Eu13ytZkE0Acqlr
f0Wr/nSOaecw8v6avIKbLHxhZdk/TEklu68hXqDl75aYjTGSOLqu4nr5GMd7kLFBn8+GuuHDMjjP
jukP3lK9dGqBmyVGSbrhG+M77wqOO79z9F2yzZElmK7Kj1QiP3Njiku8R7PUzNKja6YzAVW+nTHx
Wqr8Uzr0Rm7uLCRBtHJNf1/OvkQ2zx3slJ1QLKH7ztKXNVbL/20hRzm4HnsC6Tm0y6hVfhX9eN4C
FsyMSLyYBNda4W8N3ARu66p7xqZdHSO+9MEwjv7Vabt2hFDOXdeX+kjK2AihO9Ze9blqp+kK1rx5
+0u4CeLtyy0TvKz8JRl+7DaieQ+sz1JK4jjShNJLdK3AzIOgozN+TGk+XAWMkNAGSjxpW9haLZam
IBW5DmdhWwK0tWeY2BjOdCtDKHCOdoB0CIV4JqNHUtsa8V34jhZZM7aOaLNNh/qgfJgfrTOu7qQs
UuUhr+uWkUxolPQdzAaPXwm3IQ0tFfR/DGFkao/wV/irGIx1Gn3TxrskSvhG4gpTnX+vQdOSrLGD
W9iXVXSiZx25I+lsQBnLoEjZXI6YCVkBi2RZNJJ5MZ/MZwHonTwwx3TaTvUjJRv+4jU/RTOjfpSg
X2/kXemygBmBkSARnhRIWBSVJK+PoEmUnmMvSawqfyaABMHFqW/Zpy1xpKNunvZYc9QR1WSCB+80
C8f0HAXiIaKCcCKY6AYd5Vsvaluns84OBpNmylgOVGBjcJ52VAPhcu0EUKjktvoGEdz4HPvEyAW1
A3nLjxemXCq9a+quWf2FlwTa9MZqKFbNP1PIpV4WlwIt/LkrYrpqsGU4ITQMwX2KhHQS5WfqAiyd
AJhzfJ+MFWkHZPZ5AKS74kged1CXroZh1fQhKQCQPs6AXYOsj7b3Od0Fxd11UVWQel5PnGgvXhJQ
jOXVDgYiI5gXCL5c03nzLDvLK9/DVLYK1CMVAlW0HKPj5Nn/SqY/yFBntS/pzzdj/taU1DXS8ynE
s6uExHv0oyPyCAf4F+oUz6njComC8K3iavTkDlUslPPLgiEJeoPM0SREqi1hrDbi/ib576dnEpU8
wOqpZJi4v26DtcU8gyYqNAZjFfbXxHgxQA2Q9pH8DzcOt+/G6VhXvfUAlYCxGholEOLdPbLvidtK
MKMW0d/M+9c25Q9u/kKreh80fajMBbsPOdwmj3UVW6sTRJziooI3YPmSCXun6Gfp5+lDtfoZKWFp
AjwrJSl9RZtXz0IB3FYBu7CH05ss9Bn82ydJ0Q1ubmcGvjvNXX021pWun2e0eEpQ2DlobY1Cvgws
14ZPN99qeccZZTEk8Y2GIXlzvmq8OxQM5W/VYWMChNS2BgBYZIRAoXNPJmNhzgnrQFDheI+35ZDo
DpCFiNu7wRzC/NA2gAAD48c7hhVD9gIjt92txA3z41d3gvaXwoxLtAZ72VfVUYCjwJKqrEYhavgh
6cmzp2PKu2UPr8bUL9PYXhP5SgUuKQdNzK332Eel6HGKEXb1GH4zd/GyYNr0+PfkccljuhK7mOEa
f6PXfwjOywO8rGT0Lb1dVSTNymzWBdCTZlY5mxqIQN5oP4oOFLsmGXQ3aWBUEa85Rz1P8oHzkgI4
UeE8wwC668DwmIeDDi8C3xrGffRoS4AzSkkYi6RxZ6ArKqRV9nGVKTXcW1vNADOaONOTtMRA75ba
lrtZfpBjz5mNT5MkGwlrUmpdxyz0WoXi9wkP96K6iPabGzeNJmABNjf7yxVGGCLQv9o3GTu2e0Ce
JpN+btNZZOzXMdf1dOHkfoFc92PMBuR2qMwSF6pufRzPsvpGVH2Q3x8Aig2AznrHoWJVJ+dwkFgj
nf09iJ5FVE4CidA8O3mDacSZGUAE3o5SnklEUAGd3pKHaiglYiwRwS678xlxY06wA8KFGjdDfcGg
WbJIIpg6PIGfLWwx5EYBeE4WaPzdKHWJsXH2RBg/U4SIZmgKsbEqM4Y7YN8YaABUmKGkOB0qERUU
E2TV6soctJRPwsNkz7qWIpNYc18T9bPRkKiE9GKNrVn72T44GzTXZlXhW+mo1y3xShBXmrHBElzz
czSu/4PReX7vPLJZzmkrDeHv9yXP0CigJKbTqImHi/P+Q0ci3EEeOmzHnfsoOMMF3QDubKRhG55P
5SxGkgbcIQyCtym5rs2ickCyxvKIQhoruMDesuOwsNn+dVOrLffhdRR8cfranOAfmBU+3x+WCRJP
y+mvdnNjKr3LRmUWQJ2f9kG9BiwuQrtsj4Z8kjM9kTyjY300hu39c2TsMW7Q8rA2Z0ff1wC32ycf
eYxMAXoG2vQd/oY1UmqwiFOltYU7gJfN0RdoqoUS7VG4UKUdHoCP+7AALeMHH3f8fia/cWA0s1/G
Aho6jr9cWkOnAmrWBWRhqUhUp7UloWfNnB/sRvZtexVB34e2F1udt9IsHk4De7rKA6BFmJoS5v4L
u2TSZAjr51k56ymm5021U8+tQnqW6VdC79Z2YY/bjvfJHIDgF/GV87ccvBbrDW+NFLjmTRKP6PqB
DK+kXvfZVz2wnh3GSIMG5loOD7lr+F20CQVZlVlbLFulpOte3hN49xFtfGaXSc6yY7y0TwLEf51d
ysG0Sq/nyLTL2FQUWvmTyzX3pdN19p9oJOeEUq+zmgt4Bkc8ErZDF8HhMk9ToPkelbXkFk4egBCv
ofo6vLQ1f9xWMsepAyh+QKJ7myeZnCk5qUR2iBf91D2v49utcO4dDPb1lqm/eH3fdHEDo2DmART+
PPDNt8XCO29Ubq0EAJpidnkMEvPVz9hkFdiJe8v/+1nFyElaLidNGf3w165UkUFD0R9t5Q9KiJZB
33p1pyFBJXt2revvCUBFFS6vOf81zJO1tmt0GY8Woc6hBCtVLEioYZo+S1+slH2unQVa1DDA4Q8Q
MIgzNMd+gouGbJKg7jfUQ84o9NPxuKE3qULjpsEG0pk0PY/20aWAw3kM+UYzNZJxvuNW9QjDNIvP
jWOAN3Sdi8AzptOfKCSz47/xqpFspoKPqw1+3GabkSQ2IFatk9JOybqc7QdNDAyEadTu5NvApkgy
SP6EeTznEs7TK+UzcOJiv2g/awM9sUJfCJbxUx55gwiisoSHzNMgxUfj8/yfq9ipJwaLXn8KEaqi
k4Xfr3s2M5iS8MrdbK3FgSxOphEqoiH69oNJKcBo9WlHy60E4cvXppk6Vbs5i9PnwJbvnBkbJdyQ
0+E/0mKYXxsYyiBuNFw6+hLZJgsUOQUUdLAStTxc+H0HzyuPMzhl09RJHpl5r19txRFW2tedE4R4
AcRm75XbdKnI5jP6YIGP+0RPCW2oOyzNGgsW4aH1j0FRTqFCfmc0QBqh9GecOgpZgMUWsumN4VYk
z1NDOHazyV6qpxRkzj4hf5HYYw7i9lSorymjn+btvUA9KUiwABdEaGOVIDXvBbNkilDP0sTnF8Pz
bxwNllo45sGDPycuRy8wJ+A6K0KkkRce5FlySl979GWJlVUzcwZM8PMQuz5vAjJiheD+EFGbM6KM
8fZ5P2hBYlNlONsP1IGYdqq5gcn/eEkflyfSluUc+ln4Z9tHX26Cdzw5HEuNqrazCfXeTBYufG5f
JTk2qqyX+nEuICdAtxVIN5xEg+3ERtUIQvwkDgQSFF/Y87ANRXlIWf5cN+o5qtLarnlje6SbKpDO
RWWeXc6FFC06JBmsVObMSlMj4piuNJc/oN39jQ1F0aXSKz1XjraQB10JRBIBrdBGieZRDyTNgnP3
VXfVwo7905lLjdNGpZu25Jb7zCADnKuVY9Z9D/Hs+KQqi6aPX9LXsRNjxWzhVmjCKHJN1sQ14Pfq
E2D4vGOreIZPnaDVLKTX4j6wpOw/2BaOwIcWbqUKrIPuvJKUPikwG5108ejLuO5dfeFR1VErctMq
4yAWjL3nh9GdkvRFqVKMWTcRekS+PJfsj8tg2DtKYZqy+U9PMtWwegMX32Crf/GFN70BDWrVVdbG
OQ9C9/a3Lb9tZX4jO3ufdGYRLC3b1+BGlrkrb1gt5u0TJkyimFlzkX8kYszsm7bNomNSixFjVS4A
JhSQr+HxD1KM6XqwHfVeY04dVrr08NphvI6LLD5gvMSF+2sXnbdSnWSAQ7glnOOqbtaF9eaWfZR2
KnSeA/RaDD6E37BX6ETGhZ2emiUNqRc0HgQboB6HkPC71rYmcAdpmvrUGsJ6ahLVZCqVfoz5reNP
2abCXUZ2C4gUguFT2PLLa6hltFPa4WZgrkghOw0h7EZm85tvdZrYWDFijcvZLu+2ss3TGQZqAjjk
oJcnVzuqvGl1lcX73BGmEGH2EaL8LueMg1lCzzROoA6r2q+v6v4GXLLJCvD4rAbC9EXpVeckpTdg
sHSBBersv9Mj4088sLN0oVO7sw0dZo07V2JRdtJRNWClnl5RK9VP69cSvnvnYXaEoqUzjOXPvINj
3uOYnZ5DJ6OofZKTb33X9t3NUohFYdlWYWOcPspRnRAI9yoqV1X9P+dywLpK4ltB/x1xJdqqxOaw
F9fjZgeINJ89z5DmcGte8pRQzggZpSSaRMPtQyqPIE6J6UpZf2e2tE7APSNnfcdTeDu86rMGQuTj
RyOJMzWqj08p3IRGsHVbcrg1VXgMAOiutI1B9llIaAVzdC80hv0kFJInhZ07fW9uoyrcr/Sca/mQ
MdSxRJX2OIdyQwBAIm+7hBtE02geoKOhh+Bq7GujPssWry8f7EniHNK58V1TKeyp3Xl1rxszE9jS
nXFbF8w8h+kBJcYKFc0g5w4n0unPJ7BU2Wn7xZqOWLH4A/jbxY97CaSLfuap+XnuenZvaJ/oWIkU
NtogrYCifdizP6DbWDO9+n7sKbAx7QLbmN1hhFzGCItaRjdAVLTpLYQamAPhQOTha5pKstY9lf/O
fxyUnEn5TPWLXhXpIbRB/YKVAOUW9NQZRhe6eUJA8oyuohx5lMJ2U3LSFwgBtBeEj1hav2UfxX2B
MvGuTLtiR2FbFpjEStTpmuqK1H7kdhPMn8Um8MPMcJ7NKHXzfzY5i1smnv+WhSBcMwWH9X5qqXxA
Ls3u8o00XtW4RGSuwylzGYOQ+wcycZkbhgwj4MCB+I375tuVAOZClrVJABjR8R8LIxs+DThNvcoQ
SAlIuOnIXxQdSnrX9MzOxsRK4aPWWbDFv6HJXoEk5IePjgEfvwKI/PPvMVKt0hN1leIKFhuTxdvK
cuO7sSouUTo5qsSoytWUdPwE3/wxn0mVb7kDGTI2EXdjw21qIJL91jAroZdlcCdwIKy4S/OcVgIR
mgol2BKbh3kEKf/HenumkcEndEEbAB/8U0G5qmQYIxEY2mT68SpMlLHgbb882FYFuvhkkh6mkpi/
0EIcmLhnPG9XEBiWgGtdTQ/TD+9T0gRDS+7dmFRHHgK91lL10PR6VFyrttehrzg3L2CER6tHho4E
0ZfXFKbLWk//xGmXr3kTOIhCdoxQ0yBP0kgPuIBAaH6u0T0QFAvAMza7VZFBItDMF+LPkxbOHUhV
Fy1Mrwk7vmV0DjDLPuDHeFWt+kzFrgtJq9f+LOjtYBxtSqjMljU6A0IichLTRDcXnO3JiLUkAQj3
rxAyp5EXoUDjtcUD+uOAWleOTVJo066d8jxVwj2MForpQm4zwNwzPJcMmAgGOaFBRFgJ3SsTptkv
Spa439k58bNCeIjXKIVqPvohnVzA7xScQAvEV1UTO8A2iUXH/t7NnSRs+7J78iKF6ri1OEKLaC+J
RypGr3pj/PUvv/VHmkBPAvVpsNB+fZ44Y7Ykr9SA4+Tlxl4MxvmyZLN1XJFfhnCGCJc7mNQ+qvH3
ttMqyU63db80sTS69tmBSHV+9iWvAFKkheX/DJc9DF87T8inDbZDHE2I4vyHC4TmKog/qpYkTsIO
+aycHU6v6U7Unp6Al8j36/X1RLhxXnPP67syPiuQ7CFWwZt5BpH2GUFZI43qgnr90WWiaimmrhgV
mHGeSXX/vW/ijFvXe3UDBhuuUApVN5hRk7VM+yxN8mt4Ko6mpMXUbtVhlWHXDoJmiorULEHxPwXE
z0XTDnqEW/7/P/pvEn4i+MwjamEZsxAZycaPByZQZgQhUcRFvq4Z2rK1b1ZP8FaXQAHwtfAWuF1k
g9WM/DQr/MfAsDXu0dSjmKrFLumYzGjnOFu99/HtqMmYhOl7bilVDoCMdx/izG1g7Y7BCTgqKpIG
VKTpb9CmT3qEyYNOiOdcEacYHS3yp4amSzKQvlHk8HmGTyLs3Nxk2PugWaWCvltBmjrD7X1VAUgo
CwfnE04WcOs/bbJ1Yn14osDL3OmUKt65XYjt/8c3t6pu4aoQDcDnx2kmSZebg0SZZfhBxXQUH1iu
Hk0/SDlTIph59tio6GB8CsqbwYjXcNDff39w39QrPFo/IJcJRFLPgVFTk3cZNjN6qjBXV1B6H729
xj6On5/ejQVdkx23XmODVoKsoGnMzOYh6pNhQBWlzawGigv0gHb2QAmoPywK3d2nSdHn38+le3Fe
qK7pEJW668H9GCp+5E8HiUmB7aM33ORA7+Y8LCC2a/qdlLg+VX9lml0PRyiIgIi4+95ln17dPNQU
RChKxN6AIg0A8tNNCE1G5F+iUo3hrsPWlR4fMDdb2g5W3z1iQqS6Sn9kkbyZ/YkKlaYjF7jhBYJ0
h1f/afhhPFljw8b70v2J8qYsidMxkOQhvGy4xvCKdH8xI/3Nb6LoUhozI685Iy71CqKc3OeppQC4
JLhPahmVIzmvPRl/H5tmLh10A8OWCtb+JmGy5k8FP7qD4Z1vtUPBWRWkadiRintdne9zPQSx+CGm
GLmzcbLZArPtNo2OqWROv+XBOpbdpUzpSIQOMwO0bURohhqr/rTgRXB/xyfdr4Q34aS6Fii6kr7X
1cvc0fSNDIMBkQkO2JSlQe8zp+rLbO+X3vrP6EBwMpWVE3qa7Fk042iP/QT1hAH117EWoMcHvakx
EUOahdx60uwLJfpChhk9paswGYSv4icx6D8o1Tpocm0fdH4anCKdte54VI0sjz6EQhQnGGnTnFP1
aOK+HvWmDowZbSsnvyV2lBq6qphDVuTmFTgWTdPewF9diTN8RYBTFZN3IF7L9UyLeDw6MevJQDSa
96WvcvNLDCr6NCH4NWnHDDCaTfa8m0qVpA+3o8rAqDBmeAAIC030uhyzlNqCiThTIDHuV4T6mZd2
BTqkeiR2DoANZRb6anwh8ZTlXGcErfLmayjshi/sHydmmqWLIhYlUb2KJn8kI16vK4bMNB4J4JLD
fa6LqNb+zxGng5RfLg39VvAcRDFVEMwrFO4s5RsHjLr7NwiwxRNw81Kko/tckb84Ycbo9wnNq2VY
ofOO8IKiW9UcfPQy4lvxuufI+5pKDr3jzYMTtZeeCsD0gdkks9VctMB4g1BoIDNtSdOvKS2ZISQR
3fReoa0yvXe5escxkaGtxriNc0Zu8ST7mCp4k4rWK/Nlr8rWZ+g6BfgDuiwr3XWqLJzldl/L45u7
xKEWqtCVTJSOQ07gFgwe7BOCKtVk1n1siJHm+rwv86uN1245G5cjPn9gJLKzp2l98G8RzI5URVzU
NLHIyL9U1JDFAAfWZOH7WPtBSB14k797q9Gtu9uYtxtS87M4ZUiRoaZIoy5wgOZ6veL/J8Lo4Ulg
rBxGPL5h/mtuhsBkkVBUSbwYVgXFYT5SticuAUfJ+891Ushl4bExHsRbICZGSW7CpqZTxukEVNg8
h6eh3t3D2nQOJEI4zI4FIgc42nvI4ys7EWRPSYs3pQmVKlSmBUL9rsH4uzUjhMRv1W3ij2MsP808
QBzWOyLAA6vCQu54D9KBon3owg/18taF71W3Fmgoi7iKOR8Xfsf0Rt/Rf2yKLEq0dQPksKNX5Bap
zIkq1fJDmAXG/S/fQAlTDpabRe6lgBDbRHu8b2mjjb0FyMDz1wIiQkmIs8G2pOKSCSZFx4xJnfaw
Ail1lnueJI627BcRpmFlNvSCx+FHfy5pINVdyMC5+45CfVgYbtPFLnc3m6IE3ovFqi3gbNKKH/yA
nhTdmtOOhPi+OXrT2HefMJfLT+/OUjdtXTifv/Ow2ApVUcWZebiP5MrW3lwVQiHo6498TNsIZMBL
0rN5Kq2rR9yi08kxWXckLGsLmNLklMmsQfOcBfGkEg+9FcAhA/NedgbITF2F4aRn0BPPGvD3f4yT
eE9ZtrwEcUaybr7LIYJj8icttsGVrWZbGFg6CaKtVVncTpNoEl6Neqfecll06LS8TIC6rT6dAuOJ
qFp7/MNwY/70ZLJ7TZhfH9+s5aUjjvhnZYdzFXT9JiA2cEe6x2P2p5NNaqlGuos4QfGd1XDg26Rv
le2lpmrhmgQ93u6ac9BTYT4p15DfVVOBPXYC/qbypj9uuplY6rGK6Y5bDm0PbaJfnllqal3V+Men
d1mQQO9DuzVooTgk8qovc65dgwY1U6tC5GkpN+ixs7DmjhXFJ3G59tjEPTx/OdtZw5WieGYQ6bNw
plb2/CJc1Vkjw8h/EHWZ/ude9JqD+IjXe/0y4tmbup0b4qpNjE+S8E8S1zUYshxKrBQN/XywlBMd
L8Dhu9qbK+SKWXaq5cqkCHQjbI5OdDAdXIZJTWCR6U1wg/oTX0LQD6seVXPdHzQDcH2651NXmhGY
kCkf2SkjmbTHAgIy+Qx61Y+TiZ/lzcQgyHggqqpuzPgRtQLvwWJ0Wy3njIaV8nRR2MbllvLQze43
vgCt4e08zr6hOqgdxHHR1HCjh68BCO/3Pz570dt6pBPS3a2DcLqarRzg6CyPzpFOb6XGLFB492uB
4uH4zabu5FRni8FjcgJGd+AZ13QpwxvL9guxOHRGfjkQYrgNA3J6O+11pyQWjWi8QklZgzE5t3pn
IwXPLz9EusovvEuwXcJzfa31WvcIxQc2JDIsa40T9e66bTZ5cGQVII8wkSEKYEURpMM0zM6SmpYg
CZyCIehLNLOLelm2UyPeRxeZSWXLC/81jKCzxbokMMTui2nY66Z+M9i6OA0TJZHZKBDeAYxoR84b
goimIPT0gjc3TqD7lZ7u6t8/y/yGXu8xNhax7xqPTw/NPsoJvkdXMsRfvqJ4RTISbBELDRH7qPqq
4WRrWeAoj3SRHXEsSfL0salmHLBwYk2N0V3kyglVSrp7mlDj3Be9e3yiIbByPQiz4mwXivADNFn9
7HZuEMW85CNKfHYXe3TDLT/elzyq7piuz/B7aEZOQyLF41akVMuScKM/gBeebS5na1e877K3Udz+
YpsezDYQNRqXCiq4KkORnFMIZLNn/tSPEkWhRssJLCbkmnhlVfX/WevWpoJr3RKAUaGCawecCDBM
IFN0lHFsmJ6OclFj6Iwtk+/ziSithkk805EJ9Fmtwolu/fPptL5yN5sNEy3P6LsKUYW71ObEJQef
6gl7b+OU0kBCVruUBVc2dLIrcVyTxpSzJIcJIyjfTJAh531ncIXOUbsEPrYfKDTZwtosnW8i16gU
JcbkxKNSCWQCb33AfKpbVjzFOXGeb8HLd2uO+hgF4adLBOSNPs/0Gsugtj66XaqJmNaqioA3Ow9K
Dx/7lLvy4cvemWNSXY/DbG2MqUh8fa3Pdlj75O6kyFE9r2o5lwun0rJoAIyeAaihTNkjtSUZ0ogk
Nnh0xFZto1di1n2e83IsSIuk3tteuScjjYHlQiybZAlsK5D23BFe5GqwRFlp1KoymxCJbQfbPZDQ
SvXspyL4d1kQdVEL/YcHaVDd9iDkSvEVj86QkU6o0T3CYze3Bm6Nbl2XFvdi8wjsv/z+ZcA15CG/
HsguuVq9WEB/37HeXHj0TmPPpJYo8y23V4+dbOKFFMH9L2RKFdv4XjP7U0PCsbJ50IZa6cWKtxvD
KGBnTX91zonNXg59H7OWuY83Y3ZgN9BFknJ6MrAWYXUnn5vZcdk6SVINope4bgmcNKMod6WAmn3Y
IN21lPvdu8Hy4kLcdFRZLmyAtcnPgPraLSm6uSPByanqdTBDqGdZLjvvZlWsmkhg+XS1ehi8snIL
WhnvOhgi4Muiu2ZBry5ZJ3e7j7+QdsYUV5YZHhD8lBk4TF+mVS89L87PRFF0Brxvu6LcAgkNmqDs
UFJW1MhtUgFeQ560//kpkcBJzG3PS7EQJE5Q4ioHMFHdOi4EZYZDFKsUK/iQkZMIokJpj7Xt4AjH
y7hoTjNPYBXzcgS2QblQp4kfeIydIqs1fUNsr9hkJFRD3TPabdBYWLtcgWjs7i7ZHs0OS1N1giPH
S5/z30fPm+VjEaQMDrZT0az2O0ZaTOYUAUlz14c92/FgfkK8EctYz4fPsSZPMre8ENHZmi3317kL
a0PZLDZk5cgWihdKx2wUSDDZStLRisgdb7pG/IooPLmHKQuaI9RGdTF8xQxUFP6vKAUbgM5XlZNT
q54Mk/czWWN0Bs0d3qKGRhZCfyJgWdszxBPPNAopj/j8G7KwwsNDZL9SIUvOV6HA6XRMx4LtLsM5
nhqJ2ulp9GvQMtGehx7Y1NTBFOlP7epQoQgC0Gg6DmTMLUvugJK35KWEnwdvxQMhzwMffjB/s6YF
Fz2jBkBRitG7wKHJUoU3pK+JpJRyKc9TE1NbTsMd7qQEDPu5u4kzUXo+vC3dSXGgb8ZK+cMRl/F6
VHbUQokDKCgwgHKrzL67y0T+gEDlpuNHJsjXER7myYe8Ll6cAl8f2cXJzcQ0mW925+G8g9bV3vxY
tOg0UzM3EpyR4VIA7S/YDoxcZmdHzpIEsRZi1Sk6JSifUFSForxKl5NCJEztImI6NzGw95RNLqfV
2t3RSle5SaMwp2RlMdSOB77dHRfPjgybko9RT+rJVVYNEJ1HuPgAzZi0kyySiXg4zgUq24iZuGfw
Iynsbz53EXNVpFfo/BrrR7mLs9WcuNqXF3nJ7dSVYEIdtps8FkGzpLRUXRKYCnDgmrMcTN9xleAX
PdO5bbz2RtzNJT5bJabB6xFux4WaigfeFyx07Daze3muhFSxQ9TIXxWGPjns7UImnjWsNgfhEJjK
7sOOqT4pEhSmJUJP2HU24Cb98AGhFsCqAoxi0B0VRFh79Ps3JFP7YCNYAKtB2N2DlAjKo0bUEyAR
+Eiu92XS9QR4PPLgiXNgKDZzat/6ZslqEvWScpc8MhEKowh5aeZg8LbSzMdfoGLIsu9lo4eWShnt
n68tJcS2jisaMRP3kJcFd9YUrngcS+gON5ayA8MMgSTmQM3zbuH83xiRZ4E854wkHF5UPK0Hiq5N
LeJER1Jvm0vnaMWw+AdHZ29jIvyUDSJZUuWHsWLZvcM6x3lZ2sbgz+/vXbm6VTAQ9PYUrmzi76yL
qvoHeyB505/aNGASM6VCYwiXp+YTMhy54kd2NCBXSOScm7pWCsJ4iIATiwNsYGdR5U0P1eYmkNcH
8QlEpznlGVMM39S71Hiz7BpvN/c+HzErhRLIU4e5pnHLbjuz0/7yJ8n7H4TY0aAkhtUsFumTS6ZL
lEuUW31zrDJBBYvIhmJyr7g474pw/x84s5udSk4WACrv66tHa0ZlJh8ox+objw5IPk8C6cuCkW9Q
W9jcUauS6WEYLte89Cxo6qKExHxU9aLd6a/atV/sNHLoLJpxy/Y3fNCIkjOBWFqsBGQEb1RfHGDX
NMYshhPpT6VQT8MrZf5LkaOokXcQY4zxAKwx6ILiLO/1tYNt9DMDrga9kIDcy/6cxDcQJ6Fh5gCy
7RYtYNtCA1cSpRxpMUbozGfuiLgJQlhO1USRWuDWw7DrIXuS90P2vKJ4NwDZeeZsFN7HMGG8Vibl
jYFQSGLaQZqSXr+YjeGNhZk95uWJ037eRqaNJ2ugNuZ5gda06v6a4acb42PloyjFQ5NABpweUaEd
J9ooLbnsr9zYdmdBPsPLQCfDga/sbz/QHB0A9Y8ddjwwP6f9MIiuO20k7Waj9LoL5ixX/EUKWHfE
YUpcZymv16FMTXM0A9tOsN0gSPVWazalaGEu+UXOCz2f18OlB9OkzGcyZRTCXxhOZMR6rdAkQkMi
mkjWAXyI1uh8qIfmYlMUZafDyLFt7A+S07vY6UMrtWxKMGdhsWgyILCcMQbU5JwhDtBTDkVqlFOQ
iZlqBlr0h/QB6WE0+4lffi1xoGi4fpBxp4uXwcSK4+VP6/eZRS7GuBGDHm0v+xvukD6RNRQLZWw4
mKsZENMOkGAnPyiQ6B/+Ep7K9x4GlSUXc64WHrSUJVZTxGCDpk4LT6jMd6PPdc0+uiZV6e29zLQc
BsgMDsoNtenAs8caGwWke/dOUwLMegjezZt6e/2pW0S5QCsV7CvZ9Y8KrLjyeAxadniWNzqQLDmO
mVHdaAB02YM08cMV5k00gpyZc6RRyyDZmIGkOcE6fmpAhJhtzm6N2VUAlPzmmAbWuh7MDGvVX0Ks
9L3QNzBeHk6kzqZV0mNtkw4A+uRA2nZ0yXrISOskZTf5++CpuuDu8GjIl+m/UBuw3nxIVJUws2jg
LrXeeBcQ7wDu9J9n0ZhB0pwIDE7XX+J/fTCo4wAjKQeDpshW0Ilxjze5veVqkXI129rZPs2VPqwf
EIdeHJ7BhMBBMhUsrBgDA6zn/b1B/xxwXK0yIJ8bl9VVn1kr3xEY9uvhXJaw3d+KW0vf2znUEZxn
JqHC/Mjfo0Td7p/VKQeNBc8eELz65tegFz3GNjZsiLfkKoFs8aAwKZe2NEc51EXu7d5Bgov91/ji
otYeBwyjQRYPYAPROBl2RkmaniQi8hxPrOPMdEDa5AT6PAXlH4JUFHDk1ikbMdnbweumL4MDOAmw
ISOPb8oJClgPV1x9Vd6xGFojriRf3QmqEG/6Uu9y/n89/AtfpbXlTJuxuprSQxi+sCl7N9G9tbC4
iLZjwdA/+YQxAa5LcNwt1UDFCHV4clreTLuBW6WYQ3rTP1yWibtZTwBr8YVq24q3wWuEDxwacU1g
CEu8AdpkUv7EPfqkxYxT1EfrNeB8iFKD2IAL26zSnkg5uITvnmhVwOD4ntvBmA8AfpS+3Dx/ilPe
IYZPz+y8T8ZidLHrTNm4ZmMvdXUc4w2lXzld0Br6egBt7c7joEK6raLYBa0Ar4oya3VTQ0Qkz5Pz
0jJsXFpM0olZqQyQcf+T4E48e9a4kwwewaYzFr12+VWmTuBou81btfHcOJ9kmJujVngRS3vpvyWr
71TFAw81sAT0KsJ8yLNNcbd4UOC0n6atNhRQyeJmpFqJbJEvtqPqGzuBnKXMv468ppVp54K5mMXu
XPQqf4Z11fnLOaqnCMRfs5lrmtFxGfUceSkfLG6nKvh5iGEpAf136MddDimFhb+vziQo+qqokwpF
ZKc3pO/KZYNZ7k+e49dR43q3SDyQ0175AA+xwi0Ya1tMl1UEee6mABNszj0+YeB+oQebO0LqGiEA
c+QaVmPqJdRMj8VOvObw2G9zC587abDeMxfVmv/ZrN9r2jnYNStqBux3ujnrn+cNZV6uzV8btazz
OwdNAhuuQ5jEGYO7ScUFei8EbTIz2F7tVR4T6CfGQkcD3NIjKkMhU6/JQGOh7StgG/S7xqcadD9a
/13BRRsSgX/QxF7oaYfV47KSN9zqrwHLftVcBSb5udetTtbnSn9KGD89jNivOF4THxjRf7ms58xp
/vM45ruw9RJDrFhtdAl+tOd+qYMrqu2eg9Jn4HJ70Bc/svZ8gSMYysxz8rQFxx6H+KRULyH+7jYG
ta2AE4gH30J3XEgN0lNPu5x8/WsuLVFvnun6A5Qwk3bUCAEeJAQzpe+/mIpHZLzfOFcTJ2Nu3Rbh
1/ygn8ds1is00AvACqyYOQ8YiM612k9x6zugqT2QZFoo7/fSMDFER6UMW+NS2C7xKEwGkFqqOE9c
xxPDJ637JS8PAQcF/FMUfiFbwQfFFoH6xZI69mgso0uPR1xmHyWvd/cc8LS8syBL0UTwyAmaiQFD
mutbsDJ4rFchOwmgqdh2giL0nXTbw/W3JWsuOcLlwG4mMigit/28DwxLubxeZtpfKcKQiXBJpPCX
kZhXFtJ1DHGUcN4R/StZ4cslRDLh2k/yPVDXlWowqZMUnR6Ygo0xwWS/7juWFs7rzoUsSAbGZXiz
+7yTkVTAtt9FBbGapE29jg1Z1jPBZv3XOwx+qUgbX2hVMKkH5HpR+1Kq8eGInqv7SqoKNBdUtKVb
suN3oshPksCy2bJib7rEkjY9G/c0olt+36hoJqllsHVMLhjXmOZzRgp894qxLUqr9rvdAzGjpgrh
/rL7/W4vrWhzwlViJcykofWqxDYLi43MkNVJf/x5xeFCV7+ne676/gwrvfNWg39WLiwCD/RV0JLZ
iPWHfaiJ/PLuPfIG2fMJaFQyVfEIIUzcs6IwP9eC52XsIXWnf/0h9fsIBfzwpHMLA/pMM4a+eDSa
tWRHtZyHgSVZzBSG87kb6kjFnqo0rlEBjOxATyaJmiiySA9VTf9uMXUs/e3xwJ3nUR+TGP5JRTSc
aiHAvKK3hcER+a7pPN8HtoN9a3cC0aDtHYD4NEmCyIBPGFo11YjJ52Z378fpUJshiJ8ARY7KmmTh
mDaBxTeVNppPDB31MqERNIHTviFy1wiTkuS+VbhGkuEAMV4ASFKG3EI7Rp6fI5m91wUJRwR2X0fD
7mIIEwAr90WxxXngjM3y2B74RXAL2jYSE0eKt0G6PWK9Gqa7A2Qa1fB89Y+uOE5snYqh5in9+UTv
mEIZ0Xwelqi6bzArUnDzyNduFVt82uHPFb/McMAj6b+NthvSp5cQoveTCCDhh7t1LWtPCxo0imTa
ks3Eqaibjppd8Smlqiq7ZaOstjVY4TSKmdIjXZ60A9G0DIIYHp9ANOGuvKXVsFryTL54qaaWQBeI
ZPtHhy2Bsz8u6DMbkIKAMhYSLVIFa0JZCctk660hIg/gqf36UtivzOpsLHcTL/SUiO4FJPvpUJWo
tTHAts8VPB/YIn+2kVIV+2rdjvfY1FsLtqg9fxMPPJAloVZB9wOhmrDvF9fAmyWbS1asZWdigprl
Mo2gEYPVkdlzwYdKAwb/eLZyAwu22Llsu51scyBdhQRe7SDFmC6TNh2omhpz/jpRysb9xQZoLXNK
gbfL0wOdW2SokfINciyxlNkpQd33ZuVeLqOnA93gTS9PMvj8S0n9UNuomDktEicbruFgURJfCgvZ
3sFo8ze1cbA/DFF0KUaLsVMxJaw7H9wjKADg8+CgnQUxUj/DkyTM+tZTJ7/SBjR3b7FfdCwumzgO
3gLMkInbuTGerQ23X1jsf9j8VBkpEE4zfjN97ylJnI6nn4kh9WViuB62Dc+Q0jnOzy9Fll6fP1Zl
QkjCjC23A1pf/RFGhTFUgK4QlPFDq2dLxQ34hsfVz1Y/x0cp+kXR+BVJxnxCor5B89+0MnY6VohP
oRWy89zmt/3ott2pAhj8JO7d3Muy8a3TaC5fCKLqTZzf3QneUctZRL1eJiBUJ0f77T6VwSYirEeY
6rUX1Y1Aa6SOt+nq2qWOf6JLImNhY9bT3VNWfNfLrDsMa4qW9+k1+Xsbqqa3OkiZbUPXoICoCLY7
AAtqvK8WLUNCfOvefU+EIedz+JQ7qT0gMEW0LBhJX5S+Zqb23pq0Dihn7XwIqUFVu2u8xX6AKsHH
mKr2XRK1UoMOVB4aqKH+L24B3gRliBqTNp1l2krcq+k0nB5lt7+te81hZb7GMQsoZKTavqjQxcAX
7lxUj03Cg4oW0U8uYmDrn4/N5V3G02kBg19hSMDs1D5iFPbbT1Ma7cDfgN2KEqihcKuiE0/M0259
YFlkxodFQ4xW97OdBtZZfU7ftKVroVjG6Jiw+bMyJ8U0glAyX6bAthpN6PrsriQL1pfkVPK8V3Hm
InWDSWXioCSKZ7sNZTRR9ISjFXBulSO0W7WsQjOVDbvfRQqxvROpvaP80rIDGXYVb2M/S3IR7xr1
QrWdg4bD6dtfaaLTdPH0i+h5lFJaqz912A3nSXPRTpnHIuCRT9F5WLThGQf349IJ+OWsa4T4OHDx
uOlevmMtXOOmdHgffs9PnYl2hzcYp4MYkzMhrJoZO7C2TM93NvcT7fnIgu+e5c7gtEBTtFvRvGos
shIPljA5VpEfDF+kO+uoLqVy5ZbFC0OSmCLirbrDGDEJluhTb4WqltbpCwWzvvPxf7RZ5ns+5221
Q2W/TEF58EupJF2YGQr7XXm0s3L7gqq/uUNDfsfBOOmhGe3gw2stCCgzP5ZdDzJ1wY+HSLd0qQuE
BTxY3royWXKXNClp6ByavsnPj3v0w3Grtn+3fS5tRSGMOr9xd4wI35HGY6LNadQh7HXxrCw+dwn8
y/r+7YfVLYqmP8QrLByG7lbDCleYKEApHzssYplCWVqeQxz1QQXaMNMmaSvm2Zc2u8WLuyMHv3c/
B6LMl24984m3aGOxFsDkGWn98HHbZLTaqyPiNb+xY6HqlkJX4cooLoRJT8PkVMJs77sqZQq/NzEA
7O7rWJFsoZWPySyUmVNMoo4zSpBZPtByMvJ/C18/GSnufEWbpHOYkt4M4E6jMOLLnEjcJROf3O8j
NMnDsTFD5HAoS8t0v1jaOAVhCmJu9ECNBbMEF2D6R87X3X4294EvVdIig+IEtj7r29hYgI+YcAR0
d9cDeUqOVSAhybC2eY9HDI6mQIK9V2WpViE/iDmI4hCeUM2fqy2PI233j5kivY8/72C+DKX1Bk7P
N+YFbNNJrySHdcW01vzDSnIUmBMpBmIyXrWnAAYRJSdn30XIF3xzh/+zP7c41dXH552I9X7anpVg
5TPKJKYJZT50wR501MWOua5FEg0RCUvlWqT7gfvz9zha6smBWWmU/oH9fD6uU2KTp88RXOzOHfII
cBuoRWdpf4HekToD/F2n1XzKD7/5F2uUUDFHQ0dvvUXfi/s/0QnzuHkwya9uhvV79NjNSCmsAxfD
hbf90kM2VIxETp63IOgzRV/wAVfsTMLsqPOqefvNDmSkEmiIRVMr57cS03B5/+uH8dOSNX0iMhNY
7cF1Om4PkM3gfS38+sdiGMOfXiCKgoiAmyxY2jFm1AO/66ms+ouD4wZUOuMobhF5m+84CjoVZN4b
FE78/vF2gru4NlH1/TtwumeEbmg+hH39+9iOvxMnqJFyAIwEIyYHr9bfROFjvFSvGtjjyqbznfMk
RuM5Fu0OuO4NPtVDPlYOdpEbz8zMQaF5f1PnbNLFat/SHKlEarvBTp9tt4BlllstqteW/0lz1n9Y
H+HRXWr+wcVv47qESlrtoODo2CV2HSseJyrhfpe7fp0zdDaSCdZMXs8sdJKaYu9zD+TcdCMgjX25
29Qd3gExwPPfN8CSXtMNbAKptdSyEwbxwpBUzdOgzAGvmen5lsVefVkQGH/T/WunYEXiS1T7oFaD
iBgVfmnNL96stdyjfiougbzVzYRnkedXvcCXua5r8yQUgsHmkDyxUpOZjRsZYJp4sCr29GH0pLMM
HM2XajxfOxe9EnS3mgI70sWM2vXl1I3F5ycajKKalCUVK/XtYoLTB+x1T+FU4e0f7A606wTKb+2a
XbNvQpcultCsv0FXjYXG0B2x3DBitXKGDtr41uZvBBxjNHihwYoYR9j4MQh3SsoP3r9TN1lUsmHo
4eyoPaHAR7xfz/rnDtGLY1aVG8J4JCKqc9YewI3krVVOW2Rv0cD1dAIMk78+uwqQzUs2RaY0x9Fe
xImmY9OT/jcDGzqiaBS6VWdzBfpOfzJbpe0HEsd03jB0UHw8A2wgPr2FWyZ3PimpzUgIAZO9oZvN
GbCjOkHsTWaofrw7AVf+AFQYODX3H5MFS85iEFQO6uOaLmFjkTqYG0A1KXb7CP5QycaTJWFjJOZ0
R6+jsU83UV6vvx5Q9gIOEtzFBTiFbinY/mkED/uGcgfeqiyf0S4bY99yKaxYheBwrOAbmP5GpT0d
2C8W68oikZ8yE0m6F87Vb4R1rgy9dECIjioML1k0t51fG0NGpOzD/UeMiK2CIDWiQkOU+9qDJxHd
iBLsG+Abn7pEQa9rnmuZIJG3CZJfj3Q+JaIkz+tnuYYK1csSMDKTHq2GHbfR559yJP20QotrbiRc
fvDNnrjKPr85XQVRgdvFEp3lDXYZY/EMtadTNwpIPAguuAXJqOTbA9dq2+vpszO9R/WSab1NfpLB
D9UUNnBVYhwg+Rtz5dD0+Av4PCTO5MEJMiziecNDH1ms1r5v5fljCv0W12//nSazn9ky5LIumhoS
vVJxgF0SlfVM48cZQHQibTvRQWLG6+zgSLEEkh8xIz+46sC4JxLkH/X+pPqG4VRo5v2bk9nEuM1C
r4A1Rx9aczaG346HwxiOMTPQimPEK0OklLU6PwnipiWWaCC5Zpq5sGQeDZg290oSl2AsNlc410PV
DKmKljWuBBvfl2O0a0XjVK+940aqxlXL9cdmwx8yHl53TJQ3zNNzDle3t5upB6zYQkECX7x68VLG
KWy8istcXXdRUH/ydSd7I4vN03ypNs0Q4j+g0Y4a3DayP1EsP599ifhnvcHx1vdZMxcD9kgMNxID
wgRUkazverkFkfjzL4L0+OlNTCF3+z5N1xjsSn71+Av4WPHU6X/i8GN6t/DJNoam8sR/f1ZvT/v6
SWy949qQEIyIsR2ZghOClN+4vCOSX+KN9dqjQV3yqcCII7AbRPOusTWE7se11Pd04Y3LUh4qdImO
PZZH4sd/rqDiERdh4hNw1bwgxS5BLYKKINMYtjNmPUy2AWmorTFOXFnBGGnvxEK6gcGOJb0eGC+G
AwdZrO1R57v5t7i1UAZ555baj+Zt1QAkjs6ayiqW0t6lG+TjZ2T2DvmtwnOUYzedGFfmZLjfATHo
Sq+VDTHDkfuljBcMc0EBII2apubJ76aTJ4CMne7rA5QroOAbY1nCnT28qnUYHM7eYs0gynBBTWq3
KYpu7efOk3oJ/+d8rm0afY2OOSMTQj+SKuCY5OYIylTlr69YuZBGP3tJshtygu4P7bWQ15osaWGX
q0v1tKlUUHBExJiVNC6DE01RO6w31GNR8N03qbCafZ2EXtxGilo7iRfcqBHojbNRxuJxn6SLD9c4
mjH3MgHTQFZM4C1WeZUuxZqo/gJIgzhFzoxVlkgfgHyESfE2iLnxykFJPx1b7X4u/26C5h9cI+Cq
HfUPHqKu+B/20Ruloxx3NOViQbvrL0W50rUCj98bsQe+wOrr4EcI28Ni1DT8mbHsf4gkcD31ECHz
xWM3yesSROA71jPyTormOK41G0D/532UdiABKvQSzzM5wcdETrW5hUz1zBOb1Ofb7T5+SGaQ/E4n
YrRtklf+jNLzART9tf2mLb/GPAw0J9E3l4lE2f9S3s6VLArXgrqUFo7X1GatXg0FP8Ex2XPOEJko
KPnCLsSRlaaHC3D/IoNK83Brgshp4elaoXQ6w8k9isJsfuOf5sAFUjcv1pyKbE5x7n7W8QvY9RS8
B+EeA4GL8UFwr8AhxCYT3y3P6UGmdrrVLCTfGWjy5vYaF+ui4kk+h4JKy1jJKDHAI82V8TKCnsj5
4DcA/bkip8p4yCr5bTItVt1JGV/dQRxQ1UoVbzPChxhRvdFoTr4VtDFYOQVvYEVt3ZuPTA/xBqf5
6ZZZpZWI09aCCV/dNG/nFUmHh70V5ejwmDYfD8rbcdLmRL465QoBSMfkfB8ivGIxoNF+LdqMVcyU
Nfvea6cOLfHN7H9Z7yg1J5d6XnVQy+rs+8kOc0E0kXwevNodw+EMmUm59Lgm+AOuJiOqaUjvP6F4
9IEuQyAqjlfUEBMjcKEEwFA50ad+IKoGB3aQRsLLOMXas85T6xx45jDJiAjV5O+uBIK6tmPxl2UW
FavSiId0pDNl3cZUnQHwGmBzJNSu9uiTdCXAQ7FeMG0qjhHlqm/vW9i7JQVAqaeYGQ5JI0JpE5WL
nK5PZVgPyX1fgs26stKZchntOOHE0EIeimfwqXoMQHeRfIHFP15fZsz2+rbvnUHjqbzEJgTrgNCd
AfGzZbeuhVVTr6J+0cw/lv+TyGUmbxiREvS6hN+OJOwpamuSX3SwYQAfSKH/u5/OaHKAJFE2Sr8B
HnL55WrBX86UxxOZjr2DSqKwFqRi7ChjmmpP0Aw/5EVp6bcV4W2A4IX7NROgYGDEL4yLPfMFWWRW
Gr9FGbBXMmOHHMqFMibucBlmCAP01Br4I7AXCoBQyvMJe8iXb471vXUZMeVfut0RnWLdl4hqFBpK
3uXohjyQ81kEwqvqB0CIC1rn4Ks79f9w45pMnMs6JgaUtiONtvfUzY2Dl8T++ZSO8tt6lAZozzlc
1Scod9CplvsT7Y30aV36F2AyN2W//cMwCV5Tbc6x54NUWX0IlKX90iVnxHllVg7voAHGkt09+NKG
apGILZYNCp/n3df5wTKvCxOTyyXZTIrJyZwmDqc8ia0XbcRFy7/ObGnYLeK16N3ObQvxzgByM8IS
9PDuw9yRW+AXO7CTo/zam0dyKxRDjv+LYkusm69rP87JDRUX6rU/GktuxmLJJ0OP/Vr9G0RR1Hql
PXViJXM4zNFOUmDTnduqVuWwf1vq2SnH0waXLyWut56ilazarpevVoAq/TcPZW2JufE2ZEdo98HJ
XscsmF51b5Gs3CrnFlQGBkUO7s7JN19L3IfItoInt1Ex2Yan3W7AY3y5QrFD1P1XpMKHc6CaVoWf
Z0DBQcbF4u8lFyGYg2kGzJt+/6dY/PJT+43k8u7q1culVCVDCKPOn/HGr6shkFIjAQQAmv/tYbsX
hLX6VMrg8X9ztc3t3XskdB1JK7VVg0Ed/d/txboxiMgGhqKB4oHR3Vi/p4x0ZJdGgWlxW8tmAZAY
EpvwiT9z3qekaPQnPKpxtQT5yWPFM3qAQGQgt59qE2X284E4SJwR2lPpRgsLBfFPX7KY4g4mlts+
MwuOaJiLwKgaI5z/c19LZ9mUrTdrPKemsYTCZiJYBICIHqgIYLMfk2C3NxNno5aRYxQEUuwQmjW9
q6/sSr/HmgExHhqR1craPETH5ybrrGTP2ZRTeUqemPhJQX9yo6I8vyedIv1imGQqZLXueJOCrK9i
NPjpvAvlRS1HhJwV0XlgUl3K2pAbb3FA0I+SChUrAJRlWfugmYRAqU0kgN5CkT5wvUteWYzTxCUC
spqGDyoLG7id+6NHn91yNsudfda0P9qLEpk72mEWudlxNYYhYKIoOSPkF4Qd8SjtWnR4NMGoG4YU
HhOJDXE86a8XFKG5M2dJof4m/8BsKaZG8TZjQVPALlphBuDLhXj7t9El8f4NfGdDMDcUsZLGptIB
CkMG4pFb2E5qWSoswQH6w070ZEGGoF/ujcnpeSrzz/H9qdM6ZphDjX1niSavOTwF0XQ2jf3QhIAb
hnmVujMQ/hrDTbh9GpiipLXTAwRCcwT7l9XLEGqdo9LE+0VyIgLHRlwmlnWIY0/o4W11WMj4pDIH
PHh80A8++p7cIRm7dG5J1F+eifOdYe4QdZISNOb+0uqXrn4WHeSBv/C2GRQnIk3ltQErBogqv7e0
VXMtWN3G3DYLzdjKGb1y8quqDR3LXz76cOmZrw/6hQbI7o1y7WrxC9FJ4PjrerINFsztdft5XCUf
e2Zr5mkuajklde5mL2PxB4pGCXwoOJLTCMvd2H7PzH2lL4RPGV8YZG3Xih2wu9DjnpcbwQRdLNiD
dK4DTqbLLyadhGTdngFwJ1NxWvFHzRJ7Znwj2o+qEoi6yaDuh+TDeY3Ya7Vspk6xdCP7ZrG7+NSC
XyQNXxztvKiRhasLDv68sFVuIj0zymkwHEkzY3mcPaRVrdj5CGqqelhumGEmlzLcTAqv31FmYLHk
THOx6VxwBwX30CplKfXq82CQHorNw1U0EJ7+qmajl4fPa509jYKD7vTB5mvQ5g+h0Cawyn2yDutX
bmrIU6TllH4Oj8MDg39GB12GS8RwIPsp8Hmkcry804eRqFDx69nPvxWPxQdV74hWCGgKkVqo+ftG
m1fbqjTKqeGIyIXVIn4P1gOc5UGvgtB3FDR0Af7TsZv9cLub/NEeeGV5ZRsWkcysCUwn58pBl4FD
qLD6QEm57RGsapozcRXcadyaOXNwuKbVoqY6Irr4i4q85lfEyk74HUNW0UhiH7yFP5Juk5BLcRrv
jgTQVHojOmlHOXyrrz6Nz+imOrco4ZgGq6NEVChUcZK5Db1NxVoCHUxrYX+7bgRB/a+izEpvf2zV
I1rKyHEysigqI593aqNK5wSfZetoE4IMWvEdy4c3PbXr9Jqp1B2H3yZqdsJ4SOuNUJhe2eF69d7j
FuOPfP+VVi4JD89eVPiLF8l5MFkJ4accWmg36uG11dIJlM2skserFHhdNXSHJ5bWtrni8sb2ZgEl
xIzu1dmL6eMJj4/jRsNzarywZ+doTbL+CLEtSo0T0Mp0Uts4FNvbpuQu9f/mbv5a3o/yKfthR/+n
rGBzXa7KTlVrhJBYjO84X/D18wPm0axAVhPEsc1YwFBOjPNx8DCc0OSiOU+MhaZvvjjU/zvAUAh6
HMMzI52vdY3WCKI9hkxk8OIUAfaBXWqpJJP5w9pVkn/tvDSKrVmIh65Q+kXZlu3YJb/WRiXp/NUK
e5lDZBzQA+BiPRPZCzOErpsRDKbfGKMp0FVMGDEIFAYl+kSAvKYCyHXV5pXey125u07sH/K3fH0L
DNBozUcNOSCxuPT5czVTLk9mrFJI/HTM0LJBMK1LcDnBoPJuKyFim7jcjT2HTzx+eit19upoQfya
VSdFhcxlSg0GQHdNvOAJZl8Y4kC9zR1fztkCsf8AudpnRLin6+VW+ikeeaxWffQ18i7jI1q4e4DE
2DLvEilc50+M6wkl7MgMw2Qgl5qC6hq4mQE/zsYN5Dx/R/Fn0eSC9cD+mI+t+UaLGJi45P7bg4Zn
+XoVQRbi5Yjy0SaIsTqyj+tFCkWBv5/HCj/NgM9cGiCySCiC/SgQxPpo3OhJFeDHMOyjR4SGcpQO
rOSO0mS5EjuiE6RbPv9mYqIpyr466zYdCDrM3ViouLhNMf3JGzbeo6OP5ekoSc8vJzAjeu6DqWBf
n+aP7QC3NIw60nXoBhl/necrX2qjgSntOgJ9mksKn8LrNCZqktOSsJbW/VEbFrcLcE4F5MjKuzJY
XibBz1k0SWsk/xwBGW5tFE4eX29hBj2rgICuuYDtAZtznyUyE+NurWIZY9ixsUsey7E/iyKbEZFH
u744tpYwGclOMzZjejr02GyYz2pIQKpKNhQ/H947Gs+mbmfZvOPrAGmvdS8c/bscaEfau0q83Mqi
7dUJlaI+wdm1r0U8AA2NF4TeEIFgWLRUfNB4sksMudGk1D1UhyYZKMNauQyQe8kVI/keS9AVvs7y
RpvKTMa+x880/raOp1+BGZIR+8B3P07yxpUlD0JxFJeLznD1IS5f55Ah8ksYCRpu9Npjr2MWtctn
JHJmt3MRCwqpdF77W+/ia4as9KCGd7V5UxMOg/x+40hrQ6aiPL0+51LzBVwDBYekA5GutJkgTU0M
hFivFbA1N6DMWhD7Mx7fLo2Z/WqgWXosgZwWP9Pvj66ajvmS1xdROk7PYc5uLR1/tXcfnigboZgQ
xDwY0iRqTu9Y6sxLVE1VZNKQPwJfJmRBKBot01GOwchHPdEhSmrP9uXZqWqUMAuEabyzbu3jgP5d
45KXT0XwklsBALLb+HO4L8rTx9OJQb80ogboeaoRWRNd9e9jkBnsFFBthDYdDU149R4wqdrkXnFe
CnH3+WPS0DQYOQ9MKNKyVMdVwfpPFXZsqOgz/99QyysCAo2/vDFsiBC86LePpZz0WMy3WPZ4cY5g
hYPD2aNtKWAjEn9JkQyCqsSSPfHgMw7xc5L0KHNqrt5oiCwDnapykFzBnhmcfi2dgcCMcepUAIEw
Ad5gyMba7ASGk8j7nknyhFwxIL94gfHAOnQfjBfjAUC+t4a0xSlWmReEIVJixUNdV6ExidxcDSzz
pAB3VEUwKhUtupJ/pT9UgME5/MPiZ7gkTebAWjSxyhO3Xtp/VX1Dq6T6YbFW7CRfK16a2OWe0RZY
r0oCSvIb6bLfh9Rtd7qRl8T/cI1fwhZ5IwYfWBuDYvh9ZUszmfXNk7b+5GXDt/BVDy19wTYMwY0T
+8wTVIJ4lVCoTL4oS+xj9LpEQhMZlGKTcXW32Q1xDsqAQNR54gAFT2320JcsohVd/hgO8bZQ4Jcc
L1EPSMcQFf2s7LTL05oJLwe/tmuKJ3r/4oosYvOTXKs1IMtxVKxS0PzXn/ZRpNVnYE3fVVopq8mu
+CFNQts+/9gqqeXqMXiqiujYkgK/+QTFx9bDvINtBzsCxkEL3sz+SXonFtcq1pOzFayIrn3yRMWB
mFLOSxZzzOrw7FE/NI+6dHUHMtOdiTyaY/0vDe+CCIOCudOfV4zqmzAWqN8EXkLGX5Tad9V5oSf4
GblI6hEWqmuDss2r2Vyg4ovvdU3js9zbkm2Xi7Arg+i9IFw/AuQNDQETLjsiJfS0uCGugOnsnpEl
m3KsYZcrSsyOFFzuocjC8ez3Kp+ARap6Rz89hIu2drNyElF89d4amg4Yhd+UbcbSYf2dO+BTFld5
o7US08YwflvE0dpatCmmaJ4XZMz4tbK2XUCqvAJsdpsbH2PPEtZGCsFW8KM2YXkRc5Wa1KOF/Teg
KfuuLcPBhbWicMmCP8x4bzTh9VxxKFbg0jIhpTCUgAwNbj1rmqc+gtpEE9M30wt1oW2a1f9QnCJd
Ev5yNW24X4r28PEr04WgT0yYHU7zB3cDq/H+GvODbfWS4GU77lRoOqeTCr1TO+JV3zh2HayI+/w6
4zu8+wHuRkgp8e8rXhlS2Dsrr48s6wnUv1lOAZvMHOxCjyAILK86gP8iexPBpHf6/RkbSLRzczFk
fIJ39Sy2tTGRs/pl3uHGAStpsjBZF2nfsCxLgNG1Wx7KA//0M8hT1hEC5kuJRbYwKkkpgiTAj5vs
TN967aDe0WHp11BU2/xQE1YmHamqgKcm19J9sqzmoOShxDxWbGNESPFxUUQKrasDnQh4NVOS9DKT
Lg8hLTVcMLP7jCUNwaLz4pJW4YOd/ScydPgJm+AXuPB9RSY72yRuPpnfTYW9OVy6by63byJjrC7C
xr8SITTe/7LTkrEt8AZCKlf0EGQCnVbc06N8JgV6qLfeF++pZ6ekMnDopLzzU5lYb0unW/PZSfZD
mk76G1DFJA3EgEuCzyJXnkL6A3IGC88vUCWp51lkwvWpkV7+EhNigsMirVpZscunNVohmCFkMTHC
KnPJv+yDIK1irlldN2qRJ/zCXNUJEPJ2Onza5aLLjCPUrEK1ht/+RiDLGY1xTc8iozCDQCSe2+jT
ASQJuMJYotamD7JVkVBfXp+EOckWNhLmchtnAAxTqbJ3ir61sqOTZ8/M1IYw97o0SdVOkpJvQo/C
DmY4bDKVKTfsJ2fHzZoM0Vel6XySp2DNz64LB/6z6Q1rnH2n4nhupbP3rgVHXoGITgzb5QjWodbi
1SA3DjKzRwg1A1g04Z+Ekhiz1DIrnVi5Wu2SqCESBpjIs5lZ/jsgemqRcZ/vB9J061tkp93Gtjol
5iUoWXsCiNHkdelOKV1pcp7OWAnVQVxra2Amau757IvUaaqoEmMZCylDIF12YVlEOPLSIRc6Uaeb
DYXEEgZlHPGzU8GRQMObC/kFMiUS9laI2DpVR1KYPVIfrENeaaVSUp1zZ0UVjI8BDUlh5a4d+WHt
+RJ7gVXTLuH5LMBA0WWQ4FylVYgN39tfAZH16QJN3chc+IOS96n5pNPLdS9WGxufv6SsiZux1fUQ
gjTKONeOE6cXbIm4nLePH5fV28496A8SiGK4dH9m+zBXX958fT+AA6PGpvi82zZIhYQ8wwzKplHG
pcOJqDFHS/UClKnXATkcUTBYViqGxeOKVYrYrhDWyyWcLr5mJLPFB1LMSke7IvL+rge4yztjarCH
K58spXkVB2p7zJyqfAOuY94BLop9n7Ubrk14AlyZycHTYP8b6f+Dzsn4LYUgNozBwOJ0t8yWfmpX
R9RyihHe/EC9NSzza6xdYVhY5uBH26cH+KYQTQ/lxyFt8i/iT4Q5fldW1X8afiibhuZ6Y0+U7cHV
g/CU6/KCvxDG5A9QqrdDoSIw07nnDOtgF123WCPMDBZ1xoHzPNe7s1gmeIlLWGgnf5IHwDO6iEZo
L9R0zAFJdRcbmRrGbpHW53W1EveA7aDlg/Dj5p5fjQO6dEtnqbJj0YbHXjmTz1nKXEYVIDgLZ7NN
Lsey1MA/rk8yve1/pv867agPTPxEmMbpCZxGR40wFSNCugYYRK7n/9AFMQ8OnW7t3BNFTsoFIAH3
N50+YZIXFq7iNEWs49LE7plKgz3+mHJmx6OWIpyc1G6uD2xYB7cc35gbxJAqjc6BAZleIgdQDya9
NBzwkjW0QiyXXcnysDMkRKZjssgaF/ccXqf47neDSSqG+veFdPhyHuqpinbJuRECw/HO/qvs1/Ml
IfNp/OQgrpu4PBMKA7mjIYXM+vZ1eHZ057q5zeG6YrZebTd6yrJwFEhg0uqgHXEBWj6oB+yNTbJx
eguBtI7NgJFt0ptxjFRMbIIJqK/70eXxLaEUUX02TbB+i3skED0xcF9B7/Zc3NPYJ0ACCOrWREsz
xTIVM6E/2S2lYGHkTHlb/r2gWwmyO17ZBAMIb7euNCJEzgMphWG7QTGimfPdLf01l96WYxkRLo07
HNFyqVeVQGkYfLwL2UkgIQ1NfZXmaMWH3cc+oYQ1DkjI42cJz7Ad0zFmkA5WiAxzJFhhjvFhn/ev
AMnJXF9JOI8Vb3u8MzM7Vjy97fWHSbjcdg4BPQ3/pwb0GIfj4yu7D+DL9ysn7M9HMuljG4H6l03B
lxstqQhOc43RmivuGk6k7jT8L4gT5NBo+hgnNM/zO+bLGaeEwNESulS9DnoM0Y3ILiJNqjBzx05F
zc0E8VQ3kCML7c6N9/ZSbQDmyTMsuwKfZ7bGcpepcxO0ZonSVMM4R2FC7QiUzMpdgGM3nkjLIjI2
Hrbuhi/f3G0uhdYRGeDthGqV1YX+yzX8YFnuqayvjFDBdPRKKhJ5I4WH8UsDJpyEYu2McqRhSjP/
4MqPv2sAil+mvBAkC5zlKqxCD9Yvy0/4RnQkCXrQU24hY+L1i6VLiZcc8TNKp3VVMxt8pZGY/Uyw
ZOzQ1wW/hHnVBVDAtjP29rx/2d4JCQ2cct2lcwaNZUbfokMGlt/0Kbh99GqbxLKM699qU00k6Bsm
QfrIUR9/vYLPvI3pwP2HmU+2hdmo1kqyOD6kSBZsTmcxEe6MGeDw+j9quI6pTBvXRt2/owFo4+02
9N/XcWV7n0CdWTPm3+Y6JakByGvGGs8ikEWor9lFLkjzOTpE1Yq89h5P9wbgrpnjE7IOZarRY5eV
jATTYE5QarD/JDAydJuixgLZs3NFCpWXnj6TzDMrOSA4y6Qbc0CLQLU6N4SOwauOGJ/T6szPZDrJ
wYpe4RxUgZMin3aMO1JmrLaStlHCWxCejUUDrgpAErQ/Oq37oe+KuPN7U7vrtZCzVSIcECDM7tWG
6Enz4ioXl8iA1F1Xp9IXu6eaI2vfhBv+233GVYYcRa1DK6kTGQ1FxoTUSurz3V3uq320YFUbBhft
nV46ZgnKefi4FWRsoNc6kkVCiIjgkflmP7PSL00jIXC+kUfmng+V3J342uiRGOAI0rLu1fNuTHDN
Q4RLRObMQThnKWk/IZzxqaL1H3Iz2RlxqQDvbXk01jil48Z32fkyYqflot1K7LwL1R+vlTiWW5JC
0+IIqkr7ILDPirXEKnnstvMTY+IycZ4mBbl8UgtrJAaX1CYvB7a6FydJoUU/Jsni41RMybTA5On0
lNWmqgUPfT1CEL4iv22lztav8Trv44vNs2kAEufrA9AxbEQNdQJAkgFvwacP8Lj3rCKyK1TLybIl
dmuyPdQEBdW2obhkiXwNVRtWGbCyw3o4c6Y0bLy1X99FCCocvT9mwD/eFUYzuGV83OnZ2BNbvJ6S
Q3vL9c0e0P0AuP4+417v2Ki65xEBTDqEQLSR9Z+GHIKqC253FTQ1J5DQnz/ha3HxnDnAABgdlKJI
MiFmMK+txzLCYkzyOR6iTiUO10YVZTkrM1yJ1ax0PzqI96JXIfgboR2RjHsmmS+whTFQJc5Trjze
iLADM7PUvtGhjRHadxmC0hQiZAD3/6cZq50z492fwAkIKOLXNOufCEFFfjjs5+8Mam9vidZxrGeR
vmioE5opxb+rA61A4zGX407gu2Z0L0xMmancEAIqpNamhaaFsGBpSCz2S6m84mrstQ4h1oOuxdeh
Yhi0DKwtWTMtirPwO9Gm0pmHzq73KkbIPqEWXuFIeQ2gENoLordtA8YC0n9X8Wuw9OEFu2q2DuJ/
8M47pPiBJFtRdU4SDQbZZ37cyPkpGbHdgwFfTqYu+QKwm2xkgI/oqtCOy/PM22INISmvJu8KZmtG
AVkx+rdBA3mkM8LdrCt0nFJIIsFK8UQLj8oCMAmM6udU0JT89GPAPAqvIU0lfjW98I0Cum7UZ1pi
MfeVh1lrFI2yrsaEefTF+hXMmkhi8kOPqrt0v4qHy5VlYlj4/txEtYZfRCpFxReh0S6XmZDqJACB
a7zez/Gzz4txjnwCUQApRsyQb1LFzPnmoytiismyIJFUYwqe5xZIq/5vHVe8omrTjy7iiXtNjzn2
T3Q7BTna4D7/9c6mACMyNfthYwGZ5YUUkWgxh0VNBwQMjVmnZWZMUusDZ6+ZKZ6/0Y40NbcNJ10H
t31Mh5HnGMliiNUL6d0liSJ/IgEbKHIg8hl/U/xFEo4KvekDim5ggPSG0JKixelb/NwIY+58B180
ibEPNYEiA21fXTTbA/6x9FO+oQb0cFytuajRBYvfz2ky//F0q4d22pmwQwpkpwMic8t1OkXzYhUe
uy8HWlkmmqGOkrv+N8/2BxpMK/hKfx/ucMskAsErNN8wjxc6BDb+OWaJ/35RjS3fUpRTmOgNMO1I
J1ZAqSnRHfBqJtBNxEcJhGhwJZKH6PrT1lh5HD/YCYYNUspzAERo5N6NifFnrqXIuNool38UlKYc
8M9GsABmzm0jURgRjxrslsM6R9/GoNU01MG5wb0HU40jqsXVz4atJX7WI+hVGe1SnWv1iofcCJJY
tzZEdPoYkKU0+U+mfOs4v2ruqFQonhKr/++o6H0XxHVtG1SFJv3InY6rWeGTkLnqvbqXJgg5/7CO
quc86bC7GB0wPT0VCAXg5IDpLvdrKbFgLy928acl2u82hCWER6EZyVIvp8LfWaCk9/T/79OZ6AWA
J8Qx3DzNwgKAJnK7eg3Pkh374cZxJG5rQyfSVPCO3XdM7npoPc+ILeh0Jl7Z8gEJvUFhmMiorrdq
pEWYSSBIce4/yBBjMlSOdVO1RswZ7hwFJlbkGdpIfDRtbDAO578pY1qPPRLAogHlfKMpB1ODlcbx
VRXwXqDCZT32ANbJUuysIL2hbZixOLKnUlxImXj8t5NVZewBUy6fMyZd0vYLlq3R4HJCqxlA8v0L
03bHEf3wY0cVd9RNQdt0wY8LHzrzvU3uxKb9xDqKh4HKgn84xvOS2M+/Y8nhL2XHUso7cc5AzooD
jqwF4G2sQMdcROl4VInBUv6/dnWMYbHdIPoxB12+TWgKQbxkk3LrFlKXJa15/T35dUKinCcynfqo
iBX3lszZ6C5K9Foy7P1QQXDB8FMZTnWuNW3R8Zqp6B3QkJ+NGfTh0AomYxeIQpyLUaSQd8BId8OO
Ct4Wp9xNaMKYox3YysZDugjjaLOAx+WwJ4ClTvLpwZ6/qQBITUDfII/1uSjkVt7fb/7x8po2Qln8
dZKAPXJ5B4GK22HK0cdspEWmn5v5V7wLEzAERL9ftr5T6ysRsskmg2y9HMuouNPK9K15TGt08WUz
f9luPH2hlpJlHQ/acLQlsyGuvqJ54PKswehgjP0n9xAJ5dFx8iV30UMAp7OmnsRVZIkC2aQM86Oo
L2E5JA/kr6OO5Tpf+a3nRTGS8XLBWMkyX4KSXzAUaQqD+ea/Vausgn/3paVgiNrW9ym8FsYVsns0
WC4UMgSNKB9iiZ12cVkCHPxz/BuMU9F3uZakpICt2IX1bi61JJwjoKKFTCcOFjelzF59rtSX3hIn
Tjs2xAEEJ7ANE5EzQ5zi/Wpzso4puFTv7Fy+XLpqsz1ceY3GaAZkWv2waKj4Knmaehu4xeIw3Lt7
IYf5lRvj90IJZF9M7CPaoiu3VglH49WHMjyUwLxp37MWjrtRheGcqIHUgnvowRqUCzh06N2nidgo
MkPnPNGUwDWMMnOViBdswhCqzy+LbhGIGTbK9opUT6E5kOBlFiF1cKOt7vS53uVfATz2ngtVc31v
o/Chyo9IN4SU5KArLD8lwuKLA1lm+PxUgEDt6VU4Ak+uu1K8EA3EOoEgsZBtKU9QJHe23FR0ZoaU
UfbtMxEy8OCokcVvqCnTlF1ipT6skfaVkL5URpc3+yN/T70N9Gm3yf4i7jfF0pPCo3ttQAzsR3RP
Our8pOVsXeO/6D3Bdgzz9yomJSngu/AhAwrf4GxDfE7hlgP15VU4+FkOna232drqV/D2g/r7b3uP
8ryUEJV2Qbp6MmjRhMQjZaYI23Uq2+bMI3whzXQWP+lkArftRL0On5UheHFC7egTlKBIQv6tpUOp
auqKZq25sTZKiuVmNGLTIlBRVex31tB4tLJUTXxWgRRVkJHXBus7i5wnRKZVKcDm7XfdVMDeesjZ
hOdpkuGwki3+yHXxRsjbUDRD8lILOs9HfsXcSbAG/cGGH2Nh70n3RdbWN0Upp+cKNdPbAHqeSOIW
2OoZ3BIWTL94Mkhm5/uv24N4AFx7hmlJ8WmgX1viYc426G/iIYwmBl5CyKmCTvlvnsbwzW3iCJKj
OhCACXmjWspvmVynEF6S2zX+HVH0BFrsQ3M6SmV0QJrJ9T5+WRSm9EytKu9cxJcYQrx7QYVOEDaV
ysTteJD7vxxXyEbyDjA3AJfIzToFlZNJxiCj7yLO8zb9e1n5WimumQHLHnkk/8Nm7Yry1tHjbHL2
tQu/u9u6HJgvC7VcjLyhTzfN8/PEMDiroivOsd0sFvnur4oZsMYcDudXLIfRVNXkgIobmNpkeX6p
t4nSFDkiDpzNctmkHSQveIbfeYngL347BFh3SdVZ3VX++wuYPkrDctPaelYc7WrzbCviP/hBK6G+
GVzcZeyL5YToJCZk011He+cIzTDelogJcd39qfymdzJPHw8jJ0hciKRm22MTby4/FofBUICJRkxc
2FeuaI0m/7l8ypcCGKSGAWYyNAyHVQQORH2z+D0WKZknrBJblkWoJBkzttmjbTcG1x2s5trLTxfp
kACgy2AOoy9Zkioh7JWXArAnDQafwqnCwbjRnU+9gW9fvPoZtXXATct0gxE/4WLbci8pEK1vG0bB
rpY5njWzmwDyAalEuUWurxO82imOg2qv3Rc3u1+oAsbQmP+T4ffwJUK94mKEG82MPoIg1JB+VlNE
cBJ3q5NxVQxFvARdCDI5QOFLEtiakM0aEqAqr2s7nsmxYbsTCANvrnYxhKIia7uppkdtZgf/Z8yU
vKNBeCkef0rnU21e5yU52pTppbtbcaR/6ChYlchnWl0MMj7zrTntU1xGKNjP/91JxhTRAOd6Xdt0
XMvMjZyUZ7+1Je2XwTStxKE3zW/2dJt9oF2dZ6AYcx+K8Yyr6uI0W8fJRakfAt8bpg5RTCq+S/qz
dugPnRY496uai/vGktHxFL9s/iqqz7LCNgcQUeQFzHpNarfcZGZUg7z53W6CjQo5XuZImidwDGa1
/m6uhU5KubWNDsKaaXkywT8+nE0J9MZAUCnkDBSzJ70Xiz+Mx9JegpS0OZoEt3kQNX9nq/eSwJui
LDyxmS6Zh2NEprCRMnvrjNsS0/6tehNffkdzdgrCvt/IaZY6Ud5v592kXi5h7BYmQIv7AOzCEO30
bznzrzfnxbNci2D18NOH0PMj5Uqf9mYhh1hcQ5ey2UTm7va/faZ1Qzio51MXjvNSnT4MGcsyf8aE
ZjaHpfLd+HkDvcUbsScdMEN1OmI2SoOSPw6EkkyvCjaA877oaETF3bk6Ef2yMJkmQQjOFgjuM+0G
n2EwCosD6LnTDwDDUWJKMnveWG5jBWr9Nk8X6PjgJ3uDS8LKmNzDxCrDn1AlRl6MqWSUQjRrml8L
vWwTSphkPpkjmcKZ5wXHoJvxigV47fMEIafqiSuB/zcSJU+8DwGuJbEca51hKhH7p1lKcEdS8I2o
GEm15kcsMpJ5LeRcwj677ashaBHixAZCdGVbXxmiFY797zBCbOSVYs391nNNAfdj/GmyNDQeA9AM
k6qaTf6PIiJ30TikX4dHSLaIhIHGvdkGXabiVHhRKlFu9cvK9kTzuCqm/iOfM6Ca3yhk2nJFDIPM
NSSfetb8RaCWFHfyeumBpGlndFVNvV1Lcl9VbUbOCQ5L42OcLxfgHiEty3Gsr5hw2pMhvvPVn0oI
LEwbZ+qEOjjBVvGRMLzAnoepq7MJ0pz5ywVRgvnPYSU8Yqd0Pk41zloE1jIOxxHMrXMo7lNbLolD
uLFs4YUUIiTRuOr0Ziktvm0qtqNuxOpmnfSmoRQF+xNpaOucQkpx1at9gDxpmvXtGF6/ssowUHr2
Yw/kPSqc10n/8UQbRuX+QHOYM9gB98oF6t2uI/tgriZRu95JWJQ9GiKzV3HI1nUT8U5oNuiLcZE6
LXzZKusxR5N5qwQJLUlP5MrA9/79yWcBMdjgYkARGxaaHlVeEclhEB+m/dADoXK7gZCIRMTt6PKG
sdpA9SE9MB45IvzS4HUlhXxjQ4JT6O8XzvTS10OMu+FNPMExj0qDsRuYa1EVyF1J2exyDdpbY1x0
7RCb/kqfL0YNqH9oHQYtf4fw1ZKMTiwtQCMP9aSwz7npqerCPqQvVPPnadAgvPCwoXVKNSyAeJa9
ev4rlD7H1MET498voYewpRnVp4IWTZoayLkErm0qUFy8LglLRYNeEhoyPzvRo1Bc3Z+A/q00S1o1
E2JrLLkmAnECKAeX57sdH99gu/94NVl2qS1tgnUvepNhv3JoekrhxHHl5YfOQxkYAjwQW5po591k
9fECBqAkx16VrdEeZdWONGqhPvpd14K9crgfN86PHJu4E4oP3DQ7ws2PQSIaQaSk8hw7m3nRm23L
eYy17Njt7SEMxsVyRQWcyFFMSpMK8Ao2Y7VQB9wNL2JOikrX85jjMai8VaLZnK7A+FVWv/BWqm1U
Rxosza5iCrclN0fvemeLeKnhH1c9rmvRZhaY8MF6GiYZywH38cttX6JnPa1xGNH7euZsfslLZlqK
GuCYxLGrbm3SOiAIpPWZoAnuqO6h1wkqqHT59pE4KGusXNHIDoPJhAgEc1ncspIufBX1adKIREFj
2SEVCVft99vv86T628GzrUojcsq/+egOE17H6I/NZpx29FyJMWZ+010lUBr5fzUXvDnXKrAvH4D6
FcFDpYuAdCinFCWFpy3pBbJr8r4DLRVn2BCpCdah7IajkSoyx8ST6sbLvkcU34hgSc4OUzYlHkhA
7S91FhHDEF6IEA1qIPP/cXc+wiJ4ftxXU7UvxhpbSMCWL5+AVx/YModgjlmXQY6c0P+3Gv12NuE+
VNWwstCaZRZDOBxH80zabzRT1Hsx4Mr0qBOnNNUk3uw38NBNFLH04m7WESAOr25fdb52mHaBmoqu
wzShp46fo2CtM1bZfjvsP9HAOSpWD0WyBOl4Wis17gp+5rJxpdnH2a1QUPRWou1i7tjQGhF3IKcC
3lnN0YSmsC5iDDW/xL9BxTJyYZ6ewRO/+mBU1wq7QINF9c2H1S6syifhjdsEfx+2VAcxYY8qiuiJ
eDOHGuD7ZlysyNcZRNNPAryCo3UI6nNSG/ohX6xsVraLf6mhPanUqg544P73MLQQnFDE1ahGiM3s
Rc3S9Rx1t6LRO8lUG9o4Bxa1TIPhqJeFpOjcfFQ0ZE+woBI11nmca4WX2K1L9sE7e3yH+qNAWqZa
+nwTgQYocSCVflbvHzy+pU8LD0MqXb3PS+6W4e/pWipC4uNFd3K9NDeQXsyFu6BY0yQXCVYMH56z
hBTDk8BxENtAp+L67khCHiAbbSzZdr4YhXmBWQiDdxh7XNQthwsuGprwdVabmJ/Ke6O/YFZ8ZnNt
4mgesHQLPTr/CStoxBCGGfQecHCGe+iiWv8amYlcpEmO0+VCBovdzHT50Yemmal11f6PQfuvb1VF
K6WlBPXR3J9PW2TFShLwsAbpPv30LzvOXjGAjXdscO6k1VlEkemmgr2FuQWi8fiEvwMQuSCAtbBr
L1LpenI92cqFN4KOdKA3cevUSyLROTsALT68eeiFDPJl5nRjmuzSp47mn/OVfJUmbQdVHbmPlhq0
X2Q9bFDEnQiVhz0rgoYn7t7bFdD2kvW1aPAz3lwLSY2w939frgIJO/ZzOQj8yjjnaIPpLgOzvQSv
bkaA9jjCOKlLXDNeGgCW4Lns3LlfHuez5HONen0c2V8ewi80fhfjzqZKC5tDNK8RcHSc2WvXZMV9
2uOWpXhgIy1dOS2DwsZ0OoK4BuQn9B7hMoe3myGcnWiLGDIxjvkYEBQ4hvpHfyF5kJdHmmWngZb3
epTKl8SChZzcktYoAGqdl4b9yPpW//iwE+KEreodC7s5myE9cPl8iSRE7k5MdjZB7xU2FQUA8i+q
i+DMyq1lO6yNBzBTm/A4fJE/f++dMEMVg2xoMOHQ6c+32ubw4D/tCfSTfkkUVRLpbR7eWp2ySbjQ
jIQqovoYKRwBjXffwyxtHQMQnL+R3gfcpKPGfIGuB4GMEOINF4GJJWSP3LSiPWg14f9KFz+z0npY
IAx5J2QXV9DtZQD0a/Hm74nDyRpuhpFKxEWlKOuNLgeMZ/ual1l9Q8xUN4UNGNWcXbqxDzXPr7Bt
7ubzNRwPOVlOVNHQkzm6NcEFgHeAqcipnfMwOtzAAKCbBbR0Re0RKjH2kq418pich9P3Teum+z8A
El4unTjTtIsPoWPCToB7Q6mFkmBz3uObKxbQjK8LnRATx3yHKsyhfdXfHQrmbHRdr8KlxHSN0kqa
jAiHN9kOGfjfpp+igeIOv02QC8YM7hEBVpItKmGgMpQO4JiO2EmFEPugifUr+GaT3jnTCBASbAmq
ROnN7jsHT00HO4n2SnDTqAO9CYFYZ7jyA3wqznnQGe10KKBuaEMUyC8tijHeqeYdzKPoGNAT2zBY
Ou2xv6gy+OsRuW6loijGI6Umds4nbRlUb3C4B6O1U0aeb64dOUh479IqJue9JV3q5Pfc5VYVAZsk
NddK3miCOAYBcLE5bYVOM20XREO+/IYXUwIInVanckO+TB2BbTsRbCau1M+kxEez7+kRXqBnBKH6
DcICcaWRkaLA33+lNu2SzOi8rc+Fxmh3JHmR7pOu8qw62r0W9sdwh5LQVQOb0+ZzdfreF8BQNFoH
6N5DOEed/H4DHRlAvcEsjGy7TwM1KLbwgAuVkFqGlzVXQdq69f69gxPHVQgoXIJzc08H/AgQvxK+
2PnWb/OzMJ4YgqFB5xv8kZTpVwa09AYJLLkXwxegeobUCUcNsHmBkGxP1d8MeWXpHdbLFTl3Er6D
LHMwz4DNV0UZbjGkNN7tncW7hpYRdP+W8qoTrQe1G8Pr2M/rblPlU8ex5yCwfxKT5yRAj9sPIZv+
8Hdbe27Y6qYUOMiTzGPWAh1ITq8YAgDe9KQnli91MMxlcjAoFN5p2mRrvZnQ3IWBPhha+erxN+fn
bhzy/oPykhAqN3SYZ6sniBeGfLfgtnM7brPAgTB//cuk/G4se8MFrwtqGPH2ozpU6JbZeecVftmI
mpnjADizLF9d2b7ws5iqGxJPrOJJzXGyVZZYmyAf2RUpnUxptGQ0xfsfyKDA1mgUqB8KK7LkvFQa
DWAUkYhHUVTtxDlyAYna6wgfroyxJsjuSbVsLG4L19n0FrF3nIHahmk9BnvTxsc9uuQICHsWSW4R
s6GhTNZ6C5/AJ2bL9wkeIyiZT6UEgoKXxGpsmjb912Tvreh1L6TcKTJRdN4l71UhM76fG5cmyASA
2uKGRRDDd1oAsDl9pVcd+uCKBvGsNAr4crY7Mx8gFu5ILoaUgAdayfJ2wuJ7R/wwmLFz6rhIlWuc
ZadkzCkWFYvEMJyDIVC8H4kYFndNKK33xdaPNHv7ZlUKvdc4R76EPUXQQrJdyuIT8kCp494rvk5g
VlqEG3+OwmUPAZGPXowE3ilFlr8Al21caqdaBhtmegWHp9TigwWBpoo992Y8ZDuQZpRr7FE2oIsj
fVDI5cT1zLhWjhnO97AqPwaYk3E9zV5BfeCsMsXSTqM32Whd9eh8X3l+4xCrwMyFgzQBOO/Ko3QM
BiChJ2HYuBfh50xKkVKq+ghYzZOhEedcqzPmze58ES1G3/IDe3AO7s2QhEXOGAgbBfTQKV4G9Qmh
iSWbV9f6jjeUpEaAIYxJWMBownZGKTaJ9lYbv7WItlpKqzpLSnuG4p/QNCissxdkb13K28Z4cSfD
wOKrjCixXwIRJsliIJ3TsEEPl3WXf4M6wLhDF4jUoQTeuZbmHgLgMpYWcRcTAmobqS4YUL0an5I0
1NVlWkMcwH8TkaIFCNxcippfHNP0xYToMiNExJ/P3IioO4g1LldoUmJ5w56hvhlS0Jg03u7qjYqx
o0V19RsVsHy5QtLdZxUb7QT9Jz4A+ByEYdBE9uQ/A5Wnhb1JOtSZa/Vk18Xkv3ssEIW3LgMVrsm0
H/08sRIsxY5yy+QRLMZeATFTagPkVqAjThcXjXTx7LSdH3sbEYUyGSUqWH36KCOjuFB2Xe5b2ba1
ZE5Zghczc0R7QJd/ZqpPhAz2lTvklWCXOxJUgf3uKP5QU4YYTRVqibZzkyK2e/R6d8PrclF04Bsx
vbBQpihM025Wf3ACJ+Mw565SmopLxdShJ2o3RbGTCQdTphEpE/F6h79uqUGMolqvzJbGHbP9oDKr
GEz93lOHm7l4d5mD/czbF4yKUakGKLm0psowqzxbRzpa3wAl+zPPYm9ccHTB05T1VzfOCxwAHzT4
hRrg/3D3sYDm++0Vus2lCmeWueOxvNt49j2kdO2OlRcj+tjZ5ZtITifxRZku2Q37F3lgV8y++vk5
vn3tyWusPj9leMckT9DP2T5QBuvQmBCDyZqvhBXp6P1DuABKGPVTfm3e3m7iEggk3hHeqt+rPRCW
0kaqLpKxkNdFF4+JTrT1+gU5xA2pbtJ+Aw45RKV+eVXlTW7P0mJ9088aJCodp3Q58zetjqlqrZed
O1f7yvqD+oejsRAoE8IykB9qIQ8fyvnjRRv8D5qPRRdqsx7c8jJS0S2s2lRo9hJ2mQfttdtjNGAN
T4BCxJ8ZNaybMdTdAClBpz3mhdPnqBNM/Z1SFyoj5jVzJqbdxVT1awasLaLESO8+u1T/mvjdSCo6
PuKsl3q5Fmh9jcXL99FCBsXrzpfKDLghoPvQKgByKTVO7qWKjLxvZbZhlZQFfy3AGHmBHtXiEyfV
evFqRqSvQ062owUx/V60Q/77nbkXmknsvPIuBTcueFRXYPQzh6c0lT+sSMFbUnM/6QHd2mz57IS9
pUsHEtRirrQ2KpHlzUzgOGuNlDPvUPrZAgJ6sZ6fm/IDmlQnmiKwrDiTbK04Ps6cwcIwYdsjGsXl
Y8We2stsSXPB2eEyo0XBJPF31uuNiCI5yRO8WJh8PzChGytPh1SygRpAHz6SwhXfRxoy5vqB8d4r
nnTzsFQs9Ggze+6VKoduAPtJekKSDF2OukRQ5TwfN0zbonfM2pnUMrjoYNLQpYRZKtwU25U8lCjf
6M5r4NNRlk/h1eGVZt00FldEIAZbkaUQPVHbuZd7ZV7hz9ChMitTTUu2Pv8MXjaiQMpqj74etW95
2Xq3jr9XufHcELuKNGguu1Me6pIdiywv8inkcZXxWJrT0SNZaPk2JhtwTIdHjBQwnKPcGonMh2GY
cPyLTUvE/1fPcQ+89J3xrjmrctN5EIgo0P5SEBMDEZ/X+4LiGbRS60WEN1K90HBDVfAOxB10O8Wj
DEw5VkmRvRfImcZ5/azNOdKQICJddKS08xcvlP5U/4J+OP4bGewd8wD+7n/QPR2nCPafieVGTkPJ
GtCMXvO1u169ALWYTPEIARq1Sfn/YvbujSoE9rnXUHaGkEjyrPNhLS+WuIPbXAk84kHP1tr9aqH3
d3GlP9u5DQVBqUQyGGHsiscSdSXyktdG5uGmTGH3JMj6xxABtDJSuuCm+Hzbjfp81oygLLiIxLFR
H2QXNI0ayhOfbtqZHiv+aGxNpdzzDBypzdej9ZxmsvUHUBRwWSkWUEvXPErDG4LgU0yMtKq9I/fd
BMS5iphif+YlzodKxwJFF5uqNdQAItLOUV6EknrVR7WA7b9HBxpHU011C4cqqFj6i92IAtAuoKB9
5a7R2JI2nWeTdLXgAY/5bheUcAATYU/QXbtKjENimvf0JVov3Kwr2DTimreZi44s4dlGdHfW+Yz7
4HIS6EBsvtvHUuNV6DWcXk1QSX5IOiMfCi7mUgx0x71Ew/TUphtEN0N6k6G/0t4jm240l9o/BeMs
J5+9EePLvt+miKm1UYXlugCEqxWob4FVcmXcmTdLXp9W2HDRw6oej6ygPwkUJtD2BT0lgTMd8JJo
PCnHesCrI7bm4xXQmRL7gLOr3W7AiOGzxqZ/lzPVPHYRLrEA1UOE9ekq62VwhW+bZoUGjoR+myi9
jmuMQD4uZ63GjpmPuJhxxH3ubE0RfmqaO8uqXewvL5KCM/hBAn/Yu0mcQwaFckvJjvx/xZEwzHAn
2O2zrwHxRWYRJNbbkrbW6tn/laMwMa98qxucb+0hQB+5+FbB5VIa8rRk9fId9BXIRL9qtkDZmY5M
JZcoRgn+JGbF3WE93uBqkV2RqODnZfLCdM9d6BNW+IfA9u6IXoCO1baY6ewBg+G6GsrQu7afsw+5
+ik1TviSsL6V7YnuNzE1wSVY0ZJNpsrF8Koxaq/Vfd3Avy65nK6gxb5FAQfoKvKDFHQQ2oy17nGQ
Hzo8awDiPpq8dF7SUFLxoj4u9JJk+gleMaLs2vckIIoFwwm3ojpY7uYEYTq0nnFh1HywrqS5Gzq/
umdwRHuX3Oj6+fFqoIOMhpOEt3rgh4F6W8HinLgemdbPEib+FZwqaqwtm2gpVqwlB4FWZ7hOodDN
AYgEUKgi28E+GQlG8pj10hfU0BdyC6ilB9afLWNOCPtWvxV/I/vO4CFZKjbTsUC50Bow2ootN0dH
8uHHVr7x9NJ/kywqNEu8pzjhrfUaJxcz0XpLGC5upIV4rOYW8pleanLoEhGLVQhCYkMEOLugxyzn
HWoUsn7AJvA0AjgeLBXHs/kpKpmjGwKqaIZFHGGConbhZ0fMf0iwiHNESrTzudkY266763rZV8l/
4vcUaFjg0ryuhkR6urWw13qGhyYX17Fmth4aIv41tCX/U0X0VEea5CAUqgMTiUt8lqVNSGX2he5S
8Ze5C7u1/4X5AEAHz5vx9aBJWFVNg/wzJkm/xeNJsEvRrpniZJEZxodUdNVSIth1o60ZXuAHj3Ld
zE5y9jMnkvLEEXjII0lv0VCqRGPBngpNQDIlmHcZKN/5F1Fc4pegw8xdkGccpKTqlYV3oiK9EE2l
7U/Wnyo8kmW9BnV9ptah+cwPKazJ6NZ9QZ5ogksN3UkVcbuEeQ9WB10QHQrhmBEj8pm1SDMNTY/y
XPwnudbge2pnbgNgbEdzmjFHRDRhXl5HIevJCnMSZL1A9llttbWoSKOKcmyZstm4P1u4wCJNqOyt
PUVkF7KQwi5XJhKkJJ01M5IHzQDiJ6IPyXhPazwSv69ZoRf2ke8/mZeOKdBSpLun/vDvU0g79hD6
dwc0NtpkB2/0Hogd+tIEGJnwi+jH5dFinRpV0GCfz31wOR70cxqlakaCYxQjm+CNMt7gN/7vBtCX
cMdZizRj99ZMqxtzS036OwMfIaSYUqG/oVsnTe5635wJdfUSAQmFNZzpIihMFuG+PgPe724sLbbk
Zvhg53wZC1lXlizwm12tBj6GxJ96t9DICushP3JlN7vCf5wjUbFiJLyLDAeCQY1qya04qVUA4eVA
C0tE6oqnAZvMFKfG9gc4ftHgwUFZkWatf9cC496utDxW6Ejc7aLvmccii6t23QRdGeXzqPERAuFS
Scq0LGL2mEJLthWicvrWI8RVgyyfc7CdOjxinixbjLYotKbC+jqSb91n4wBTlelt7ckUFENM9CbF
0RNm67IPj4WL2Atzv0K/zvyjwzbzVKwIsfO/76eopQgUINVZMakEA1+sh/bof1LvYuef+d7O+9vy
1Hg/ZsXWAM5DYm4/Tz0wmmc3N0I2WzkZ5cQARsvLFyKwc9shFGpnZAkFRJ1syUTdTedrooODZFZ3
2e4gb8HWLmAUbLQdCwglTPZImw40sWFjdMKYnZOvLPoI8g+U8zZ4tfhpGK/cwvqpAuC+muYertA5
ydr145vLeM5qf6SIH5PEn7GmAjulhEs9XNp48L/tL+zDKq6dlsJ0jpI58lLZU8m40soEzh/XZ2gN
12KFYtAusmFOnXNoZIfQrXmWiDzzYaie/aNjhNM6V9MN3CHXGri1/pUELzBbjKMBvlMSFQ4g2lPt
tk2HUBf4+pSWKm8hmt69sSlkN2Yd4wfbI/bnzzjeUhFZEP8nJk8YMtxuOV4AMKtGGHyjcAjf+LNR
bMWx0qBMtrboNwiInCMnorub+Jq0NK3q3yYfjBxhjkwgs7Jbnp9dLRIWC8oTchBCrcWwy3ezfSlT
lFOhMFHhQnJ4CsBXNcNaJucT+o8MetHLzYWJ3Z5rZxKaGExSdTttDvw3+1NyJCjm+igQn/XIJqyS
UqvAPg8aQkhdzZZsAflF/RBWQIP6Xk6acwiWpZ3HXL3oF2NuU6rnM2qJ3aWPe7m903PJA3IS+cjN
HbwIQbh1NnJDSGbf0aama6tP7zzFxsRIaPtBxKeuesAIMCfYVICDrDYpT9/7HDb+ZguD9r+wL64r
RDoY0ZSWpggrI/QN6lLIjqM07tyDHO6XVhUHfj2Drf7Eg7Zig2TWHPW+3AA8iQzFBdWc0GW+1wVt
sjrw0V28bhKWnnDkPuysBzhfNGhJCXslcsAAiQdmAbxFezRb5uZ28ljOJtolUQjNQ0hDfZqvT2Rw
gzSiWf4HtmMNVjeB/La+lgGx3ai8g+PIenLIjT8bWqDbKMlDhmO2ATxQt7uk1m5VigLjqLKCZkZ8
eki5UcrAaJULp/XEdgiegbaAYRTitN1AReU/MfAXm+BERK41qIRcZDLz3mMcNbUSPDKbft+i02+/
bYXI6kvIyeUFHtpR7DQUyDEx8QVD2S7QApXvGyJNqmFTDpXo1Pq5iaC7EVyHoZLzkmTgSP+quoF7
nIPX4UckPZfzk+XbDlx1IZW2VqEifQ5ElcnupwFpZCaEK10jPG//H/rdPWYSVDIJUnmzaI4EGKo1
OVUSr0nd66loKeCqnS3ipSCOTyCqdUUDf7h9rVsczXeJi/mnw1cZgN0all5Q54zfmYEbzVB8IJw1
/IrWWNVZUJoagVysf2RCBlcwzmSqVbcng8maz5/F8dUAnE7mI66SVVQtjUPpgZN+bDPzUl5L/JKb
O49ro5FVex3FErjhU2DWIR3mHhpOGFyip/2lbbtJa/rEKTbsh4wlRh22reVDCNS4cnhmBQc0raYR
QJ/ZAFago3k8KDKMaECoxJnYomO9AQ7vzoIc/0XsxL5nbUJWYM1u24tDyG3um+cHBM5Qp4dbN0ka
nsZOWJRWjk05une68tkcw+jYb00zbtvgpaO8cFUxysEmfHi9+vnnoROizheYnMgurGALL6xWeD2/
Q6aWsAjjYpM9jQsRSVAu9Nw/+F+JpdwbgiZ6ptU1VegPLJ0hTa9OL0nmbjiNFFw8jzDUCb1MYtWG
QXoLBQPxcC29xC3gq8XJDNpxDkUy9yrtKcl8enHvwqEayBY816K4WwV8L3GK1lu6YTkNzP7Tilfj
kw4ugN0kJJeO0C9BQazjZdBrRk79aQ/nGGBnRRLBFZsZqADIBg9ji8ONOEV9ZSXgYKK6H4o5JpRK
7uLsevz7ijSv4t9jJ8l6HBgGsTnrj1Ww6gOs7VUEisaRqhdFzSQHxNKMNjZfHyQcW54wI/6ADRUL
ZishMq/3l4s40ztiE1OQYY1PFDFjz96w6H5njA77ncFTnxCtuJxk+f36YWrpuMdo67thY6v2EEzw
aafEkXwYoCptOV7PBMhbAx3ROkIJjHs7l360E+X9PT5q1ebDsCdzb1HHYDIXS6SnNxo1lheb4XKY
RTXSJ/g/69myiZFeytU9n8s1J0mmaljZvNG8HR3IWsb37htzu77UMx6jDwhgdEN5ThjJOGlSu8VQ
EQkdf+kuA2fGAtSogkHIBoGDyWu6h3T3pZF1wOxDGgsuMypDUZwUXlgYMvkVgXyS1msejVc2llbj
2Xit2eHCdJ4j3FFy6HZFoc8CoTzzAUj0TYKWYbneVow9VNfbUP7Pqw6clqWW/fLR9c/+OoVwK+G3
MJgLrHkAR8QsnxJiiEC5SZMmgsTuvNr86s/1kbG1G3NrVAIJNUSgIjpBv84HaABK2Jj7RBVhuSy4
Pfe4C5xF2+s/T2WIHvwBBXtAx0qI8HJUW9wZcMr5XAaCG1ZvMFOEv48B6ERSECCfNMqZCJDzIi4G
nwny7ojdZRFOOWnx6eTPMJF4ZG5+JEoMMi60aZtGIKe3E8eMvxdC4dcaTF4FnhMnjx2abz2xtdrn
ZkXXaSERT864Q2QvRHcbNxhdnW1tFAaEuQpdmbrrQcbfTv66OuDBrMlZU4XnRn/KFTTzlskOrG7n
WdC92w2BsOqwtVD4r2zkxUBcq9L/J2A1+BwRzDsKnEtNaoTkVBpidM5r1bUpx0qtfV/f8XdeF9YN
gQGTaI5w7Rd5VR58CsilWtoNqvUYQuKHzQdHuQQchhsCNcrZkfp8QBxdJDnTDDPmAq1if9K+Ydet
X1vTrl4CGaN/YpyDZdm2hTe4+CArZOq21wwYMBQvcuNMneE4qLUHAV3BQdNEoqKbONBfENNr4wNK
dkuEyikkW320LAUvSzmKm3GI3BH8lGjqz+ISpjqk9g0su6PhHVd9Vuj0GGwqVfCceEilSbWZ1n1M
PqK/Gn5W4C2GoVqCC57psCdQN9/I4RVx5T3tvlYscCH8nD70MXD8G6t9mDn7HB1FWEahPhgqezje
Uxk1qOP7HDAgE355K3AZNTLvRZoprpDxcn6kzRVW9Yp7Y/fVrBYEehNqLZLjhT/uWi5dV+/Qz6R/
FuD1Gw4KXgc8XKIiadXtl7l8rsvSZHyPF2SaClVJmMy+5bQyc007hUfLlbOsn2k+zcrX9n0TigsQ
Zx6htktjRk2FDlTPJoq4vDVK9sQgmM/ta8IVGF/o+L2IMxk9HNrSYNo8on3eycwJhsF7IK0jYziq
Hl3ht4a2R034SsR+NiGxm3nYVL69YxA/7gHix++W7W7k3rPrga4JbkKLpbEgX/6R2WFsZVxqpOIC
bkf+MuOp8eLBLODeSBte+l8XLgWURrCmTD5LQpcG/8tYo1XsTZ4OJ4dwTxxQ0M7MGIaFLFKmux07
S6UmUwK+LmLH5b63tvzbfFQKwl6Vq89N6osWF8QhbOftxzQOU6foa7Os3UKFhLzmlxsHAPIsdzyC
kKk8uyKrIt04LdalaMBNKfEMZMBPp2r0wjTXYL30HxKclqlqOk66wsZXTj6BwkGGAoPGhbBNyEwu
lf+i9OPFnme0qmsrpLvS3KqScoRR/hB4j0YGguUMauU5wtc15DWupvaRgSa+YHTAA4u2CbymT2mf
pF/UtwAR4CsYJFGErYFCmxEz3IMoyezVHvtO0n/Ftj7ZOurrdWQJJ8CgCwKMjlkn4bcX5oGeWuWj
l62iw1JTHKH3gzQAANR4rehr+hDx6CB/4ouaNAFTrpxDbauz4BRuVnu5JodXGMm6LkE4KY0LXwh9
U/WF2e/S9/kAOPeEYqHfSSA95dsyVANkC1FWhMfpcjBLSszcr86U5zNRpI8L4yK912IyQrpoN/kc
UeDV+Aun97AlmTxARV7M9z7ABQk8OujGf3+5WqqgyzaZrJ5uzFM09mHYG0t0GuWHR1MTNtI5WLyW
PA6IqkIJMT0qS6jjnGsSLW2SFWYJgeq4+Qi8Lonv9+sKOde62jqwHc+v4eupI/5vKSWuNZAqIG4N
5YjbvsOUKe3NPDQtHRVIFICuEqtUbpUNRhzkN8z4oxJDk6k8LKJpg/EwPtIPz2D5AtVf4tEhtUjY
UnoynNky3aBPb+ZTVlEX9QEvjcBPH276ufOkeLKDz8ePAlj3UomkdLP7zHdpLNHF3l8TljDNuS4K
dRPON3EXnYswUFuGTOLyjtPSSZhvk+ZE+D6XDakhJUabsxVFfHxUcja6tizNCJG5Aa6Nmo8ODOyp
cd+co40mhR0BmUisEub5Mq8sZJXEsDgH3WqXK4xXpzuwNv2qyrzs56T21O+oUYlS8pAoRLiSZl1a
kpH9XXiH9p0RxN1bg0LvHdoU5HdTPj/VdbZdpogX8ipVq487z/aJ3FGA3HrX+kEjprfpKmVJiHZv
OJM0ylX9bgKUSp0abdlPAOt8RbmZnU8AM2xWhq0iqZ7pAoC8qMs88b33pbAuQsIVJnIZk/1EDmpV
wlhciSB8RD7ZNycKpuNChlFLTAM7i6YVp8su3LQncexPNztytDfp2XIkYP0WtNBmyg4zRTD+gkEc
pGIiqzc9D0cS8xVJmeVYATuhaX4cq87POeFgahUItsWBD8iauRbhFAhyRzkt+BPIVTIKy/0uAZHe
cs8g9ODGtT+3e/son6d1TBL/R7hjYf+9GG2qq5oA+UDhf+cNlmHQyKVMsu94d59819NAwL8PDKoO
657IS+lHv5HfqVIWNTNP7VOuF01xxP3Us+l5oORoAq+mST7seJRM230PznP2+PZqRxau3uBKcYsm
dDOD+0MuY/X6p2SkUJX4QRi73IiIc7lLCMFKYw0nPNPgaVKyl4hcAJSFOoXYFmcu0k271HNTXH51
BxQcnrKEZzujRX+cYWQVQrEtXtDgCm1tbhnxTykwD9jq82eqBAN/Tj4iz5K6RRQTE8Tmdzvmy1cg
FhIIUa+b55B3Lq9GV5fwjc+gsQIQAPiUeIX9C6R+DQ33YaP+dpR0lvtZ9KYYvYN1yJu11I6qROb8
8zXItAz7beglQABd8nLwnRxr55T5p2zS98WL1wiFKY3Pn++sF+ASuekY560Om0PqII1CDmlEEpaM
gCnWIeJPvvg/qx/GFlQcIwwCCsrHKek2vcCvkWCQX+mjKNb5TQTtn6njB49f7W4dQU5YNkwiK2BA
EFsueZ6gcuLOH+3cyC5q439y+a4fwEeC2y7ZoLFJ/S16SyrIAQpnHWhP4sQudXu0FeteedgApvUQ
5bYAOgmiIbxBdmjrSBOdZH+IGGCKLaGWJBoKfyCuUCMuiGB7i7MxPtJ8mMb8p8pujWMyGIhyJDH7
1tXFeL7Hw9VBuStvEqETlls6CGltQ78nq2vZ3ccB8GMQoEM19k3I2+xgb0FtGuQeIX5R8hTbPwGz
4weeE74AhLqWlV5RhOdeOFkoezq6Y9LBokv/UMEe+nbxYpy5wDNsR+S2cVHuIxTAtPzqmET5tswZ
3B8mEJ80a8kAzVzcvGkYMb3ZwHchWoK1deiedPHBwpHfx8Q91CcDh3R25hGe0bHeWC3WLAEzvTDR
4+jXfG49mPeGB3vXLjLchiPd1XEbfm2xrF4ehIEHWNw0xjS5g6K8GmykaukAWtAi5UHsZ0T22Hhq
sh9L3ATTWafK1Hzk94a+hrhleeMLGbL0e3K0RT2F1QF3Yafds87v07XvV3HREcp9boZn6Fer1o6w
bkaj81YwN1/YNl3tCaFMM6UaIwxexEax1H4pdT7AF7KAewa3AKYrclvwymuao9rEbfE9Qq3DQDSK
Vkl9vOEStF3kASYT53BU12QYJKitMpgM1VGM9yByJK7dyrYCij8c4JbCVT8qqEyahcoDDvn3vMeC
yt2vJZpJq9JbtSlmHkW7OGT7WDoQ6mwcc5fznVY1KEB38+RcHytVXe4IrLYIVEHqZLlcqE85hOy6
W6tm6kN7fEsFfymrfqLfqlLvBYSJ0lTTZ4bVges58MGzNo2sXmYxBSJWe9v8VW721xwf5woGVujq
e+5xtWje2/qixnhg3bZRRDWU6TNDRR+2UyO13BXRRRMZQMsYUUJidF75kjVyAzhF0vnYpmCt2eJe
2xLT8wmQHggPfp3vV39Mqg6f5W9k35yyjbYoPfPwhnf7zV6CTLMs/vRqS/Gq7bcm50kKGvEd56yD
cbj94xAHWdF8wvZWYeeeLU1uJ4w7k+5as+3r6omwEWs4lhziH8tSvpppr7lPU9/XPlcjXdi+cDhC
v38ml7tR8jPgfcjSN+HJPLYHfsPKwnMRh1x8XBKUXVS/W03vWBJco1ta6SHn9v735bPq83qleZ8G
ccUabTQHBEqfuFlJYWcM+6iLTcLiWtBL6p7SwzZq0yquX2AiOyGFDNyvfgv+62ZK8as8H4uY4lsh
XERPvxoMOOIDQUDNS4+yOx0k6msHHwt/gEnAM4nQL2NwFdXlPUk8ajT+6g/ztUJLElu/7DHH/OJB
tFRwMIoDnIDHy1NV96xQmKrtxHFaxgkhkn/PaRanVcREhdGFLrtDj7980zSJPr7vCGTns3rZTRe/
TuvGmznWfWVj8vfSgXTPlzSo8VtMgCp8aESp8EvUSBgla2QLQWqEbjHvTIr80wZ0k0mqKNz98LUK
McFUIvWzdLBIip77UQOzW6u4JtRRDj46EeCz2cZhUycww31CdQuUq2uTyEILCUa6vl9ZKFspDQUU
qJMEI+WleMtL7t9iBTd14mwb1dRmc73914B5n5CUQMkbxYQSR8xAUGhB3EJ/WlpdF0VkB4ryb4I4
kZA1VCZoz9xZDTkgX278DQLjpm/Ne0Di6tkP0JMCYLpJgBYzCviDk3aeiVYdQ4+oEXTHSlopZpIM
jnYytejgocjdfjw15IYN68QedrlvR5fN9S5nz+i+taXg5Wp1Qhmsnf+MahVLiDKOuDgNAQS4SAtJ
Wc15833uetUNE+fX/f+LcndtlNmYPMrA9YevOZhQcgJmrL/wWq7+1S4wT+coacoUcWdEtbbbiUip
TYgRbgxiAM7rTEGqQCeMPivYItV8JFCws5IVLTOgeFmIkJt5n+xP0AD/MsJJ4JM+V9j8U0w/PJcf
koH2AKEcXQANHPYqVEiFIOa6ZedKS6kqUHDyjjPg9Z5ZHr2euk0IvFQ9Zs2Qy6qXnVs0jacxTE5p
IcQK3r4/nssjopNrD5dc/VXqLCOFzRcM6+sQXaULrsRBWl6cgSax+evkkjSm0SiUSBAAl3P4QSM5
m4Ao1kizuPzeo1RPMtSgdRYnPQ2ZxPnXTRfgg8//Ut9MJJgywcHOEmw3XPd/gKW2ARABBFC6Zh3a
Py7NMfLD5yuL9zAo4KBy4dndmWOR1Ht8FQsIJDeR8VTYdkzr/DMp87ayX7HXX2Lbc6YRj67Xil8r
oByHyRgSkMeq1M18NVmCMxAglVT7dpPueO13pxGTxGBjwQiiw+j1Se5ASNxw8OLM1GCoh2ismuP5
dA3VayXCUu7KswhxPDEFpicvgDicdi7OiH6c4RnPAoU6l4J5jApSi+kTCF8EM3rYXt234oOErhMO
70YOkCpfEyKYI/KI+TmJWzJQ2qSzrAlQtzEKs2inEBiafHdnwH4Hi9mTKj4P4D9ReF906f3ds4gB
UR0Meth/3ovZD/9d+38N+PN8CM2wU8N14NtnXLQK3nO4lKFUHRdpKQXseAhT1xWyAXEZTwUxXCFv
x7+RtpfGIz1U3PmuIRWJkV9l8XSbvh7cnjgLO44uLxGrofc8jB2R0Ss+3tcFB2/rlMt0nSVuDlei
jbAB6LKkqzoU7FvSp6E6olK+sreFCz+QCfh9ykMM3piqBV0VeWlwG/D/T7tpQFvQnLCWPwUtbnYK
vsrdzVCXRLO2Fbqz/v2NxFOax+I7UlTOeNATqSmBCydSZ03+ZoN1vS6UNmsBdIbJgmeMxeuFvtHW
oJPC83ZgKWQNP2dEFJZ2HVgAl+00ZKyu2XQW/c2kV5o1oGPw7FcnFtRVBFIyACIKwy758PrhTs6Q
Mg6Yn3uCIkKrnehJyboGL+0sz30bc7IVyeedSv4myzD9+JIc2sWD0kBcmaU/TnuqYboVmg1It7MU
q6lFtvcukBldzJ+0YXNd5K/Uu75vZ1huF0ZLJzA2eIz5TMxwd3Tn5W2HkFq5NJBSpC+4W2t5xj+Y
zWDJ+ztPKjyH0MMp/gKUtW8orHkM2Nrye714iAd685k3TckT/fk5hGPsZAE79StmakJOMDMikSve
siTG0j/fXQtNbKdYFeSb6UXQjbCGC+V/E0WJu3MUdgRmHaToglVBDZWh6gur4YpkZ57uWQJJWh/6
t0YR9wjoUyaPpOd+MAgdUQ9BWgKd0Cnr5GPtHxu6/NhZs7T7N6fbcQNq0tqkWqnVOq5G0kWyb5lZ
qDlH8kuJS4VI2792D9Wijs0u4tHb26eTmX67djDjmBrFsmIqAqWLPiMT0sIw2uBsuM3Uw/6GkU0k
g9dVb8th/ePft8MEZ+gR/D1w1BKi8+KHH/usncjQi8RDiKgwUoC3m/eWSbAKi0jigFY6dvvg5WSD
/klCJu/l12A6i5G6xUNvICES/DBBuRqnuDoC3rJQ/Tm22NV69arXg//nMJ9giij06dvYjuJKXrfc
IT/8CU3+CBlAgxi0Y2FbHDke1poRVGCIieXvVeqEQQN+tZ+ePBTf1xX+h3+JZj1b1Ja48LO1kizN
dQWl5bjr/VBniOk9n3TaXKbidXk6pU2N6Q5Iy8OEj/D3ivDd/VyDDQbZEtn8nCbgaK4pZEklU/XP
WoHDYJwfhrK8fpbla2V7Cvf1nuZsYrcCMx2UjqUFrtsGRH8NbtWg7XlJsv1ByUdTbkSwx/9YMv0k
XP7D9IWl8gTL/VxaGS+/kIicKmGw1M74zHvagk6eB1Vu3+OR4h20o57s3HDV3Js9abGA9Qkv7EEK
OIroE8EbeUdGM44DV/LOnTu4v2eSUGYlc6jXXqfYrck0Q3Em4cAuorn8Yk297TNwwzdP+zdwI3Bm
IkG0AgGAkVyOYJeiwBoV131/XGfRYLcd20KaGeNSFelZGS7YDfpidi5cJmF86hJD8eQXoxGneClH
SyJ6Focp6IY+RjfV01qIV5NR6FeQ0D/6iwi8knTfifGUn4UOHeoFa4L03AVtsnHwuvIv/DZb5S78
UpLmkdoicdBBMzxaCIpYUmjoi9XF8X5EjulxHG8qzmUBnPOY+dgCQ12rChI9UkRVDRnHVzE15KGZ
kG2yOuhW1gCIBEHGli3tQSHj+kTlR84kqmMV1Iz6wekKIPftH/TesTzGzxEDpThpsil2Rg+H/2ND
F9mo6zyeDDzYg++5PbAzmifmCsgYHtqmj+ryelxc+Bm75kA9ad+uTnchZE7FmTAST/wWTtnydjXZ
aBwhgBgSaJqEfGsrFszs3AqM196tlsx9CAvwLR+yKYdU/MNW/JIvgHdFqcKLQzqYY3WbjmiPNwd8
29KMS7s88bPipjgU7Lt14Cl134rMDbYyqhVDXoL9cBxq18EFSq9rgur777dRZ3R8ror2iJwBtnpL
W2AYp+UTKBdnVOTBQ13wELef330w0yS/ds6VYSvx6pw/S3fVdH/NiDaSJNy1INHatw3GJ3GXlLi9
HZTuhlpZBxjzibwjmniPxcBZGbpGlCYYND3NvBU5JxJBruJnG29Tm7vyy14oj+9Jhf0uPtrZOC7c
s+wh1id+JVK0GY8lQMOOk27oErSH6SI5EdzOEi7fgOOkiNdUxXObcuNZ4QcxpQgUB7TCyDEX5eVs
flNaBV9ym9S8nuEAGlcUahr8qR7ZgGzGQGoploggRKoPBaqHi5iBj5GUbLuggNFmmWXK6lH/RVmF
NibGgxUq2b89OfwVRnjBM8ilTJtBe8IBcMWRK03UJ9VVNX51kWgrc/6UQ5tQtWSxa1UZQKew6NHG
tZ3IHn208TtU01oDx6pQJyy5WUN+bLd5Sd+nstyobO9UL063BoLgXCCNIt8bSfEQOxA9Y3PAJ1Pz
3VFQhPtYlFfeP4NJH0ruYbM2DEZxpq3vR0mvoaJjZwaJPwZ/lks5mVhGq5bQPIGjqAwqDvANfsex
CGnSr6QySTOH+wpo9jOfSEYT635kZoq5gUrq5JQJ+5H6A70QOfUp3N8YN1czznpJpcTa60ZafIQD
wPIKpursid92NFhTG/OfkJPvaMvqONepQ2LJRiOL4HgskyvaaweS79Fv46DGhC70qTdcEkrP7Xy+
0nZLPCNcQGBOC3/MNYaxK4pEUX8CeIAJlGZzbaZcRiSAfviQnCFkozKv/rpnaz+nuZcw6KQSg1T4
Yh5P/BfdopT3Ak+Gy6M9bV+VLgPWoi4h6ELRhxuyQH6Ue67eTECDI2pGZpHYlm7XWE+CSDtgV7vG
duh6LER9sAHlMLI/BB0DWz4S9mIFwyTcKbPAW8Ci28rdLxpbFfXzMmNxPJDcUrH0TVVYb/30Bmzd
0UaKeqkfEoHvHzpLJSyQl/yBJLcxT20YmziTNpK/fJ31LtUN4lWLLZaU99O9P0PCiyF132qdP5m5
gZDhwKTx/SrbkQU0bMChqfZxR37MYzTz8uo3Ng9Uw5crGJL6y4ACgOkaYREaC9hXrEKUDgjOTyO0
c82u0EIm0chN+S56QAbcinzay3fNRtC9QfRZTCwfDBXDl8K6mANzrBWwJfRHGgJAYgjkWt8AuLBi
elnkNYzMSFnebL4parqJ6JCAN2+M90j5ERbPLiveC1a0LdZT301gnePN2cnplakBf/yaE3E7Qujb
FkxwsUF2KQTuJnJZAGpGy712JeiUfpOMaJi1FWJ0FN2hCXQ6oRDpvc7cgm6eZLO3ihqZNFuaWud/
wI04TTAZ4Rp/0dPVroq/O1OWHJ4BcvOy50xVTIgKj6I217lzuFovgSAe+6oCYem6D9p8KbuLXGIm
x+ih6A7OPp/fAlz9Htq7Jji9zrpbuKNfNLde5nIfiecOm2TekN0rzktr0Zz59rd52JXqB/tfbKzd
G52T0bV603pZI3dAbBfJEMFjpMR0xwMq9SN0ZIVfjiOVll6f30CCB3VSX+fibKMXel3DxOFS+2Ot
LydjzKWo/YSkhpFOe9GvvKMNJPbSCYMr5CqbbIhz6qB376oCmK0Eqq0dV/zgwRCXpdM03sI5r4vu
zFsY9H9PbFFIiafd2vtdfj2WL75/0wWXkQ5sCciBKPBz/MlNV6mBxzODF/v6udb/iV8WoxRtBS/X
aoXFULkn8weyZJB1fnMkSKhCo1KpgYg8IIrxX9JLGfmH5xsx39LWL45uLLz1NjWW2Qr1ZEeFp0pD
Vd1ZXVLgI13TFzUdOdWkos2k1Eq+z2tLUTCjWhL9wrg2NyOuxvZJ3gmMK0W91izkO8DrSf0UDLml
qnNJY5IjwbDgNcU2uEvCyNAJlwaBJ8IU8xUqD25IaW+LUwmYHmBXhSvuySaE9nNzx+0bepYT73GJ
pJXqFodCxQJJr4wdKjdDmtfnPPet0SCYkBcBQOgwK8XCERqPJm/CSxaRotOmXNOlGdiJKtZHhpI9
+Ixbdq9GyK6Z1N8tAyv9fLSUK4BI3Z0Gjv+R1c3/mwvWKHkdAwGnqqTv45Qyq8yQu8dmwdXOOWyQ
MtRIUQyFO6ML9wpCV8VGq5zhBM6myioOY/5A7+r1PSogejsm6NKlqNgWMMWSbLenXmq1mkMAzH0p
C8a7mE/ilJnTsltBzQkUPjy9xB6ZdzdZd8e1OlVUXeIIn2n42opze0JamLX4kWeffZq3A1dkuCBn
MdMwVcqUpv5vkmlLK7tRjOVm8s0WYLGIdE8Sexj8EXVVUXJLnqxeTzntgVbetjIBxayLCDo2ohSj
Vk/dnK1Rk8sbn/KUmKvQbT9TfQ2z6NwMuZ9hEGW3Csa87XA4bI82EU6HYsfT4JXeqYfPE8zRPWzh
+TC7LelWgvcFjpN5O1hnWoVux0Lfc/hWquwAlBsMiwe/LgAPpnqifF3fT8BeBasUH0QPOnXYQQhK
dDn83a/4hwTrC0lysqykcBmasxrQZGMnlO+11S4XhvcQ3+p+0gtCYGyrd1VJtb7EDqXgDPhuC/Z7
1o5trJLBIVxUc+F7PwhaxLEV7GIuSNKyUBvnfrozG+h4NvhYmK1SF5HVlBKtOt2EVuIANrua2m1F
MRH09w9NYz6PRLFfBFpFTU2xkZ78D4pAKMUhdix3U4asyABuRNnEEJvpsN2Ew6i9DZfQ8CWEE4FS
eliMbavly7wwVlqxbpZyWiHeuFv9yOTQvjrFOsTkVsYohlUKkwDG9r0GQpnDaePjJYkV/O+6sVII
0RYmoz+3DcHCMbrLChkmrEtjLisADkatSxqhwLuWxbBAj8GSWwdRxaGvCK7nMM3ZiKQBhNDHavrt
jomy63rvpzJnOwm9gXmkWGZmf4U5+pS38s2TDjg3vq29tWw68MqelYswcTyfHDzc+FNwtxWbQn+f
YilAT+n0/0oAQ/UZon7Lv3zj8sCop0OxrlHf67ucPWFfdr5KJHeTYKwIx2nI/wPfC0P+F45IAVSR
ChnSN5G3B2oQ5V4lgbQoDpf9xZ7TYwG1EsF9Q9wH/gv2o+RD1hR49GWRMEE02cgkGjedKHhPkvzV
/Tu2bBqdKmgjNmlwCVXc9hI71V2lINhVhGtQXF0imU5s2H0XBKwVMg5UvSTkIBNIAlhQNQbPuNgb
QCKNl9Ki+okiB9OLlrUwacXSbZASMDtXcjqf217ldF1xRLl+wBx2cvrQepOzoZcLudxyN4HLVC8j
azXo5PdNwJD7vNumdKY4ntfPKcNbzmsttdeEHwo4tv9kgGW7SyfxQqvbuj88emONOHCLM2vXoS60
EMA/GjykmEBaDe8qpy+efrBNhRq0sovA7RzkEahjmj4KV832xDK8++9MVRGXolAjdi/9g7mKLOSf
7JTjOoVu3zwFUlwVKYJ0KWNZVufn3MJag84+Zlxr+S7S0cnfQ6JoWXfY569HAyOKGbTgVc8hfF9L
CQIR4G0d29nm5Ok3szl+fQapHGxPzhQLuE7h2wdvnyTaByevGnwYUMTU/x/9o5Iwk+M3hzj0cPlA
MejjFi0vi19/Z+/7G7ynmStMB86hQgg+GkAY5kdI6B+2sB13VlS+OQFctroUO/6k1WiXhTBx2zeP
JlzfRvX41FN9GYgLF3I0/zuTjYvwNWu0g9CKfICQvi58u3kHFl+PM5obrGVxxJWTvGDBrWtrOTUA
j4QnndUVvSCVsrOkWb3yJ1rnD2Y8lKn/Df+Pum2x5ck7qTF3e3BVQqJi1lBvsLIJhlgrIGmczzUK
Vps1YQ5ENXM5yzSd80m3SzDa+vPbHryA8J5MmpdJ8EpltIKtMZxbyvnqm+dMjlUrsGCCUg+Ovub+
vMw4442vUd/Xh3FTXWlSx0h1oLb54hFVGzR/PDo1nJm6IcvUCAHr88C076lGHlMDpGCRnVzxNZBy
QQKNMGr73lgGhkS97tgPKuCaUw+rv1QnljvOQKCl6+AY8q90RbSaDpgllx+OAgZk0bC2w4x1d8+G
gOdm0rkcRlk7gYRLBRmu4iZ7s6FEqeDUVl42JvBu6ScgtJ/bLeCVZczcVEeSSzIzRGdqDTW0AhTN
4mx8kDbD9/c4n5bbMLF1KBvRcKh8CYLjG5RDbY1uLBn0kqMibinwhcrfT2ddcVqi/d614bzEFOEV
QE5yUDwO3B6aRh5FAAcgD7xERHj9P/d1aPGL8e+TMedbSoenM2e6I2x85lyBoDbJDxruR/MTZWpz
/UoKNA++MSECtmW+iyDhPBke+SVgxONqOtmQVORqRm6hkt2Gj5TZRKL2iUk+4g39jplqDUVlzfbr
+37CFv4myi5Oj1wtlAlDLdg19GlJh7zU5vP9Pq8Slq8zDoDi2ve9cBOZvPHPXPDs75thWis8SkF9
w/B8GTqFcm+fRVrEAQ/Okoel4P+7cBUBxck8y6m/kS3P5SN39FMu4k6n7DI6rt5slmYJ8SqQ4C03
BRwuF/zkCChvypxMuOub6Ceo1c+I6DgMchSBNtWe4vYmpFoyJF4AXtXhwXGMXkDVlguyw8iifxVA
GU7FbWjlgaloqHHTV0QOfgWO/0ClHD3spGHWY6dhqkrfSvMYifLtdSMzDHw9MvdTKkMBIn8GGkWK
x5Uxz9Kr39J1wtEtYZ0w1FkKkdkWlM1zlKjD166tMt9aGOkHt/tyrBYMYQLMnOjFPJ1KjsvcNJn0
34oN6NqNmhHoS3oyy3R32kVVhRrKkASQXYvFFHYMBaOumcj4Rn76L3IJXTKKLwEHc/gIMjcCxKnz
hzyh2iTX3C3QRkyPsjqPwNPFNbJZKx6eZ+h81fMuutGdqNIfBRuDPP+DOKsc+T1BLKvFr6cTe7SP
PStL2clzGbpQa23Dyj4RCUJWw4flj03j9T3sgH0EgslKgbF+lWLyvy/e2uM1KxC+bQgFvkCfOKak
d4K3SNZBAOKIwuT66gm7hH5m4gGM3DP36txtw8fdh47X/pLLZJYMHO5H3hN/xTqXPUOgTJegPrCh
BhpkijJHYQRHEeazumxhJO1Z2vVpZy8dVRlqDuhrw5ogY0KORkEDnW1qswBWbb4Oa/Gna35DqmqZ
YRMcMTtqCwFQXePRcJ1ikWpdysPCFhb5VVKGG8jdb/ZkkPKn3iY5yQXgzZvqJdo4VmoiPeL+w0m3
pPzR1WTHQWEP2V5v1dbgTwVIH5mmNcXK9Ls5YoSSyS+nNSzgUBjIHazDYOb0fBdmpp8xK8rPj71H
8/U1JHRHNd5ongDEwLEr1bpQiUmfcV/xMjL+oLunABHAhvCgy0wPZByzUfKjWiv0KqH3Bf9pP69H
4lqzRhPsaKSb9Fl5z/SriqXO/cNI7uQXNvxW76KDwqURiMQjt6zpv3CKXJWsCodtXimexDssktZi
D5HXIINR7/hethVljXUnYAqLDFITj2TpRUy3JBm179wpLt9l6xNZcTW/ZxeLm3WYtf5V9+p00omS
sv9W7N59AQrKS3vEBWq3mAuasllxYUWjG2N1RwySHQ0abC0AJn2cEVFT4SesPenv6eTYjdQOaon+
8oflwoyQHCPZJtFPZKnoOX9krBoUuQX/gN3GIUB+tSz7AS1CJmCyvIqiXAV+bCXjH3Rryiw+iaQH
eCOym6ySpj01Myxow6Oi+3QlM59aPtmiTgCYsqEn1g5bX+f2ii4DN4Pxvg7ixgpw8udjUaeDNlm0
mdW2B0MUKHL5rNny7Ke19aJI21Pej1zNrp6UnMrPd/+jTinV818a+ENVkpBms3HdMgOoSNoYgGch
gL/hXqv7cxJX3KSdy9kmixeHewjjICEpDpKCRaVDWKNql9rzTsdbUbIyCVtJtlp5NAx5/O9yBMGM
DCoz2pCfGxgtRV1y0DK9rQ8/2MjD72RX+nB76YnaTacw7zmbaw4H2NSI79qEhc9BnC8OcV4QYwnk
KRg74PnQ59XqEFVg2+85zxE5tr9FSsPs83Gj6YGcSmMBZJxmp/tgBYqDk6iTwJXvZz1i2Zd6bbAR
kFWmKgQmHe7bGDG7sJ0nUR56mZ2i6r9fTuFsIyLWQyLlBYLroojSk5N4aywt/yBzeFy105ZYXBDU
8Ryn8DJNJaH9cmFtA5ccQ53v8Us9vWJU0ddZMtUdT+iaWUtUFRr1lfANBJKeL0pwSRgqzPz3Q2wJ
/PRdX+DXsYT3X7rSukjCw+MmylYXKe5uD5Y5BMmV9/mFXPbgtdXQNomaT/BWSJKpxnz1o31xmXtq
wJfb5ACLavqr7aL6f+iFoDkYrjduPlPqcQ83eSUK0FfauGsJJPaN17oaPpv2jniV7rjjKTRy42At
oXZDvfxB61YLit3uKDzBpq7aijxXHfGoTA0YhFYryA7tmQP9i4W0lOOi7Y+WicKzfGX16TJG4jKp
nWGRFAlsS0GsiLsoXqrzwEX8JLZxwyAf4eIMkPg45r5oYZMTOLcljV7Y+diqtzhnqvcOrvJ+42Kd
Xrvnw69vrSFP3yHQxqn4JGYifACTdiV9qgqRSjslT5hnTgYdklFFeFnlGN8LcQzHonpq4Qxp3PIM
v1v4E3s0T8COOEXLpadylPbkKVIVU6rqVBQQTQy+087GaO62sUh7pTbz3u3JtpBf//0HLZ68DKJR
6ufbOgs7T7dJjmsrD4ZyVSwr/0EHJug76kn69BPab6TI9aVLIAJ/xUFZk+I/wyDXICHRh1/HzOF/
IYi8zG5ZJGVf57CvtSaPHQNdoWZqYJEsFdGJf0dUJy/kSGrOXuCd9WnOm6K84LPCjNW6g8uwvFlL
gGn0c2FoF4JjwggX2ZVwFa5jTfUWz39XFIxZKGsAl+1L4/d6213pupao9wmgXXm9ydpDBl2K4h1e
wQx9E/nULc9DRSMiYC+OgGchXQRGguLEslvtaXTkDMx0ejeXxukN/+GCKHo9Pl6+c/wcy2xhqDR+
F7rx9HVH0cZAe3Dp9A2mnO2VngA7JlP7Ii8Mxsk3FWBtqlg++YnzcJ/XZt54DBiV+v5v1oUobqqX
z3ZrMwqCxOaQGgR/x6jbBj1kPgD+JvD8NykXqraE7VEZDwOyCGkXQHrWvk7We/48QcGcQcYcwT4Y
yvpqfOXa82omYfo+Po/jA0thf2+Uxx5hdZe2rM4mtyw8XEmJ2SGPHh/1r6zuD102dxgkvaA8aPNd
TBGgued4SNNTdIddgq10rERn7XRohbpwPrreGCfkNYluk9xauTGBkPgw/+VsGSi/9be0HBu5X3W2
TAtY9Xc0t7ADfl92bil8Fwv3AVP1I9nMvZ3AAF6kjuPQiemwMVyVxzY4dqEEPX+orOOMKKgciDn/
xX/AwhRk5mVi/1X7v2i4Sde0d+OOrKU7oIv+LJodzyeii8HfFKOKAKZsMovubTEF3SzH0OMliEje
uDF9KcrocSnIcEhqdRWt022OZzKPJ/BMspRTkvSjeA1BMmFAT9eHLadT8xX8OPZfF8DiwTmwKwWk
21w9dBPP1+2DrEdz8+BgrOZDYJ/DgcC4On96csuW9RMi604XF+/w5FVsIz9123bb3sHGO0Nu7XzX
l7yx4U974E4Wpi8V3new35yaazgMs52xxKfl+TGkinF0cGVqPtM+pR07aV0nT46axdyzHdPcTtxe
3dDP1ArFizJDujQliVbnAikvMbfd0EHGdWO2AcJ9f6gJrwTmQ61djHg2wiq8v+zkV9XNt6gqpEFs
FlNBEpjcwIovLrE6ZQud93WQez72eJOjxdict3ps4d0cVVtk/ehMuTE1gPjPY1sQy5MfyhK8oCsd
ADOJidneTjU9gag0z4YIA3sptUtpgTA7NMZ0fXzJYwnLdBFjJMxSF3OQdHHOdYzhZb608gFpoBcF
x2QFmhXhmS+z6nRXvDlHUGJulEqcPmbIrbvZ4Nfo4cllh2k6U8KPR+/mw+02G1HOAjtmcZe1J5Qf
D343+rSp/a1bSZLI95xR7Kh69UinUclNVWBHlrGqrdxpvZJk/MCYGSyTQkW7VD77g7dZbKKY+BWm
PNqAbBSQdZgBsF2adZAxgEOqyoyskAW/UfjCnHaeb2WDN8Z6q/Z/qy61JmOy9HNxW3xB8VGgkv5J
t5D4hSdjRdJniDrj+rLhkTrQ4Nf/+tjWsAfrMlI5e7IGZGCUBvsl8gDkaOwGgAQkpw2EQgbj8t6d
O5X//4ozuO3zXBFvzMJ+yoLlvLbs8jLnT6x013v7ftrpUBm0XIQxX5VpFonNRmI8CyhZlL3IStVR
m2XMNoqowKQ8EJ1XVi2kGrxktSVHru92ahrSmVOmoE75hGECs8GsJ+h9P0P/9qmzwfFjF4rOZPvZ
NonnO0UGjuEXvca6KpguMHgGUj4eBVYt8FfM1bjb6sJ4dWP9ZAYII3p4QR3U5Vp6pW6YmAYYfV8M
eWlzklsaQ7erol3i9aJACGOrScYOjylIvFXORhbRtLRZelgIilf/R9vGgO2Tyep9qBTTo99J7/Gr
4VG9e2WSSLRExtrHvVRTFOcV+CXpG9bYhFHzqPB8PZwULyVqZKeGyRaV4zNvH4ULS79C2o7NLif2
Z92dQ25/m9f2RqCXzL1XIgQMdhwTlDJM9FduFA+570Px/etY3fPNNZJdcjHLTDeFeppFeKts5Vz2
5Lpg52G1OUF2Gu7ns0sBcrCi9fiv/GkOl+oHcvUSlSmH6IK+y0pJJqJpCwNPOUVFxX9NPPZRiWYw
T3G5kifd/5v9unWzYcAnGGP8dBD/dBeBdL/0457JWjMGtkpyyFgK0MQ96+rGmYErtWxA4JYHDI/c
X7BKRkqMNL4KUQH2YOxC5bDqa0vm3GDqJm5rSGoToU05QZpE3Ve6kKkuE2oiYsmDlgoOH/p1SngZ
PLP/ikkNGuWAaVqdvBRpk5d+bQUdac6DziShRPB04bSr9xWCml0pePrpRkJm/BPXUFJxzwGaoYR7
7nIjwZngutIzhz3hAASCaoDTuScW0kc9q9z4hW5Pqqxe3JuFH27QTDHu+W3bbNJgXO/+PLMqQws6
05TaP9jglSNnRMKs/W3KQzv6NmNyOtSXfU1ndh4eum1HK6jwRBcboKhpaRvro2iTsynziwXCAewZ
kgcyakSLqgBojp56RTpK6xRLbaizAjkvHD7ChZEmtD3h7epUFER6Q9XpkOOy47Xu19fV8RVewQ6k
QAsOX31SB1YCcYhI6wRIFlgoee3nNQqbsrf9D7Y/jL5qAoRTrjt8X1ZJN94D16eCnkQo7ewHSUrg
5Gf5geFkS8E81WMQyC4E7xK3Ixr2ckMGP50GgsLaGSV0JNRO7w/Rbq501uSrzTSy2OizgKR8zQgo
tsK9Yhr2mHY1XMefw+iotH4aPcgwkdwTXIytTVYbH+hCXKJcbRSNsk5C0xKsTtfyg3Mu3RR/jjwo
ANVgqen2/+qonSCfyLHPtpMgYbh6/Qorx3EH1qUKVFitTVML8EclXNInD39SWV9zdh8/alwYwU6r
Wh3n2/ZoyqVOGef+PjyJ2Tr4SPgOxpVbTzdnEMValDY1t/nc2IkXhQJ+wmaNZM7BuapDR70Xfyi6
N5eSfO17rxPB39N67QKUGESyWH/Gpc6FfBUzrYSPmxPia9C4Jrjem7EqUeHnjzHv+XP9UewIxS/p
NjNPgru2t4C9qW7rAPHg9r+RUAkuny/p0WPko840UMRgRFxsVRhuqVeZYiCuBQUhiBHrHvbtH/t/
bHcMInuusoEE+4W6RBx84LXoSDrxfSqNUSFyP6R6QEId1QdujHPiflYrQh4BLJTCi/b01sdNfbU0
HLO0turDnO8KnGVVXsAoHmvk+DAT/FhGl6l+Kgjd+TcOc2nDMth+TCYOZmIkagn+wep0n0lGV702
viEcSbioW49Jizx/D3P9rZAt2vseT+uIntovcuo3Krq9zSPePjJUDxpXUBJGiIoT7wSygKecZbJO
34anh+zFsaeqU/L/i5NTiTF3YuyrjBPS/iELtAu/OwGF7JmP80cMrHzGorvK8wiMI92fnCzXc0m6
KUDcc82TapY3faenRmtPjrK8vfnHtiUXvvWRZ5xXKZkDaegPWxzze/IlCYpB+yoVKytAxUlEgidG
z9M9mnccmRfYRr5L9YkOKiTxNcuxSjFjl7wjtzFhnRGwXh9FwwRlLcS2pO+zd9mRm1X95+UOgLAG
FujOXRakO0GlRT8AJ5xMdkNXxZOKADhLyPMEqlxvGf29mL31fT0LjWUSl2+fkqeZlZt7/bcJKTg+
zbcd7CY4dzt7IZhQXqt77P49rQKwKcy/khcuf2IjU/nchhUa88tOYuVyjNIBPdk+Lvy+7Nn8PAuz
GZVxlb6lJ+PXZdy+67gEFUQas6BW3qpCtSi6xYrQ98Y+TnhiMbyH5ImeG08anzBQmVHTIMZ1+cVL
Ur1as2ZVQImp4zBoxf8TT3dpMLwdt3VcRQW7xem90HhL69g3FaRdoL+3+IK88ndrYD9r1606p13K
yU8+yfG15tbV7e0Bbu5uBDaOLxH9JBc5dmltnvYIMLjDGcUWiF5T+herGdZD9GwLr4hW/2G2hIFc
8XtdENmkvv5iqhGdX2bUD1DpXze9zw1j464QCxZAts/Y96nD80W5BdOXR/dJZemMjlD3K1eNdc4+
SGEiDnIuKuxGuEZ77eCnnUVKyMUfmBLAskCEjJdlWV6GycQgMdbyQqFq6naIy3IvdWrJOlm/y5AA
dYEEgKSjiWqRJ31n81sjrnBOITng+6XaqpHqf0+S0fm/QUw6T288oVhk3qA9/q9gxdqtuZx/a5s4
TUWvB7Quu1WbI68qMkkBlUyiJqPfvWd41Kc0B3qhnGjvFiWWyEBBlMv6TWGBa7nZZdijAxDp+u8+
m5425TLHqFlDoRkv1jvnS+Q9JhzQ0PMtHmUvs39iLWz588dLk8KjdQvbGlyL2p/wUc2XrBjWXBjr
95acSkIjIAOBkdYCQA5t9ySOy985uvH5kFfWhfH1N6KFqdPJ9tbvJOIGNBywNaPkgfB5bsoXh8Ce
zYMonEM5AyA0h1akhUVxiRzY5gGknBaR8a6y3qINZMk8vzzR0vpkXxh++a6KrA0Gij6AFySY09eG
UVISS5P9nOR0IKbrZtqDEXdHDcsCDb4J1qf0B9futf2sfAIlJtcUmRJzrcsKf6djVC0LcCFRL+W3
P73gIee/6ZGNvz14svJ7AUcuvgEICL5kaQCuU6i6JJEFRfRfmVNOalpomb/w9renizBO4b94iZia
v1cLol643g+89Y6Wn2L6Z0++ZfIKsF0tPXB4cZS85nI7cTxJJu+KJ9r1nqK9LZSah5/ECtLG6s6x
oE/APWUEAKrdRRbDxiT+aOdUbsVVoUIAS8cfcQ6a1ycqTeqM5lnB7dnvN8IK169VBSLof3LhsRqE
T/GZ5YGq33buHLo0YPBuAwE/P2zZEmeL2czuOVBGvEAPJU2zTCnDXmG32ylQNGYMYL1rWxG92kgD
d51gBpQ1o0SWXSJhldhEU3IsByVogaIWbOl+e70EytjIgQT0zm+4ZZRd04urjkoRaE9P3ThJdZ1b
q1yBHHoA+7cnwNSk40I8FXjZUEhL1b+iQEtL5VziD23182Di6NsQe7K+Tfzl/ARwoxnDVvszq+cj
0dEgLe9Lx1itRCF52sbcC/HwVeR6s8b9nB3p/eu38JBaXMDshliI4edTw8HQoPjXWBIPTM0yuFbk
4bkWmgFDOKU4YaWMGMj6yjh3ZfrP1H3DYeBGnWQzsdl25XDoNbXwN8pZA6I4S62GTeNNX9T2pDBs
ZsY7w64zVDn4uUvR+O6u+WfphvTMGaBtgCBU+AH9KRE5NMAWT4whginZl9ewdCvbyvcAJSSvSXTZ
v32Zf5ij95z4EONk44NakU6nYoQKVYYHUUFQSM1gGSn7jotMjfBGaJtBx1OWJsA6DmMdibR1SiMx
rsSlcUyLKlEg3Jcu1OiAICnv2rDvdlQWuzMtofWN5SDEK3XW32Q0SmVce3+d50SEn5GoA1oj/NLc
7jRpOgbfj2FlNAD7BjzwcGKGb8fJGYtlveQASZVkxwsqPOzPFUwIo12NGhe14kN/BLvH+94gFxwj
vnIJFQKKT8rvoRRnUvUdRHyLbs+g0tlyG11YlnrIxuvTS19qDxkHeltOuv9IzgG2/CWx7IV1rNE7
wzR4QHuOrIqnkxCAMpBBDoVNWUgVr5zum2QhKs3K8Ga163AastyIZFRUxJclPCiRQjb5pv9EQtKL
XQi77XX3VBQ4pAztHlEX2MAsQn+B9R/kt48FrPmmUYZCq15sBBJCaMtqTULHKW1g7AHI5LumAT93
Orfcx5n4Oy2CpeXifwmEKscDH40JhG0VnkVXzcxXRvmsG9moBDg+TxmN6X0rqsT3hEjybwm47lQQ
ItS17nIHBN8rHtFE9vulAdMJSTMS2nc4+JuhE3h6E1aSHKT3WJUWTGxJVAagoKS6C8oxaCs3a+om
fhplFS27FTBTxlHCqoOzZ/I3Oua2x+ktuxgFRCqqkdTNS2HY6iGUTdFF2WylSlbyRXs9iszQC3h0
QGLSttqjTOAVMufynHN5RH1rnmgEBCagfjFI0b0qVs4ChM7lhH8bo/fwELdqn2VGYUqi9bhwwDAk
c/tDWc99T3y/ptyrdL1ackYllDNpLFE9iYoVKkXMg0R80uJSuMkankZaBx0wmug/Jx6d6WXfmBwP
zKcFbDydTBqJszho+p62PDiSn3Q2xf0x3rN+fPJzIYGZ+46jwYeAcG7Uo1frlW4fhgue2bW+N7PA
7VLD4EevlAd49aaVxHVCc3NCCZf/oDVD20Ehd8yztJ35wmr5XMpnMfmueOHnswLPDhtPXBEeYIFA
kABTMWYp5BffHPFHInALW0VMjuSsP4mErEHR/ARLVMdtOHfJYsYwIqcepjV0HNDyWa+RdQXA59dd
nCVtXu7raL27JOlXat3vmV+zbipdIlxtiol/WS3/rWPu6k3FzgYLSVlqukY2t8AlJ9n3XOLnCChf
ceA/ExA5QypzvirDmY7FEL+3/r5Pg5c4V3e15mdUuDcdZ5cS5c6tO1qoC3lnGTWxk1R9xCpBz+8Z
3N+PyzCywjU+bhUDWGbmHMiAc8jNxiC4wPcFg70/9iav3rptJm5/VkZOvpk94ILrLBo/1cV/Xrlw
7fVJP0IHQ2qacSLbo2eiHaY2/AZjANMQCvb0PQWYEEiSpbFVgxtriJsp1qq1Zg7eA/fOf+rrUvtx
Rv+kH1j1lXqAiPOlMTPZV+lw2U939GSAxhQMh4RQ3o3Cjcc0BuoBRzUMhJVhsiCjGFx1qFtes+wV
wj+DN3YiWq4dSwhbVxiLb4zUT2Qb00qUrFSsYdC8wvG3zMeC9/NWmfjNDc8dF5e892fMGMvTzG/f
YFXGX/6UTFF6Cdy/y8G8V/zVAO/FBPzKqPKmP0dEFZgrAdA4L5E6qt51eIUX2TsBx2SD+UZN6H5f
GXJTdwaayOPBiBkHWo7ROJP26V6d2hIoylg+84gV6gozZoZFxbHzJ8r35gC43p7lCBrQ0rfFa0ar
gVEhFg/mo5FS8fwT0iv0iP175Ioy9fXQNRBaEFqKZKR0KuDfZAxRp1rAC7A9sz71OOscSADYCP1H
+atglmpqpBbgP1jl2LYIyWEQMj+UP1OvWeRt7Z6Driw//PRnTY9G+fiiSTX4ZjkDCHEymrBfflXy
JQEDJZWyWpj6B4d+u4yN7vKkql8e6GyONR7GveC6QWKl+sR79gVbAOMha8bv9wSZKCQO1ugUt1uZ
hE36I9fxdos4UkIlS1kQlBBoEIwQqAijkNrtCZDD/NWv/lv8s2HFeiaBFW/lAsdvHujGHZyIvSGx
tcXgPc4UrwubHA98Gase5uC5nXT2iBwcymGm/18+YAL3QRcT2cTk06fGVG43TrKGsGc0sFLzTJsv
PvZW3oAn4IYEkkYdI7rBEXU4zXjeQSGb7Nu0JhJwVF2yQ/rOwMAGgawwd+OG5OomK86JIQx1eWZ0
hsgm0QyrJH8WbdtBpW0YY+YmUF3WWWrjclk4CDpnC0Y+n5H+hLs4KYzxwJkm6Iwy/iaa2GN0m0xT
OF3Q+JSfdQkVe2BIXf4yPmzz+S7bNbG33WiCKI33KoDCWzLBn6mYrWwO5zTKVW28bLEUNr/Lo9nT
3IFu8DKAZMg8V8eRVQtfti2ejGRhJfNJnzyfxpUwy0+j53RszHJA6xK5KbmwaCDzshveLvNRTRr4
Li0p5LLAOENTg3VU7qdsOVcH+jHY8EXAfl/YUMK+9DHzbEh3Nejk2cEXdU32Nadvc4/IYJ0VSfgy
V66C5bxiukxSw+XVavmSJd+JHwgIr165DMFuFBdwLjybJMlPZzd6/WCIbrwFNwTUt32s+aY/5Kv+
kc6nh5kqdMbRtbHUtuFBkRuHzQsdN5wsgJXKBHjC95lvuVgVsLTpLZdeJuxJQRl8gPYgtr4Y2sYn
b4LOjVyHZ5pBRYPCaIv7XhgdvFBpAKDJAh7Coh+84QqpuyOSlwyxe5WP91d508/dX0WFDlnZitEj
Q0pQIjNt1x1B4SfrKX8oRNz1CBjWKLuKZdYKbYwgyk55rIFDwtmrijYcT5cf/oaR/dE8kUuFr0Mz
BVfnPNpR34dQvg1OUH7HuHgQ/8PVfEF+jPtCFGtqxF1e6SW5RP6dbp8rRCLGBGAfq3csNqUSH9xP
Q7IaUtAEqWVyv0siBjFReAXDieegyiiZiQ3JCLY6Iqnq0Z00mFA4B5xEo9m9nf4w0XIWLm9eliFI
fFwJnswifcgR+tS4tcOYZVeAzy1nMNeJQcqmY7+8oc6i0P7IJxGIpRbOjGaeVkUqJlsW8soB53mg
IqhKM/1JXI0BMPucbxDOI4CrI0j6V4AizqiFDuHlKSFkCmG7BK0cwwB6gYIlJtQti7Hoi8qmVmux
fvQPaR/N5DVvtJKCV7SePK4mkwP8HISl8Sxb+3X+rhkOHYJM3AZvlT9NDVCuSoaFcQ6RqdOu6xXc
5vvEKLUFwLPFVmr4dc9R399wwvZZ7Y5idYypwW84bV91MQyu1OX5Fnqlqxwo4fNla8SV5SK9ppL9
7AAX3gtfMLIlxc6C9u65xcCL6eQeOuer7efnxwXr1CY3awDEW5F07dRWdZPok7i7TCpM16QzNbpj
OL0k9S3WbWmWNclOJGN7WMh9zTmmasMFyOxTq1owOfOkTOCh7k0GbcfKl/EWk8CPDEnEQEZ9/lH8
hXMrm5T8OZZL0/KPwVgf1/jtpVKEBKfA6MR3mz/R7J3PYmu+70Slc5SKZUl8fwi3xW8T3ZLH6mwU
DQ773oF5o1+0RKEZiKDhl7SzkhKRQg/lJH1Ekgh/l1PeuE/R12zIfd9ygB6ZOQQIfF8reAjSqyQd
JPT6BHIT8MtWz233UVpmpUk8Ea1oEg/eYnfwseh1Ib7r1jNdOFKr0WfGagaITaJPdjm3Y8/w30jk
V/65muP/UENha9HM3P3BiIQ1k9Wf5gV1Vc8cvPK5uOHh9sNvbnra/G7whujVjx3h7upaDIVvaUkC
i6/XFIaQ/r9dOC8xf/twY6VpJ1SoWHrc7J6y40GRqCQC6OIpL3E3UjAPEeC/RwyYQ68p9tCsLOYZ
glWqSbfa0UiOEpbeQjMQR7yayn12eIEJruIrtJOPu2L16GQCnxiF/fgYf42BHzUr0VmEm0N+3tkX
Vtlf3tyjQNte76M3Mpwllg8ACrzq+0x+Wmc+N6TxMYh5psTMNw3tsWI99Rr3DIdJNs+6lpF5GQ2F
As9hGHiSWVUIbA4PRCUBV/6R27g9u9GSpvqA5V6l2RCVS5fvqkhlxlBE6ductuW9GYTf3+6D6xH/
TBuFqzOmGpZT08G7zFCpzjH3J+lMpx7hRr7mFnW57tKE4FWCar1pAFUpGyEKuJlXYuKugfl/Vl/T
5t6J8f5/HmaSLLXC/SCH1ulQj5FJRnKPD3FNyH4KPW5Kdzd1HIxFnre3MDUtQG3tMyAlCTeOsJ7V
rrNS0Zl/C1FLggB1dnfiu4fkpWP8cXht2AOkBhxYENTl0uOSDVWGFF6otoloi/z7oxe06+UwwhgT
qZNgcxJWuC1CmblzoPWNw/nXD9yuRepqAQWUOHMM4u1t9EjjbqHXEjaE38RM0/WryK71DWOMJ/IP
bH9c2hzjPL338BNpvL3aLePrxk4L7tWE/zET3TWmjDmsXUSydIHoJc2P2pRBW9xyxTrr3JMCP/sW
x8wKkB8IpQz69ega/jIRd5hp7NwRuelFOP5oDj7siWFaVB8QsEuZeuqTtmD5tVUI0MrvlxaIoDin
wiGA+2IRS5e5MasktLrPpawSVcB4QSI7ZlmAETmhGy6jTQAVOa1S95dNS5M290Tg3QiYHCUyasLM
YDEBogWa/rIDs6hsEGuWkUp7TVSQbNWJZRmTUNBnEI0AtvsPz8Kry86UEClJNHX62tdkNF0o9rUv
R4Y+CwN1gBh6elwfe3zvAWiQaYsrLbykwPriQjtPMue5zRK3KydQd77+1NQ6hFtkCQ7taDTVpyih
t3NSRerg9myPLXl4ghrh6pyPQsTqSbgOh+Xw5H8erpZcvGEOcc7bOZULYy1xz6VrC0bhAKNwEq80
1jyJ9EtW3BMYvXy46JA5v0HazNVG9if9W+RTn/X8rVjGfzby1Y9+NIsEDPYW76XHRJh6TXZ4q8Kq
7RmdbxXI/rsKThy7hAdo8zSBWQ6psyhLOV9W51hdmvuX/+NJJuMWqz5dqdc+n9uqb2kXvft7gcTW
ppyvVU0OZS19tOAWadih2/QKc9LwVP4mU+QKhXmd4z0wjUOwzWTrkQBoXB6EU8rsD8Qn3jf4pKWd
uGs+FTl09FwZIF5YuFp7bJ5DYKmF770YFgb20mPpnbxws5DyZsDfq2BV7w8vtnV31d0Q20HRRoPn
1bU4bp8gFiN/VW9p7mfIHG3uw37PIdnnf4iT41VsGysCuGyCX1KM0ydk9MimsNXd66VRZMFZac6C
YwZdlbWp2Sx7CHA3M3x2KPBVploTY+SpgZhE0YsLdnhAATLDoh0sbvw7c/AX6KCRFwuf/41ZbJHP
XL1Nndm4dTdr+tllesL/1igDzysAqD+yTxRuju+M4v7TIcq4A7xKNwJtXOcYt4YUBPKeUGqngz1Y
C0VbiXmm+6wgaY2WAaq+eWkIfRj3ybzVnd9r8RNW5rJp+sCPLLIhmWXGUpet/X8dVExGIOZrU8N6
qMWN4gJVFmKhmRLzSs6/343yv5MAEPnryp6o8PgSeG2bCjAKVeqsJ84KigcWDenuTyR1zlao2umk
rPmCdqGf1Vlvi4N97rcD+dOmsFa7hy/jLAa/HAm27j8GrI3j+UEImm6+gZxL71c3oomsGIKhd9d6
jacR0e2nzXChXQt5RQ2z+zm3nwDbCV6Oed5ouLi5g70RvlLWHVoeROR3yyGjnPYT7id/ZkTE4P7c
9K0CYQCJPIqqbzCpPJvqn3V62qKTDwTzb51UU+3Sp7g7DqQ+AgdmJPKINGLw0sEB7xF7ONCtV8kN
pGewprqbHoC5QjgFhIngFG5qyNRRAIIOydgTnnlDSYpRuq1g/+3gZqbjgMthVPmj6ehddxODARt7
akwFNrljfyTox8iJwebPleEaQFv69HvJRiHYSPlhsYMUZciq4xd67PHv++xHPRhUGI4kTvVxOQeH
ZUhbAlFelHu3/PSpfCTL3pgFPa+02vazSBPeP2pDSFgIOSDL11LEGyOGqeG3YSOhvuoneYYr3wHf
wgLhNEasiK78HWuTqhnaC4lvlBVELt0WOYJlb7MHsIG7m5hiPZH9oDcBKluumhu3P53ggHkbBQit
AafF6+AcpX7r/hy6Rudzd4vUWOneXfYYBs5KQXjws2kAXW9qtXTeNyyJ+p3il9tkfGi+G/ELJzRa
o66S36UAw2T+erhjj3Qu3wm7Txoh+CAkawoRijQM0H1qis4GZ/B8NY4vyoY/YkiUhhJGk33qB9OQ
iRyI/vLEAIgkq3wVvtMI6fd5EHC80fyVlX1YYnCyu9MDDJ6mo2yON5fGYuNhPKE0D5i/LSNCAJ9r
VwTwad0VN5X88K+ILdRuaUKqxkT7EXrBEr0bFDwRNtr797o7OPAfpkYDULrV9OEG49w1k57hTYkn
QfYfC2EEF12uNt70Ch+wTjhcqGMTRJouUC/90L+XCDg9bbT/FZ2UNHdevHpmHbxrHlOY0x55rUeu
5j1tVJeW+0V28wa9soLnASEEIsOis8pDCsbo5xiMR/R7wlNEFx7Mo2KjEbOKsANcxd74Og1RN5TB
ywCVVifnr6RoKPlnpwB6lDRHijLsBCFd4BL63rtwkKmJlhCpVwzpQhQ1I8oN4r4fHV660ynsQMl4
IaeK2B0pK27FtUqpDX1Ga9imMR+17fyX8oTbXMj7eiQfNHMlVa6MsYebErUq7NVirAZKkNdjLckO
4V/wT1SfP2Cce++WVELck8w4XU8Ft7zTospwn6cz28/4YgHpNSl1771FBatXSlyX4/lCfbra2DPj
MCQEWR0x3a51sg6bp6Qr43pvO1fG1X9eqjrgIHQ/BmwtRMftn9yigUbMeB5nHexFIYNPPesdvTV9
bZRFUXtMud3bder8QH7gvTf0z6AAjkACz0x218Qct2iRm4UNMLsgo31GH2vFoh0bIoNaykXP7Jnh
S5GAGR0wjtsE22QUQoLvqN53R4ngGau2QDLJf0oSBsJk8EoO2SJYo/eyuLZg2SE2+1m3CgnS+Qcd
XJVI232ijGQUHZ7yUYN6KsxmZOa/GXAcn9cln3cCrMwEwHI+wDHeUzeF63PWrdSxZc/dsgJ5G3Nd
ZFt2s6B6eHMZIFUGBwj2mw2w0k80MP5ZfcxJED+WgCsMDlzaCncav2fb4kW6z5IsTNVYOU6NQ9Wi
mZNH3WdLwnNOWdwX4viq6pblVGlO1wwhoz7b2Bva4ymYQEbFHDOMlVitNWb+kAuAtsOiIkzLnSd8
b57k00a1jho3hq4YSBGUZG1TyY/26tM0YgKqJHrUqr25b9anSAfEXZ9NUX+YuFUNDqwqVSXb1Z8t
VtcVxQbZjYh7ZPr3lI2zZp3tRXLN/l7wgZqtLHdUqpu/lQoCj7jEAftYRQM49gtb3mTharATHSsj
j+dycjHZn+t3bfO9vpR0CAkdKQkRUFttINfsxaLj+HWnDdbeNdcqexVwT4c+Ah1x0BlzDZIiZQH+
DiuZBBVTeHofk69j4C1gW5XTai5l4PaGgIvkAhLqyAVeUynZQY6Osz54Rbtv9i7hTkMaOL5zoAps
dYywLg306/nhnqCzDlPyGK+q8EnyLnqOfUi5+tAfAeALtivf5U9S0jMz1fOrVcQmkzQ/tg5fJNr+
y3dG+f5de1XYcGrhVhs3lo60818SsKYAXle1f7eYGvz/LDukPuZpeoNh1+phfziefq4yamNLu2XF
sEHeay8m2XAdjafQDXFiKJ2jgWnUdcUQwix6XJALHO6GZ6F7M+PmkzBRuEVyF5l/iYUzsmHkHZK8
ZKL7pVXzdg99qLbc7Sm1lujbUqchsadVVYcejqr1xq91NGr+5kZhIRKZQw9y9/hTA3wK39M+CLYo
Y5YNyzoKFd8wYEY5imFO/O8ozyp8O2bz8xosi8vgQSNqxXd+iZZxsrkTKWDpGkt0+T5iWuWohyjH
NKq9DOHw0gEguMJ7mH7DF/GPLX94if53Sskm47T4zb6XyQuvwpDztmHXTLKkkPBh8Vps8J7rdsy7
3MXlB57oQkgAVOLqTD4D7NLwF8kHgwwHBfSP7GKx0ZHuqKy2giYfWVbXCv+pzWCNBXTxhh8dhaG7
oV20KAHk0FTtXl4IH+6amxDuh1TqgBU74FusK0rd30QYu/ZZ1LgU9YjiF5RUCm/2aLXTbRHeWABy
JXtOSvAAQgqfudF5so8xdF0v4g0cXR3iPzPeplS+jUF5BBYApILUuKxwU89ojtcwm2flpiN4gqBT
cRUQDJepoUmJi1QH7l4Lth6ucdxPj+TOlwjpRbLroldbEDWqEupfZZ4PP6jG4pULZyftZWgsbJhj
B3A0+kk0yed+gP30diUTW8Bh7c+Y/RmG4l7G23GdHb6lCcVoxnwWh/mpYVliByZWuh/z3fjtoLub
lKLS3GwRJ4juzsUWuZhxNYDZZHJNDtzgPiSIo88w38UmDBUqz8tCRF2vWpoCtyyjbhP0DP5BX3di
j6OcNf6ViLI8OC5dQ0x0SbHjGjWOWxFSfpqb6w5MCqnHphuwgh+X5d2OR1JvnTmJivbOWY7XzUv1
GDjgdtuvhf+UfHwou/fMhUZGMttGnTkDct3lGwN0DcFx1TE3EZPP42gpLiwq8wFD2RPQSm1yroYW
uaUHll05WW5dSUY2SxKdV3YMz9Qnlyvw/qHwEXr+zbmOBBx+LmA/OKu+Mqch9C8Y9cUkYKDBB8/X
lebxgBtHntiLWBzb30wcNJxxscBbzSsPPgB4lJq23AEJoI26tSJUKKEJWB57BnWwY39/WLhSW2k/
dDVSEfskG7UrbZvfm+GJvNw9GC5UsxL6Mt/Gh2UoODb8KkgBn9dsvM8H/YXtz+IXXzWSHs3osPZq
eXX/VeQIckFslbEvj5Vv660MoIZ7JDoSQ2G5qtxxBlwDgeiRRLrnZROxJHP0xSJqgbs1aMHoj7d2
8NCsi1sMFSIUSouQdnVZG3xDtv/WOk9J+qhZOiNXzve2wRNSM+Wf2Bgr4fVrYjDf9PRGyLFkIBfH
o4oo2vx2xWH8M7qij0mUYMs2VQ3mBBYoN/bFtrKt9paCJEB2eKvE1XS98ylvVsqlsDmDoKQfKpEi
ZF0ylS9qsCMk1I1JLodpyou9aeCv2HVPYa+yBTiQ9FR+G7bZVP9scooWEzeTFK5NpVzLXwlpWH6o
T0gW60QZ1vUmdTA1VZx0e0On7sG2ZssADdskMAtZo3Nr5q7G3ZR/z4mHOCpGjaC7mfT/hPAvo93k
mgtHgmZ8NPzbM3NYurlMkl7wYZN3XsAmbHac+yG3wYLJXrjXPT18J8W/1Q5mgEy1U3+g73aZ6lDZ
YzURCev/zIzpXZhtweT8KnKftuIoYu7xTsMQTbbBaHz4tnEYlr51dkTHmIurO9L12aYtqXbeZb1A
4er+Jt0WaFZkmCnf6KCywbjpxK5BDRL1hRR07e5KB3i4Y1FuyzR89EZGHj+HCpHLAGGeaoUbfTer
RXEEi2kfTy5tiOY8Qldm8glukNyt0Vi10Zx+f7UQM1fM6OImvzvfYOgkRLWqj005YIcgIMgoytTM
hldLnurff+8sYArhWWBb8bNlU8RgJ1JRzD2o4tPJadndSFiXXvkN35kZh+xKBmoUJkIoNyEibrXg
HCiZiLPo9YhuK05UlPuqWF173T0lxlN8VRE78ERdDv5lh1CoN/A2AYd0g1sL87gx3fn+CLmXhbpp
rfrZztdxW/RkuX1pZEnTOSn3sVwJ/9a9vTgmSrop9mzpY9FxWAeKf/WnckkpaMWQ31qyhXdvbpjt
S/5qDg9uF64Sc6dWN7G5XLDmSSiVydhoCIBKZ7SRwu2emjjQafNuNzzIhTnY8139hJCYeFIhmHfh
Ygenh+5P8uCehxnEfYreOn/qNonlFJzRQrVTAvWZHhVhbr4jyJ8vjwbCSCrUTW7rt3F0CYovpu6x
P1rvZLQJefc+29hGcpaF2DroRLS4cC+Uy3rUd5zyS704YtTtVGXQId/IvCIg0iwxKffjZROfCs6d
071U2BS6P6GCUlEcGgwe6+k/P4i5J5M6NGRO33ut89V5/r0Ub5wscKUP2bqR+CruW58Mn02YCQNA
vY8zBQSx2k2EOLwrRcYXuJtODdfsjfTvLTT98rL8Bck91MjS7ONLAba2v4OhZLEFfUk+8v81lBK0
foH54eRHljRe2juk3arYFhXLy2pHxEYnCZZNiT5R/crohlTJVRz2IqWvyz7in26smPCxY4KLSxPN
4BVD3ITUipFNPFtQaJDdCIPuxisP8G/Mq8LVah+7rQcTCjL0lLL6uO7BdHQnAWQRGgAG98R6Muv0
6YefJux46nTSKLRo5aFmcIORYjOhas0rMdGcEE7kUAujzBGFvv01nCJFHV27bgX2oNAAQ2YcJhet
/ixw5e7Yd1vtXNEv3VuY7y9/cJPotvoPL6NLhBONtiq6qGLFs7qeuXDaxoI9X8reapNpx2A68dbC
0zGG+Ne+fDd/h7HJRDn5xw8cwODxhNDemlSIVQXFhdyPNzjiAerlRZzJrc6Z8TFmek4vc3WAS513
OZ7svFCLOlF/5C9fjwX9CtR6bKbXPSxeSG+I/u8EA1f2gP5EcmGXEcii7euST48bL0nPIZ2FvC/f
abeDDSmjcErgALg8qkKU3seE02Y+Yr53bnzpjyFF/cczEiKdEU06EwL6gWTbuQKnxsRmg8GdeJEy
Zk4jGFS8KjjhTdYBwxzIeakGhWswsOUwqzwOLPLKYSv3mfKWvZU519kIQyV7zPdr7q0OLgELqcZf
tLTE+jpTFgRGRihJJsvIgZnRxXjxdB6YBwYabpcSczI4usAvfGzQIVmko9V7zFd0W4N1SyPIrD/M
MkiUzXiXJ6Hve8ixcYm6RNx9AWSrc/6/YgzWRSrRucVmkzt6CPiNveLXqg7/3AjYVN2oSxB01cBd
3U4UkKoT6ULXjfYgpsuBia7rCOE2/2dsGml82ElMrbQ0S3qmYrlzpvTnJd6eV9IFcVdeoxrcHSY6
sh+vtY6esCg3j56vTMd9MVRFgH0iafQHyimRoCY+3yvNXWsDIGw3cp6NTLVAx74yOCy0fv56upsG
NFBGw8ypvJrCkuZ4NQ437Z3zJwu3iya3hubyY9qGHyhFV1xrDdaM1fA3mCgXqFf9k/hBbzttlT/z
kRpKEoMoC/I2C67MQxurTX03tKqJTZGD9pr6Bp7FCk1nftrOc7lo+dJdAT3fc0EFmJYhkZs9C+aD
iQl5xYvVeiO18B9P+0NuPSu3jerUajjh05crXx5kCXNbwRjo5kmTAgoJzS834KxejZ/F9eB30cn4
hMdMU4xCoUay5wb04FvaxZo2BNCqel7/+hFrawFiFPJslpfZ01aKRYk1aj5htAmGWgLrtsDwH4yp
Y/74zyjRnffvPp66b3hMhCNyZS4Z2fxpLPFeRobecw/toL3F205LkfUtGpzbv0uOglMU6wVR76+r
PNqKqBcFNanJDTl4GoFKBY4RfWnR20zvJZlMaDrHlTy0j2X9Mljrx6Pmzd1ysWCDzqQpd18uT0YQ
23n/cAzACxKc1cK7iLmbB7ViuFLBDaNLBUw3kYs7MHm6PloEchdcwBYi4bedZqWj0e5IVnkotolh
gLbtTT/Tczyw8GQ+AZS8MbfhPJbBzS3tjozHHzTB1x5W05WY7SZDX7OjZXCJBfktfmEFm8U0Glna
JJeiVHxPdT4bThWB45Kr3oLOORnoS12Qbm65x/SNXIKmUY4q9J4D57s0048n+rhPTL948310k59E
tgoDDHfeMhvgGSYbhir45pv36dfNOIFy/zTOCqWVsViPTO57KsNzSDOn8xF8RlL82HcKEnknO2hi
2oA8GRK1XuM574ypwn8gVUEP4B+SBLiKaxiSylrWLZUIcrvezQEG1wXa+cXIh8ELzMGq0tuq2mCW
xFegvrMrWdYPF7tLyqgskVC2RhzOWVGjrs/5Sue7MwkLPF0xoE1ziAupRx+usJGlDgkAx07Sf5pS
YaBdkLBrXivH9CnMRoYWMUXGxZhjfnfalv3s+9sKArOWmHMp0pfJlCeaujJl7H/ywcVTLbn4laun
4LqWW/lxQnmK6xkZj70tGzVbszKLX654NZ8gnCmnf+9KrT7wU8f7ZIcOLzjZXYpdJXzRB1aO93cR
AkHQ/IvzLlBRaYiw4M50VBC/JGbrZ1fYc18NsvTvd/bDbZ/43t9hgajGgfUGuo4/CxJlYfIyJ3VG
y5aLoBtkVWQ1301j5HQdWeg3dijBzKLzaczOscLhao7N271PPvJxwWsLh/GSWSLh5SBD+hLG/bFi
kOtJC8fyM7fTQfCGQPmliN9zdJgjgt42qJ4vIrgFgmBkbSDsqV5gokV04FDlSpE57s0uOqlW4VnG
r0DbYKWIPSkPR7R0rMv51e1vlAoT1zqIJqmPSqZx0IOo4U5gI9QaQWhbtEK3PZYAmatxzdMl+DLc
62HXlzCgV73eHYTPx8FQsFFaStcfNiSiqD8EWzb0FrEMXDNkYH09+44WRhL+d7AsI9z9HaI1F63N
8jZ8q2mtpaYF+mm9/obVOCeMEMZ6Ot3X/zvSb/VuKgmhVaNO78HEdTs1OckAyFcEC0xrkyt7/L2f
hLMCL5rfa/RvkvV4C06qaWerAEEj2urAb6z5YSmLkj1yi2CFm3flBJJXUIKXAe0CEMtHIs+YoVTi
Yj1A8eb1wIHJdd2Ecw/c7U1dwGDWwmeoghuo06saSV4xjl1mHsWiN/f4n97FGGKxLrApXN6eJEdg
QkVP7IhFZFf22nhga9UjZ73RFfnKlQG0usAmr2uAAzgaB+kNbkAAYZLR2V76VDdqHFxoI8+uykf6
R+S+3rK4EGkCTSOHSXIi3tN2B91nQWwa8NGbYm3WK3iXZ7bTLCG016D9O4eFA0Apw+pI9zFL40bW
WA99eoCFuRcMhNh4CoUO8TcxTUo7DQxrmW5yH7eeL+yQYSTKeiHuvRlyYdFRIg1tEMGZcbLXAv7j
ztED6EJj8r19LkeMwTE1Z04wo4U5Tz3DHWjMPdB6D1wbQKS2J3Hj4bnewMz6e554Kou7l3d+7iJ5
qxFlIVp9ilKItUsDPJlY8uEKpfsVRJ/mORCYdbSRSdsBC+2QwcCEhIgIfpDhQg12qrjCA27pJ366
hYlWitKCfReuBRwWbsnB+aVHeQezLPKIJYjhEJzMXLdvyUElTPN7UbO/EQ8wJEJwz8UslskQXF4R
cz81YEmdMP05Ts9/Ekx2F3kwECdCB74MUNXTORuFimZGQDhgwp38M1n1ZUsIKYJx4mxUNxgWLtN8
mkjpsDxf1IvuTSNKdKvlgE34VmeXuTWd1hVVVeBUv4TOa5HtUlQjwidX/gchEngA8h2wzDD0jkgR
zJzZCirhm6gdFDBbvHlJXgWxMqAvbkHZBQwZ1DtNB6EE8+23Kcj/1RHB4mw59qms/rLurJnItsGN
sNUi9vAtWcliZrN1eM2EjPyhg/WR2/arn2/W/xWSaKo1W7jogg5uMkrHVpgjOAdG3RxIY4tQ6GrG
v3sliP9wi8k7f1B2Z7n4KZHGENp/DZU9YmJvSE07DHEgh4vvpQjCwluRgYDs+NNQZiJQGFNeqjLi
wUQYytwBdHPldgRpULaW4IqtPWe0iShGSgrrWUBGBoP2uUkaevKCt8Pe7ugzYVFQZl1x+v9irYby
VtIwLaxMZDch8a8BU8h4H2xVhy3Lb+0+Z/CgyCdSJ1TCnPk8mMhCzTYhLli6jkhjFrp7WPxUb2Ho
s6vuXYuvfFptGf3SSA7FBAPdAZGb7vV9Qk5YXbQ7mV1DRuzCDYEho13FA6vuf/hLgpxD3rFS2kT0
1YlFSojAGXU2UgPPK5CXDFcFIOs620kyeSbFGVLbtCyhA1SeM/wp3fCMfR4sONBFo0rtbCgGwMlB
3LQYTsE8VvGR+a7Mxn1HLI3q4icqRAkRTef2d+Zw+p+wfzhEjHFbfPK1WGrWyo8pWurfF4ziQxzX
Qr4hdYkSsILwGIPtrJF+KyDEuDAZpWbEcshFvLpv0fV1//lYv/Q12JAN2vSKluvq4gKVCfPV0ng6
AkPEDgc+DjbUCjX6Dr24LsEgSaH3OlIYYH1Iv2heg/28SzF3/RGa8Z3LNHQKBmpOEBH6eHzPVUvS
cbtgc+hlVTCNfjUGLZ7+32hD1iuCgJe99oTXMVHDwsJ+0wZaAfFYdQoqL+V5FB81/n3ZbyyoSW76
oYqNzfiJRYSki+MjOIf1/mJt0Lc554inq2cN7Cb9Ut7P6EAnfltX5M8UDgwMebSQKELTiRm39Zmg
6UlcreJWYAHy9ojoGm4Sn1fxkC6lodMFWC93IAoYLfP+I4K5Tu/A4++78Rws0bA08i4Px+2K4kTr
SRQ54GnIbAe41lBYyimjhAkmRN2Uu004U0oO/QUd2hFAwCky7nQI65C679suzED7+7u8y22J3Ce6
CLpwqtBN1+SSGpab4iuivpuRWerm8MjRyu6OJLktyTJQySXq2H+AHtympa4qzDxPRL0U21Z/gNRD
dvGgLWa/3qN4YyrNULCsCBSxat7MNHomcZQN2cLk4Axv1f3bYrCFcWBB01Ih9azX8h9zTFWW6zI3
y6/WchwTOsuVOTlgfa3LsMTskFMomN120/60IvPMOlvl4xKv9+D/hG9GOm+yerwFqTN59uqtwnLM
jh6j8J/TJMDnUqYJfBkqqmfG7ebMA2lJDlJCBOe3ydIO0TsMe49UjznoeSw8QVhoWuhNVSh3Ypq0
jbQSQoZaa2KKDdgsmUR+htfKv1kOVtKInV308W4h8KzNtvlPUfojOYTiKh8mrM4BFSwZ+9qTq0ZG
EOzyW+Nk/jNOQrd2yhPK70OQagpKqeFZHQUExp989vVsKIFaNKNyJTL0B9BRP8scLFg9Rd/Eegsb
aEVpONzYQMgEtcO1Y5jOS8WghxvKKZXTFPETJU9bwgnEEtKPEzp3f1w1noh94oH5rrHQZsoCYsHx
Ojgo/eWrrjeMx1XBxGp0VMuT41ZyIbY5gXglm8h1MW8sNh+nz4EOrkpBDaJGiDWtA6GY+V4dvMGv
2/fRGj134imGVBl7KPXGV3AoEzWuc9hG6UZy1k8RB+o1gSW8Zkab9EAzI11cCq9JBofeRvUsuPd2
EUSRfIgdiIRMKug8GMyHX4n4YUCRcmO7P+Kbztk7PDNwCv13Tm6y3emjR7+iVKTr2bDNek6ES4LZ
j7QUt5EUSxQz0742GfIz0e8mwXJ0pdrNutoxaXtGBz+U4BL5pEHFupZxw6M8fPdliMXU4kOSmc0M
e/E4RTIVeC94+hblMyPImrtes/tm0EZZvC88tIyJqH0qEz1u8AWG5W7IuWXv2CDVML/yEy0e/hy+
/BOQnOCLmHx+8zn0QrytAMB8g2KexAqZRptUVbrz8mIBPcp26fHFrsxFIkvVNoSIwgelJYh0avEB
DYsLLU2xQSP4HoLU4mUW7Fr6uZvjeEOddPWlIsoF+ccRIVlrWgfRgP1r45WxCn760IuCfvFf8waQ
VhSldZQ76ZRtIA9sRnIxlQL68hEhhPVWAPu/+MfcrH2bOaxpbhUsTiJP4MZJZG3GzBYuhx39AYCV
N/tQdWm5fmhPKVCkz93vY3DznBEsJoJy5PES0bdk274ihhbf4drTCyTvvBygOCedg3hfOB/+02M2
n1O0jH0Fkkzt/avaaKkiIbbV0uHu8TNaQzgcd0heNTegWxV2WJp6hNFuC4S2e95K98D0QQonXvzQ
Vgz+gy62o4/A7rTJAAN2bewcAMqmtzhfULalI6Hvhmwq81AUhVO5CM8BXsrfoIQppUHvD7tFw9sa
zGaq4ZEwLvhvJKcIw9Nu+UDg4gAJy9mAYxLIPyj3UbGoc9V+0Hq74VK16HDkYqaByz1RinyMJGYE
NdfGM0yWF0GE4YRLsDtH01pXJ5OSibhJ0bEsa0+QSriL4iqMib8VS6GjD0MnK4ngjaJYeOy4q0OD
wV/Ua7ExHAMLf8INQN8DG4RYgRuDnlGDgHvGTtjA34ZSX/PUY58VAq1jsA16MGJZReSL8useYd+P
KYzWhouXgydX4hWvEqDNTyAr/SqWYcZkWINQ2oKjl+xn5r6uu9MlFxYg3siVhs/0cQv2vfb6136v
x5oJtCv7HD0A9bPxQSKjdp6ysGtNl60PkTRw5704xmltUu+QwLGNNfAfLyN+tW6eJFPXZXxwQWNx
k7t3jXPeGjeubPos0uzHK9uqJJmHBJ1NJKsQ7Vsal+Bta5gMQQ+UqmMOJqBVTGgiRXhM+JVhQbGH
x2Eghm3uwPJN46YOwrv4KgrmiwEh/MEA9Su1r6373MpPkiKcIhcCbd3BpnHXnFdCkbIXHU0Y4TZo
WMeFsGc/jwMFiGCE9gzNlY+lGNAKSRv82OXbMHsS1H1vnz1pQu8JF0rFsusV75zcWp8XmUEjD6gJ
z8A0g3JZuDRoTsZ7HdKWP5PtNZp1MPS0c1I61UYymurMD3epo2B/i26PKJ+/jEDu/uXRIUchsghI
b0fLCYQaA2f0cewuwsbln4AUvi+v6nb7gFcVznC3Y768fOPrmYROIR+YorwjLQuULuEGIQIcRuVv
AJo+BSRmj+qX1bJ3RmHlJ8ltdZL6Ly9kdRseXtlHtEkbvudIrUBx7yikSqIxwk+v+2cglN1uWrUU
AJNfEYTcDM5KjQT3/1nsnw1EdgWnq0O+CA6nD7/JDOHzhoxmQohckzzzjrKymQ4C5A1oWU/MJlgj
A8g9jZdjI9dv1uAnHT3dBiMB/FImF+YYIm9Bj0fd+nBhM8HN4LR1QjyZk3Q3T5vL+dnMPTsU4X4R
L4P6wEaFxEGzQE0UCh+WrJEAE08V9nIu7sfelRERMtPUMoEWyLlJ+pp2XRxQaotPR/uFtcFbC309
jRTlRl5THNZvdlREEBUzsjbmNb+XsKIJyBQMD2QRwTF1wrrpD+6NRbkRoO/XI1JiKyg5zRJNRq5c
iTekAot+Bia7rWr/zfhstrHAGL83ZemPoOPs2dJx+4G3mMxXGBFtBhcI1M5Ph3j8BuTkmhY/s85z
TuqkqENQOFNAwa3AW8gd5QhiDEJpfYzVAC7B92oQG+iskQgYOgkrV/QtHX3yW1LevN1g7Z64Eret
jFqQonCw2lb8yRM/45w6V6HscSS8aCY8yrUySwXD5YaEUH69QfSFb7DVgJY7O1Egmr8jc15skRKX
t8uU/8JFtfLzpaf5JXN8MtNu1eCGNiAOgjLsJVP9rAnrrsRqPAx1dWUbSI71r71784fJMSFF9VtE
H2isrusI/MMmYoAsX7mJVnKJxsmU8/hyLBWKMZKhKXxF4SOXpgeB85uuyuEPsPP0r3pTgI3o5Mjk
aZsdPrsZj5IMAq3p+sBzQwvNlLA+CoQldlj/CfQdcPWG68Bc3BDnDwspyN9WS3U5WaIjUhs6vQgz
fCbNTRDKcrUekqBPrsrndj8hlyDBsiF6hPPmrPNIxKuGKIKm5aOT/0WHHgRtZCwffTid7vpilvPH
WL15oY/atCj7HW8Z7k1NfoxOaDNDZOxAyz6i1lIL7z3zbmZiXe8sWVP11/rgC95E7kcHSG/lmBLR
2rHL9AwvINsMJXYWfNKkKa6L/rfLJ7ylN9bnsRsMCGBbp2cgiMPb1+n/OP4Lglqhn/ABlPXQq8Ma
JF9Pp7qkL07L41Zz8IETlC/kpVongYwrCMkas9rYdKnVYQKQzfpAKZEvlo5bDFoSbqNjdGbKBjJc
eE44n4+PVn/hgr+bjq7Tr6nF1miXo4cU2nme3LesY/3Ukhj+HfvmoaaKaQ8h+avnqul1LNVhLjd8
cmEdQFXx8AvwD8dsxdlkqeOGEPxz7y2SLMAPMyx+x2rxrjDinPyp+WtFG5SILIjNTd4ZhxumU56i
Gh/Ec+ariMIypaKC5P79ihdVGAFc3rEb2t2F2lA4/OSBoDbLuxjbaJRLVmiOLJsa4LbnY77saN8D
UKEZqhw6YM8mlXK+s922A8NuKkbDtP2Q7YyUXG98vPfvLmaixmRAB4mrBF4ReRGtFiZV6NprJH3M
c3z94pSkt5rjATgv9JL5jqkTBfDpKXVyhZEj4LHxU+EnJYQumzD7oIApFDIXtk0kvHgprOuBcJw4
CpDaMQrVvs/1mmWIjcXa+YOFTwZbDz9zNzbjvvrJqzE6/4f5RZ1YMoQdL+8l6h6NojfNtrYKfKB9
dLsdayagd1CuFqi1sgun8ybzg+FqtNfrbYFib8AVkSnJUWiOf5aZGb0usEpLPWlldYpuJngQW8TZ
UEsRY3TrnV5O6ZPVbOlPpqV2APrqArel2MbkO3Oh5EKzrTA8vgaGUf4KhQxHqrEMAJGw1Ld0dtvx
VfKmjLIhN+nBWXQkW46tjMyp6H0lh5gTHAB2+L0yAlcC/l00djqqba3ihHXa0Vlb/Evt1JUhbZrg
rjqza0lSkpYzESLJRHmiG7CcDXvL83P1nNJ1nk7Z3ehis+yBiH9lx7NTWfWML894rKOyf1lLHl5P
iQBug0GicE2IHg+2pOcj5LjrXeVw5J1A0NuB1MQ+I8eIC4Ue33y6+d7D/JFSTpwLV/qTVhyFtSe/
uMMezBW09AejLW1hPwQ/bvEFzUVD7skTuZduD2uuYwOCvprBoElFmXy2v/4kub24FrX1qmhQ/eKm
lti4ykSadPME1tRwq87CSobRXL48FJcCxgRlAXfazbUEtZ94y2A4+E1RSNnK/JRcR5vRl18vWdFB
ln6p9GiZqoo7klbJ97VEMxeUfirnrYbzUikfcAzD7SHSsxYhqf0VWDAN2jZBMyTRnpl8UFmb2qyV
etWQ1+RCArpMArEdu9SgRejMspRYtD6wXgL+edKn4X1+w6bTowzbXj2AG6vgsI0JqxCzSj+9hU8e
Ojfz+jQybURhbe6SEjsC5fdFlUlZWTBNvPKOtiCP6QE4xnmGXI9KGK1fcSJGvRCgAA9ZJ82SV5HA
l+auSVT2zHhnyS+37yDmerelHY3FdoyXtn922M51dTgcwJUkNEHtLTZWheLAl32qNF+T0r85UyUt
vjVOPIdQesnwKRETq4cGZ6/TrKdvSyzqifsBxAsI48XEHLES9QqxZWMhtGaK52rSzJb/bbiBDqHT
NYb2cFRk3fc7peWoVg5ng6Cz2gZuQgTH2HfTXb12hfh9GmJQGWYZ6PfR2kwrmzg963YL2hmyCkz/
K0dvW3rlfjFpRUeYgwqapjNe+NmCAPq/tftEx4LtBhwTi7pI+fWM11veQicfLqjnnc/38jHpGdwJ
rATvEKYJyOYKDkOYduBgwkFpq4lNyy3fjV9yzDo17ypDMFFIMgyAJvCUd/KEs74S2Z5hO4lGUKw0
JgmEitoCUI94rl5jIxEZbzyA9UJZtiHdf7h/bvb1VFe9Phr0kF2C9uHLAbhF4n/St+VV05msVvOC
hEA8RQIsR0X3kKJlesHU2/JyQPXB4bcZ6Z9g1XTQcrs7VtIPajIWaUVi89wel/BR8ugLFnbnu9tm
K5RWC8doQtNUT40VDTFtUP1t7gS5liOhbRWonIUqnr/fyrgWyS3EEvTSUA+j0m519d0NOhqNi0fo
uSDEbDz2Do5jYYQXjUTQA58fZc57sohbEWcGn0h4Fka83E7/5KwRLE2/NKbI00edDLCexsbaP0F9
LzuRqV8WbHV9vKxmD8Ob9xfhbIRjMe7Faa+9in8T/5UtLa2LNX75qFavgl9Cmq3FP0JF8oJZpicf
fPGDyWrMcZ2rTzjiQnhitloFVJiSrJy4pCnb8yaer/ezpnvH8nwPIliC4LUZCsdeWytvQsY02SbB
/BOK2QSCD5/vcvVH3E3720t7ivc12zURYhWArRJa+tL7MkaKAnAwRbOim4gDMylFVpCTOQLvKrVG
Qvz1myCEH7bNA1wRvPGci5NKj4fJN01KjI3xkAlIoA64DLUEVI2za6UGvPV0HdvsUxDLM6UarHkS
TkL7mbehfc/V2HvBlzVrR+7QxEdhKljpU5SDryWtipWGQZJIwC6kSf43LOZVG1CRs2XnbB3jOdy3
vgE5Bxy/eh/ia4SvRNSSm0vJkEisqhHJ2vpud8fo81tCIEG1vesszXj+vslWuMfl5ulFfWrN9uPk
87qm1CW3jnBHPkgKArNlkpt1r7rFnxnVgTZ/4zmTWWXbvzTVIaPtigmlttapfl+VSc9Cg2xmYcRe
7GfKQYGubW7MnEIeytSLBZOs66QncTpCZ6lIZYs9Jcn+bSwHkmH0qzB+rVz8npoqBBoqRbeupfEg
DNnsnNvelqsN7LK/40VI9SXZCRBPu1AHhRfgrlS/b2XEeaIQrtpwFRPl70j/qkjQ4Z+y1H8idQyN
WcA92mEt8EeG7zR/yfNS7jgVDEcmicXz7X0hbti9LQWkbWN5yuNvWOkEtuVrMdbF/wcyQYo23Z0x
olAlEjz8kbLEmJ4fYqkYlVWE9raDmRTPZpXFZatEdCWlW1Gz5JcfV2QSzQ0m9AN7+dxG7J4LHrC9
k/WiI9BryYJ1hatriZUS0W+mtT2teAg9RWxG323DEmrUYETjSL7EM3uf/d+vOa3QfjDBewI5o5pg
772fPW5RpeKlXZAgdC2/K8JGvC9Bpipias9GrxevHKZ+UuANUknkPkG6R7ycQlBVWI2an43g0UQU
R4pWDRJNalI93nyyUGsRaYE1Ri1vrNAhWP/2PD/x/cxykO1+An1Nl7sEcmlmR04FN3NAuK2LVj1e
2UKyqP8c4SamCEBoeD5Eb6Fr0JarHRxeNP1PiGZeV/W7U0pxqgaMhKFPuDrd3Bst2FSvjAr234WM
X+/esVozcDVKipx3gMWd4soWSr5Y/7h1eYmYDjXZ00D6npyngoGRiUovvsVt6EpQujpaTPZfY8LV
ZBXQ9yaiKcFX+jNEZGTj6/qMA8ev90XaJSA8rOzvqIOc/6WZBcDepv6XUA+n0a85tEy1boEnsHjq
HicSEDoF0EC3NnRbJE0zoe34GI+xq+NM0udPURvmd7xUNLYVVuBC1r/YbMHNzzJhK2nvQSddgf4v
OVYJ9WmpWWw25Zqh8LGYS6vWf6j6THlWjb9rghnXcz86JNuL8jFGsiAsj3xW7IKjg7L364YxB9N9
07yyGwu7Uo0SE3ZwoHttSpTJWO1zpMDS7zuu7GV8ls71oQgH781utHhX73hgWtz/UDcgKEqORPKB
RDdjQAzC+h2KyERtRCLbuwwbN4ugWwHbzCKf/ZyDwB4EAZ9AkECKghcp0Ye3ZeD5sxgJq5UhETYb
5i3IKFhAaGG6TN8d4OI7HsVMsA7FZ51I/eRu/NoDGqv3LkD0iH3BvEtG/IjxH8pOTMQxyUqkQuqT
AWdQoR/4UE5hX8SSw3Xv2LFFVOOAriI5J7W6AXjOFUvo00KKG8+HLgYwyOFrx0fY6m0g5sCri5Em
2IfN2361MjJF/gt3zoL6FJ3y+qua/btSDaHRmPIFklTAthgHliCVFKEzx2WFSIWCfNJR6r9Zr44d
HGbQPsiScFxAlSIIVy4vw+hDqA868Na0PzlVyhUTtMy3HsciCl6ZDxoPm41chmUFW+eaB8uWQXc8
pbKPU1yIuGp4HpEN3XIe+8tlVc1M2XmRRMU9tOVet5CKRVemKMYvhd/6OxMyXHRSs/McQh+M32sw
oROKx5sTv9HoqNkDPNfi4yImBEm/yEkSWaDTuLQOCzToF1P3FrUVGWEfFY2ZZKJTRdvXxfPAiZo5
8u0CGxGUj6Q3aYMMp2jZwM2kArFheeaH07bEE3QNpoUaQujoArlGVpYuZSi3yTTLhGYMarETdsbQ
m/Y/LDtEfkIQkjIXcwXnzMygDqqFK/ea+S2hTTBoXR6g5BqdFdZmVOkxkeYoAUjTM8QlDZk9LJMd
59+HkvyPJcusXpxSQLVwPHzoe4ioVt3iuLSi2nRFdB8Zm+IokXjKnRlR+wrnpfz9G0rpt2FXz24V
54m3prYRe08McyoV/dflPZec51v4TKtL49UULZzESZPT0LGYUXB5T4byAEml8KMixwriP0uWoiiv
qqdkmZHd/AGbovmHBRhv4L4ey+0jN3QC9QnM6Lo6S0SaZpUykM+TE89fJvqgTlYQqoE3qxKQCjuA
VV1VxIdRnbTn9qRPdbnBmmolkVCLBuB4TAdL/onV3m6EvaGgq1sp9bI80jorPuNNxy2vfiIndHxJ
62SDIsHU5/ve41mi/OXutd4s/fyCVKeZS9QRFOc5Diw2zWGG+GGRAsbZnNMezz52HZcScePzJZPO
5p2P6O2qP+FaoEKLI09wHu2fOkQQ0uSfVKu5qlV0mkdiuAzOIew+s9FozQImetBuRu2fGmnzWaJo
tq/B0biFWL4FZsbAyHto4UOhSHZZWcxdTfquylVrQ2uBhjefrkUptmXvlrJZ7aZr92e9xLypeKeQ
Lh7PXKdmi+V2UdPZqkO9x31uJSD5Qei3h1Aex2BQBcPPpNU6Mk/JJDVrRT1Nry4VM6nSF0tpa/FA
jjAbKPPO4VVntxIc8uLTb/IdgVC0Fe4TRzrYxG+cdtvFYdmY8tvCCSSpjbBYZkJog6mnSGD3sQOX
a/oZit1Uby5AiIcY7USRvQy+Lnany8tq3PRcaR+1hlluuDhSwgDJ9WQ7YydehLD6Q4lvYIIMdYm6
CYXFWibMIGyorf7TJm5nQhB/S2aK/E1UU7aXMSODAct1ZKDn+NJXbTnI8oxm6vaKXP/Lyr1e2o6+
HAi13CpqeQPrhJGHXd3SLc9PUd/FzSvxYzYgJwxUc0gN3niZLhHBA4gtwVM03MaT6ZnfvTITjTes
rlpujJpdJfZQkSgUhAk/Ze+u7ot+b6+oFKdIPxg9q1cEVIXBcOqStNWQXgbLacmw7OGwB8ULNp7y
mjhxIgpRiKOejBKYPn4QLEFB5dg5mc8jTs9XnKPIvapN6b5d8Evlge4zCCZCvW0be92y9tlUzcgD
FP9aF0plg6LG2FGnTXotKuJR4JcB45TAyslE3x8uiBXVLGycOWP7sU7yPNraJ4tPKbknTO9sFfpX
IswuEQqFh0k7SLHHhhsOwi4HN6ai/NIfdDFT0C4+qo5uABKd3rDPkWCvZSY6TM+YJ6BRwoT32eBV
wC4ddD7pFrJp0iRvzEo+S48hwa9L6vR7yp6z43tmUTZ/fNwzlKmBTPr5BTmenc/mO/hS8J1sByIM
m5k5lyAVZ213GuwSPwmqtmmUbhIEnm17C9NVIGX4m9OzG5LYm8NbEo/Hf+St6tkAKPPBTQ3zm8hw
QqqkhzFv0CE7dr0OKFr3DlLPcgS67wpZMcKOAbTuj4LB5K8NfEcRALocKCA1zhw7IswC6AQ2iZ1o
vO5crBFZ+2YqGiX1feCyk0yJC+8fzKzszDmpoZAi17/MZ1h6VC+Z8tITfqAb2QPZRxGz6wKqM0Dz
JLJ+FB/4OJmvTwLedFQ8gwpUKYrlDBuMaYWEbxAjRnZ4FI3QPewyKNtDiiKPyt16qAuA3BLlkBww
dQ0BCzrskQGwBqsYXFiuG2SvKeUE7XCu+zrS0X3VD5CC7tov87dggHYM0G6TrjmlYWVJgnLbVR1Y
A7mkNYJVNLhqZKyHXCz4yj4cxE0xUgdMuOH3d0LfNSWuFiFSgUAJnioWIPgc4XlR0QGb51CQY9o0
uj9bTQ7aiscVf4DyUAAj1MROp4BGjxap9KILLDDRoDMwMzrlviAmunygUR4qrdTXW4F0QHtwT23e
mRGhUkcOMRszzxcOCgee04qES/AMK9hyv/bSOJ1xcrzpzEiZRsCaodTdk1Q4dUTSiMgzJAbb6giV
+xHEYshJgb9N7B6/HY6M8mVTkDL2RZwXLmtchsQbVC8n9ePRrgWECCclegtlMdRqiTQvfkd7oT0G
e7HMdTxINQiianrWF2Mm3NCar3UpblnIU/Ik3nhvvh1mZO1yp/mG8Xd2nNCRSBANKjgBrL2Njh/1
cp27Wxd2cnIlGShEO0T8jj7W5RP3mZxG6Gm1i9RNk6rotjVVUFO4/uvbLiuPsf2RHq+dYRI8qOn4
295miMKAHK+/9GYCQgTk0d5DG2sXpM81uS3h2cDL5G+/sLseiE6PXfKX63B7fzyaOaiJwvLRAWT5
3ZmmoZHoficVb/w0bxV+I8ZovFd/A3mfjy4e0ocnKL6/c5XAHFYESfSiXLIbqVInTivHsN/xjjWt
51tolIDn58K9LmegNx7selW1ib5LZjmtMubGkd2qxl2aWGFFfwfUPUoYAFm/DTpLLr79tRnRN7Ci
e3AGheKpTaykNS7HFZyPrQ+xRgaTGN4f9HA/UWWvJ8spsXvhZBzAxZ5lX8LUgTypoufIGOojRh9m
m9f5gBPBDZL1Nsw7FfC8SOMBZx1/qW3zKTpwiOSUltD8Mkdq/lMRxZhL5lhflRV4YkwTSRFGYkyR
IhxiS3/Do1+UsmulbviZq3Ys8YXTuU9LUfY5+UvkSDO3HRiNtFM0gFoOzdDkFJi3RCLoTi7F4y2h
7dfgw40xOh3RQ2bxxQYm40S0jrWgisTtE0eykRTN2XGXhz8k4EWUfy6O+Zu2V6fiIVJhUzi2R9DO
Do764IHyk0k8RcnHU1GpzMEMscZgESy+iDLetVrluAwflLC7NU3rZq8JhQzCBiPnHokzInwRHv1J
ayHGb6CayGuBTGeXQ0m1OFrflyJRrUvX+cqIEvGVRZI8okxh2tWB0IGPPSLOOxyYVpHxPrvfqgv1
DyzTumLDdGN/u9cJ9AWb73B3kFpinqaCENJevSwapsyz2LYkqLyBD/TTpGRKD3EG4yZBSTwudbmH
4xXYkx04t8HuZSn83AGIVrUEZ4aOc3/TwXPlc9fGXvG7tm41PO+unzRJ1UcWeGMZQtmj9PzkFHlP
Sbyo5fQjKN9VEWufY9gYfocFY0io9Sa1gt8wGLjqcgXjewgbdkeLtjqYhJ/VHNy/Fn5bvXjBvhNh
RN/q3m6gvJ/DJLU6lr7E0xarTfw9Ri0clY2xPrHzqcGpsSybQ7UWZkLrVS13v1de20nPQSP4QCGf
n19g9fd9bId3cf3qLFVU4KQPMs2U2vJKxuWuELd2AwPTssVtbHL3Kibo3Hd2gWag4YXBJ+Fb24eG
ulVjWSVqoEgS98lNoSMRsSm81d7yYC3LYGBqF8ECVKVQCZjRLWl5kszYDRoZ5jxTelsDmkVZ2Zm9
eZedaGSv67aQ4yDuWKQwK1NfEQsV4hnntpjKAeau6MczHuh+avNrF8Yd1NBc8A5EEDTK7zvU8srH
xUhiW9NQPuccChctoSzVZY9luls0TGj+QbEch5ENOFzHUI9yMWIb4MhqwO6z3TRK4/W/fSYMTyTq
STJT9EuRdjrIXWMaXKPC8MxaWRQjB+rEuVfx9p6W96g5E5ke+nLu7yA38LNZ2EWgJAnkJl8o00t4
marO/75hygwZpBu7JzbPi9RNUbRk8w0KRhI2cDXYqqGN8rWyHBJ7oS8FS+EoeTjvr2IKwbGwQd2v
r3k2P8CaAvfji1m21phNPAY9v9ATFQhtuoHqMEpTKNgZJ1pNtFFD01cL1r7YXWgVDX7n1ePkpyjD
lnmNzabm/zhEzo/z8xqsjfHk4I6eOmNLDIYaOqmyoY6bmvZXDA5gy9X2fDON8hRo91Fz0tJaFp73
/7XvCH4yxxhBc/CE39facO5MiBglO4ThbWNGdi6AcgADDTY/tiZAXeLFTVQz/5Y1II5x9TGSv44P
lXOdmr+/DnAhXHJTfFbM3tru2KdL+3h95sKTOIDq7A7GIs6vvrz/O5t4cLI5hx7Op3rXifJITTWj
yWVl4pYhRVJ6pqiRwSwHhDqlmVQU+C7On+26HK1Xfu72oMIMRZiIx5YiMHwgvM/5hkxT2XtbhPVT
B3SPYlmFhp33e57a+Dw/2Hlqh5Z1zFKA8jCbklLLR08Y3NkTuIoBDl4zspTPkujajF8UOBxObdeH
BxYl69pr1ML8O/yGJlAF0QUw2BZLihRT+Ck4Uj2+MVpGbmHLg22t3eycuthNyv/JAjdpfIG+KJ8i
EE/k5DxczcWkDmzA5Ywb0Re3pV6wEY9A6oeDl6DcvpYJGf8w5cnh5SjhS0m/RAXjaJPYsNqiOZzh
BkLmUKfKVmI7UwhkUkxjpAkxWZZwgcsfqD7kZoCOC99er0IpMXCF4cIkQ2uTSNsGOy8r+O0MNL2b
aPlSitCfJd36lAMZTGX0anGq3ZOJ+/Q+g1iLiwLqCiZuHuGTKA86gF3+QDqPK9cXoOUOTzKRs9Kb
Xt0q8oTjKBfO9DkEUrLmZcBzgg5CJxcOE8FGxq5j0si0Uguj+AyuL7uxGCzpLDdaQNJN9stUlXFt
1ipqRvUQI5tTVpqPjwAX9Ep3Bwvn4ig/kSkaMP945xhAqCE50r3DxLe9SVYs1WVl8KpV5BPo+igz
rrEjlMWVMIQTFcMrAcAWR46Vy+ZG0dtMnM7Mrl2tXhNBADtPwuHqfE6UtjJGOgZ793GQmp/qDgve
QSGPG5KmNybjb7Pq6Qecerjdz3TIO2dNULSzM8OZJ5UUsNWol5kWKgsU9cgOebyQyKtAYAB8xCaF
cvQ1YzO3tVHsKUWaJso0GAhc9onwwhMOZOANJCCGu0oYCJ3uNu31RZyFYQsCDAjfMDvKaY1UIOJg
CMtSj9aXor10xeHX7356BqwJcvCYiaG40Xme2ffcLbP7LkbH05QlY9hT3nW17hnyr3BmmJkNM6pH
UUgK5z57vQ5VlR0sln6ma6cpmY8acEnbyzOV7hRlkBrHzB1LAiDdfUtiskF7+JvnSCsJjTXDFxPn
SmJWj+YcEHFJiIWqlrf8Ys1noSEjjSi+xFosLN7vmb1ZQsfDsognh2cJLKu0i67kpDwvDCTrsYgQ
/tQ80peukr5M8XIbWLp+IMdNBg1IpmrRmsv33lmwjQ4SB2+ROaIBe5kSlFAS6IHL/b8C/0rLphfx
9qsnzp49TIysTcUbEhq8msp89CXQopGE5/KbIy6ntSEUiFTw8+pGIVKPcG7wOWaC2FZHm/gLDDkj
LgGhcggnx8yN4RJeSCBgakhlXc3sd63gHxQ7Re1Wgww/EhcF8jek9yE1toLgFoTdMQHDjnwxoHrl
wxB9jhPP5kgrapra0u48TwS2lx/4OH/Bl1m3w8Rsy5Hh9oRcTK4cvOf7JfMwlR0LK3mhM0SMQMI4
ilEK5eaKdNz43hp1EsTD3lKUg82Pep1gdTJFYOTw5JhmaNvLDzg26BMSy0EJKZNEH0moayGbEiQ7
lqWoyAsQpFiouyqLNpSEJ6kyqk5eYj18Y1bPtrNcLuhAP59AaVCaRyLyB25HLQPPHTNYXGKb+a9M
vqlE7L5uv8/0dGT9yYeoQbS5Y5c3YIdjxgmC/IsZqJJtL5YWgNnlcCd8apKqy1jV2Urx3uBgPO8W
ddRv+fcC8m9m1q+MVTg0HO4WlNYg8RdP3hxa6HCzU8Bdm7BcQmXtKxoi1fDOv1uKIw64dxQ+zlag
65YI7Sf04qqlxMMzsUxGdHdQ96AwIfD4EudUNyUzz5uKU7PjmZNIUeNfDe569yfrvorrYi0kV7KL
Gt/VdmoT9LRNKa4piqoycxlqVrIFzNUmjWm3sxDLgKfZUCiKaUZ/W7uQTBPA+jRuE/mYoTAryUku
9LIH0aKQeGA9Fk9RfWgbgQGKYAMIACqMwJ+UL0sf/80qxy5CZLxZhiLS1F9bFLXfJWs6mtU2GX+x
EXbtPfyN1aR5u5C4bEqq0NWE7iLpTFsDX2FF5SbvFqxKZS14SFyRTHAaPpIrkIvkFi0/TpNrz9Z5
SpaDVpAUt77mL9CRWqNmcxcBAAXgPgUpM/V8XWUHrsOsuhwhY3gUolb1KZ6cq64vT++vnTpctaic
IZvFDhntdjzShZx5jQ57756cgmpJsLQ1+KiBPEEO2BB4qfO/t+iSRWaUEfKoGoa+Yu+b/BUxj155
G3iy1c7unQbY473ndboI84ms0oibv99WAoscZieT7svvr6IauWT1ET9o1EadYsR9XQ/YM+2d+NYP
UGxZv9315DqCblghXiTHyiJYzH5werWL3gNBEcuw2fF5iItdSEamtdvmgOhm7LfMXTMDHH05hNC/
X8SbWwKu+rhLwaOk0eU7OK2Lsoo9XAPhk1C64ZsEt1yFi/F/+6u5Dw7nH6O3XxaC/81K/Wzn+GSA
QftQ2ZJqOyoE8WvnzSbe2AAoEhgSuPqsH+TmdI12eGmQBbaN5phlC3uKLITeT2HZ0Mob8GVAawuA
UJI/rFIvWNyA9zDLYkuqClJKNdQRhBKKJ5pIgzUdd9dlKGPuRx2Ga++RsHTP4NnXBXHVqByo6ISs
FaFKL9B+lmQ1kGpLYCTazfI6GnNT6PPrNqZgMqOFeNrm+86ZlKthJqlBZdVj/0j1ZW+plmr496Dn
6fn0LYm1llkm0Vp8X0ZH6TnpnZXCAo99QmIQddFp6NfaikE4w/b7dv8gUrXBd3tLXcCWcCt7o3Xk
Nr6mnq7jwvpQfuSOyuB1xrjGs5BeaoGq81bEKxWCTBnhbX/2HN2Qbo0ifjyYP1JNwgeEYMPEwfyw
wCcgNHxEL9VeKyFuEbOkxFNtBIlFQ/VDbXfxErYMYUzb+txJ4VvUwJOFYTmYUk080BzoYfNWikB1
L5vVDeDngmM7n7EZGEgYpgng9MccVfXaoNYpuRq+UnZcjx4YGn5gA/73GipNB9bSvzfnwACR58b5
L5vJJbVAGxqIyuo58/V/y3jXMwi2tkD0FCP/A9LgKnQ1zbBP3Xx3dN23rXhchx1pGolDSboqmo/l
/LgSgdTEpAj//hCcDH0ILGgt/wNOHKpLOhz8vjWHy6MSTu+67bihilnfv4vxYBCM8SQZGBOkNLu4
FjqNHlGibs4pxsHwNbbc2BLfrHE2bHqC2MHw9eCxQJo9V/HXAdGEtZMTCTieQqUv7WcEkN/qEcIl
FxJla9p6EWl/cNRmRQp71Sl+cYhMfFdEukXYCyK1LKmH8dotQ9s7/69MZcnzzghrdA4RMM2yCVXc
KiqrIFphJ508KFQa9mpHEyVVR9otphE9GoWZXyrxh/79LK6d/KQGfcLKOL2Pod55P4pRXdpMWDB/
JnvJf1a27gXIR9MFe3VMEdkzbKJyES3cycc2Rc5W/O7Y87K8laCzIS0TQPJlRBqbByzhKSTI+Bzu
KRYuYmpL8+aL7qV6/m25pc/MtBIkXLSsDdY0gEy+34IQCEgD3rsdIQYZnOXJ69LTnsQs9fUCF2+h
vdNn43LTptxRxRbotICJtRcnLGX6z2fCO0G2HxdRWK4OvoBVwuOWwULitXNoykU5PKztd2xlCKbf
oXO7GnKUBQvyzdW4b2D0dp3qanY81u696Uqzq5FaEJLvbjppdXW+GG7t7HzZ8YvrUbePh/edcA7L
eWm5BJypPOJtYl7b6Dm1gSrfueeaNGBPkTE49JhCVUMD/hrynjn0OjEXdoFkiZNSIs549cduwj5r
NLTYYSI5zBgWyEwxBkDeLDR2EmKSgBfi91wNUWI4LhsZoOsFYPkmxjpXOwbiVbrVNAz9QyS7Q8EL
C4i0O7q1RRKOBTRc7IXPYU2Ml1xefr6sgRlQ2wP08kGHoqI6TBagdRGc0qu+Btn1fUy/RiDk9kwi
GcbyQLgD+wqKPO5wz5yZHC/ALnz+fTQFX8Oq7n3cfdB9PEdgszss88d+XezbbqyiXKAblZb4mAtN
UOHLooBIQHAHCJHMB8yxqXhzfyZ4f8DJog5ANMUdyKTU8qWoQQZFaDt7nJQDV+YFpVlccACNXGKp
8dyyLRd5BZTPikcC77teaPXd8PYfh7S3gnXBHSgK/R1jL45D15q2hItwGlojj8DhicDXH6RtmDE3
rg4FGe/lKMC7knTiOdg1A+2nini3SoWUc1R/m1wQ7YdZSY9IFCXgxakyAcvOomj2u0SRBmxKUt2k
pQ/sLgrkxhsK7yPPL7wVxU+qdINA3lyZuF5f0JllfVWcizzu7fS9rK/a25VRbz8iC4Wkvh0kyF6Z
f8LP4KduuyFO3VfUAX9xpcQAUK1brPftnP9xKs1wdmHYjK75XPaNJggPSL9ILmL/zdwnDprfrDik
fr5r4Gx5fV+ytgdFJCnkWD2FbaHjSR059ED1MpaHsQhps/Nfws3xvZ/MudtGussM6eCeqqpZ1flK
WF5c2mggY4R+gW5vngoj9dsSX/+3Mg7+kPQKIGCZQjPFeomAr2FbKSiWN0VWEVAl6PZG/JdLloq6
Ku6HkzfHeA2cWLWogvK9uN9PYzeXMIRpCkX1b7nkIwB2hF9+ZjlbL+3SecgBHSKVuJCOI55u/hsM
YmYbdgr7H3opP9XzpGPX0k7Cg0deHCb6QtBnlFDQLFf+/ajCAhUaw4f49bhbnfSLkPZ6NNdyADUX
ly/EtLG9R6OdhHjh4GQX72TIa95wsbOwzSdEfvSYmsFPHnI0PCyq8h3rPdaXwi7UnWzzUiLNYoie
/KXbB+LamDu970HLi2bjjhhciXRVmHBmfaC0rQesz8UBUDq2Yvd8tfguHv9EhWTU9PpP5wFeTE7C
eXCqGhurpvOyQwfmH24DrL0zSEN9ZQB8pj0s8gCnHmd5/eiea0kBqXDYxQ/3lRiN/qciKr3frRR/
IIrboJNLLZVDey4QbXqhcYde9DI90Nmt/G3ehUgdujYD7lYybxdll/YMhJTGU7yTbdODl6v3FRPb
JuLjREsuNrk6Bjuy9J/fU503BU8wx1uwJQgj/VoedsCM2Vz5at2jI4cOjeIqcnXiexKjEYGCLeZO
FQFSw8IHXsnIbv/YWV/gK8bhngYoLD6YRTnc/4RZ6ykXRug+3NO0s2SZAPLQATFceMcwKW/MRV5y
cqsck36zw+3x9Maoc4bzxe++acb9NUsOz/Hr9tovp4cX2qNxhFT5wjcSUCmLl/NY4I80da57pEyB
k+O6Dl1j0ipKma1XW6VMi1mbYdYROartdkG3PTH6d9nOQaqlfud7uCmWHycWs+d3P+6tb+BcFCNC
jsPrZrTvW0uO4OsZxADPOXKgmIsnrljDm3b5HunXB3EGeP2eE99i+Ydeu5SdkSz2bgFMUbRr+51P
gf/37mKwHWKZdLrkoQfB0a/aoI1PmSq358NAgbU233In2EgNJ/PfIHPN+Y55FOc9V76C+UWsPM+0
qRr+an0EIdCqJmLKVkx58sG6oVghOiA8+Nvu/D2vbdReGgArCzJKqP3Z6F3xeOWT3Pafy5BZuu3m
gKACcyfgLwXbxOLhpZuOKhDfMpkdWqTdW9UAONlqPwuFFZRfAGSOgxelZltRSPF3VpF9rrp1jkvv
/lgABaxc5jNEegiGX4z423y9jDju1VRBWReDdjHVU2Ws+4/wfJB13QJWzRuF9yDH/Iu+ezCZp1F5
DwQi/M3IvvLyeCrn6xFOSd4d6HZ7aPM4LVI7S5B0918+bWodArkvGSwvjoNuqWI2wNCcZ74a0K93
+pa1DHOOpXVR/CqpkQc5AxmxETxevRRaeDS6yyaH8GMHFsIrwf1+RSU6Qu86c0Xk8Oofda4nb09P
ebJcoNAqU9Ifnr26ed7YQM+2ZzXNB1Zgw4l1fF4JvsRyTK+hY4AS4S5aEbJH+MO2CvwYw8iODo06
u6o+65kLY3Ms7r0C3euwZqZCVY3Ee3GnjVbsUhxTmZ5QvX6Xg1/ojLK9Uznts44rMo5i8xneXwT0
WW8O/dvkLb0NUc1NAvSdbrGYqwsH5X5MsWOJECgkE6LJRAi2wz41wynvfln0Z93KD3SAiXAkUr/Z
cPPyhT6ni2FbPO/uorQ1qD6jBiuoGVY6typkGhBPUZqMJEMCBlkvjojba0O69JHSOiQlGka9nVps
IBwt2uyNLghdy/zQKGeBlnTJ/ik7aRsm4lP6J5oICesLzoDr2nVTX8TT3+Ci66sewQCqp6+TMjVd
tSTbqo+F2O07N/eKxs/y9swl3lo7zweqtrlvsk9b8qQHWk0cb+Ibl9cFbXe7chH5k0yqMd9MT5yb
l2qXIOxNhf5C6UjmhiVpOJnuEMkyLIPZOD18NCvnFDqjgHtBADN/2phP65UJzz9stuxeRSY6vlk3
3+Tdv9sNEkrH1J+20c7kVv75r8Mf3LTLI3B3z4gzac2wSdqQATUg7vj6EIJWQiAH4Itv4X50ypdM
7zsUDuVqdB8ZKKplWJx6BDdadqeudwGlNhP2lrWcaHyDApDHox/aY7sko61EoGKWEM+lpEYXzJ4n
jDQ6ui4gvmkLCx/yfn1NH/rRMwdfbtAb7hG/wmhVw50y1S2Vo39/k/KxMsyNdClVsKQf9Wq+JWbE
FpAzFkQeuoGBX7SE/RJ99m55xpnYmfjyx7VQKIaqsgwvyNhmheNHIxq3S0/d/dksYGgLNrE9by1s
3HuSyhzO7shzpPkSZxpYrSV0e5ZXDzM72DLl1QroZBFN0CBJaq36Ivf6NlC4RWAiC4ILgcIyLcB7
EsRcdZdV6ay32jaywF2pu/2EOHVi4wCmfFOCK1oYoegytDfTQ+PiBoIwRbrHrIwU4gq0Y45/BW7F
C4VDy8IIXRf5kZVlxZMqa6QdUXGDMkgi1l5igAEOzvUdCAS5IoFTcy5gFZK3UbtfqPqTTXHaM7Kk
klgh0nQuUdUcp2kPZ4MoIMSMPmqBCfbgl8MsffYs1Va+aexmPIkFIne1xT4klGuYRFWg6UIguYEl
xEW0UVhbg95hgWbdonIGCTLEzQar584YRsrD5rPsGeUY+2ORCxpJeSTnCGZh8dwP28If6H6J8cIQ
SnK+uikbAa3l6dQ0+nqinf4muXV3D9aCHTXp15B2gkBdnUaAbHDJJLYEJ7UocSGE+E2PL9EQo1q0
iPj7INo1fgIKyVAHAaLKyQ7WpmTpSMDOPHSCDYcRj1Ydb3NoTVrvFhg51Lqx2tclYo9cKMCA3Xyz
cybNvjXyzV9h+h8kaZcCr2/ekbwqzhMS88algPN36fbzwlRAeHHTtK6fz8sakjtTFiSfN23raKgQ
0SlfXsoZgVTFKMYt19OHTGioP1oP9Ow2GWOXUy6HijyGIMfRtJ8MDge7uYVioNA747KnzmbLNryr
k6xDURXmSovfq61mIZdtThd9xu2t867Y9QQ1ZAn4TQQB84CJqktI5Z7ecu8bgITb05MFlh2pUJWO
nvJnLNDgLqwMhKgdthz8JTMwQde1/XIyDkl8k4yVJ6c+BRfV6X8IX6xdEa4qkuUn8CSQb8/MlA1C
UcJqtJO95ZdYkTFPXB2GO2XFoxLXsdgsubiK1D7CxIH1iHsxHM7PYJOV5FgDveKerRSbC9qcWAuV
J56Gli4xBUymfRX6aZBvvPaoOgdS+P/n+BfpSfikv01uuJksF5wfA4nAGvK0BF/NHZWSA0vGCFpB
Y5iZPgP6IbTzEeYXrCKBzyz2LyhNPwhYwTKfc4AL5YeWZkX1R6mhhFUlI0GUiJglNh522wkiIRIf
qNa5ZHNwk8hLebcO2lZwGX2z3GbeEiOkwk1icZQfBsmdyRKa8bvINxef4Vt0UqL5sRPZgZXl51YS
Vr31HzYEl4fnXnbKA9IBPuBtJmS5bdUF53qv5LYLyWdzqeTputLe1OqcJLoifjEJlehtBFIUtNxO
Ekwjm2RGVPUNqq9BsptqiVOV0JhTG/kUr8R/pRL43+B++WQkmWZ6Y7Dn217Xlp7uLh0MziOPcfeY
3NoVuDFbyqgoUuG53eoFHyd+envxbuOa6LoWu/NWmVu8tV96o3Aj5MglJg9ygwnb4vNffW1hLF5f
PgJBj5jwXS9nrdFHSRVUA2zzsg0zaI2syK9t/RUYkO6ef2PVlYy42d21PBW7xNj2w1dTJ0q0VN+f
oFsK5beXiWjnBdM7KXdMzHu/yvkzIETXt6fTvXx6s8qamoi/Sj+QlHH2ebWhCza4eT5G+153P1wg
F6GY0RcfhnxWuT0j4AlLiRpmGvoLNnJHg2XHA/SaEyRI0i1XaPaPyKp+iujRBtpb44Yjdlj3KNKx
BzZkQ6RdUXjejX+LWWLFRu418MC3sJe7Zegr1NjsSHZ9kOQrvxDCrKQBINPIl68blQVLw5d7Vmum
3EuTxyKCXdiUivhJTLe8TQVryG9T+BedPoGIfkYPtd/vSEiq2nLd8JUY7ttPdG76IZsQo/0fQyhe
heHpF2oT+hRa0g0pOoN9r0S8+Ul+08IsPxntVTDtnQoCcyDO9y/BE/H1pAZ8D6HVKvUkRggdDiRs
L9hK3qPEmUQgBzjyMvGFrMrm6XZyFnURxdwdS5mu9gUjVY1ZDWOo+qDctrF8dk5GV31Rvoh3IG3n
E/azqhb/H108kAGYuhYGHlNinn5+da+cCAbT0jEjXELi/ls0ISeYCGo2bRgVAdJzCRR/hFL328dW
OasMcAaAUIm84q+OArC5RhtJCG6LjhZHW6U1mthIQNqmjR4qgC1iVEkiFU7GCpTyPODoMmTUgMMT
sknxE/P66daXneZkaujWcOL5hrvZJWZrcDwf2fhEEHphqiycE9OX1VBlxj61wVF24zZvt9mG6OsX
naM4TcKBwBQADoJIJGDqvGaxFaKwlYgbHbsHpgvGK6F8KRd9wFYvMngx/EG8Zt5FBWkz75lz5jwz
u17I+lGlhGUWaEW3bigjXmn6U0vV1sbi4MAXpL8EsqGiFAYaM9E3c2fbwTtYXdRo5BLMMrf40Ay6
yv+HiSEN9eegCHGiVHHR6UkNwdovr++jmPi6ndgOEL2o/HL7/q30PrA50GcAHqGGm932qMq8KPoE
/rafinW1ua8NaftVWOjBtpfhM5L1JyQYmxHh8/w49KUJ72bL1pb5ifmx0/fVUblToSFYa7Sw7Sre
646A+d/t1gYENkde84bIv4Ji97/AFyTi/ODtOcN37zi8P9VGs9a0FamC1+BfY/cN7+TbrCAdBfz7
JKlx2x5qLXhy8V2J89tAPioOm/I4swTUFwWhj7r7ds0Hsadf4bNPNrM2kDvuZ3p1lkxx4ZpGezoV
oSqESPeS+jBndcyKSnLfUOW7/P/YpBnCIrHhGLPpqfDS9Xwu3KntqDAn7MKfDx1vd4C3UbB6zUkO
093kGv906RvAwl6DA3zKde8fzmzVfaeIOKD3JgpZmYCrkYty9vKU5Bn4TtPy7K/F7VUDEKPgSo+k
eE2gwO5Bqed+9b4szSpTEvP7/1C28uwDubpyRK5koPJWZxd6CAj3+EWJHy1NJpIpoA/MMdpWwHwG
xG5zD/ycRKTnEBIr8jl8OQBilLmuz1js2R0sawWtQF6yTavj0RQbmrXwC/CNUOfDb9E2mB1/Oyel
Adug+dJy/PfUfsxl+ufpneFAgr/bL2/2U/DA0M882pc9pDIDt8a0++nqsoT5bT0RyizuSAlZL96C
NsPlpgCWIfwBK+eLSmQjyDIPyfGp7rTLbxkvYINlLynGTKFFHcAGuXyis8NQEdk3TCH7pYO55wgL
PYllhjYiYhzMmTHnUYUluGGP0xuw/C2Bk1xGiqVO2l1LGUul/3Hzb1zMXd/oU7hWzfHerR8KoHbL
IiRuKoeTjXxY9f0UHAvVBkyCQE7BvGe45yrbrxBKipxhnpGPO9q8XC/88gGpe8m8YHUjxcGrrlSM
1l8TlyGbe95njTWLRc0wwQ6amHh0nEc7fUnTTxeeOOZGxomFumQ7S709ZLX9F60eJ7dNyQqs9Ndt
NWa9h1MAGTxfclteEQBvqqDM+lkxO/kp/E8TPg7rqJgBNgqoe2qCfjWwUcqISOz0l+h8gAI4WCmq
nXW4Zy4ZAgjA/A3eXBFAvP4lPHkl/u+qIDIohmUfjoJwmD3rLGcUdjpDXgHGGRMTWehcL2nEia+a
bvep2tiiFDPk312pkAriffdWUMFJUSdY0fIB58W/0aLedLjJGwM5jzfkX5zBZ4oEEW86v/JqDFo2
1zBEleI9V57eIcCavZPosaDzK37UG3Q1zNZDdTn5bonybIxZpUrdjvWuyit2/nNXAdsrCghNztXr
Em/iPo+/mjoC+j3w6rxOt4RZR9FupH/ZkEtCvsVr0tiJf1BnT082qcpx88SXLRsIwOAtkbdisp4n
4bAk+CPTScAecO+E7EWC6peqygixKX6TqytvRJb3Q52Kb4RWeNkcU+mXGvT3ZY6RLl8EZ+TRJVPK
wzAJpWD0hsYP4gP3j+Lx1xAWLxO2GUEjLNfRlmt7xnEvfJxigEnsw13OuxP6Bdn61s3sizJNyKJK
iU+1YWjTCBsYFNpBod3yDSGVtk4X5obQDm83BT4+D5T+EvkFiNncp7tlndnfSvbxcYsjSLrToqgK
jxd3yO5PCvscGBjymxOfWQtgkFb8LiEc0VtzWE6dJHF6ix6LtHqYh0Qm0K2eLCXrIOjIhPA/Llsp
EmjrvrVopMaVjXW6tOBpSi/icSkSXI3wbZPrWAheQ2Y0RTMXvnIeLVJxf0VW9l+oX42eAZ5eYyLE
n2QeSSF8xEcO4OzJ4ZVoTVV4lZWLvN37+BbVXnr4qVHIsjfeO7NHIokhnep3KSoCp4HfeZJlcGr4
FNNYst+OAxG3LBxmYYEzpsSwhmIUrIA8MflxNN3n83xMROfKZDNGibvxsXAq8o8kqi26dSdtKj8k
m6DxwdT1hjSfiMYJjSl5dWRNFd6FB0coyGJa9B+hTDO/CK+n920QUiZi8QW9crcoYgEfnFixnt2i
LFaR62mi6dtnsvQV6BkbMDFCT3GcM0ealcoGwAkERTHhVpBlPqlsbeL/m29WqgYODEPVNs9oy2Ja
yPE58yYS/+StfmaI4I7PMsxayZsbNRJA3dXoZsqUVmwC7yJKKJ9YIMLQKmGwImvAOt3sp85dUNIg
9jbl5LctJwe3N4Nd5E8wUjS5g4Qqrl6TYlhRa3fQU1XoUtMoKN60xJ0dFBXV8uHKd/Vo0HSMNat4
qENXHe15nqKXZk42Dv1mv9Xt20bcnPipff6rQ4FGt6lJnRdFGJpQfYWUUcnTRlUSu3jXVh0W1VBJ
+iWn7z3uNNTURtFblY8o8+vR2mBoQaXcoN06V+ovxR4BNU9sCTKEvLiZiGCE86PFYk98imppsNla
BFAWgDF3YjshqMZwQjbsaXmPxBxPOoPFKpWER6yPXulnxwCDt0AlOb8rrsauzMkChox6e93noJer
4HAD72+NuT4q7oft+6oejDSVRqkgryjwNzsNM3/q/7Xs3XfZ61xXZkQbXYoOgjE94Agh+BnSjDDU
sgDS/N5ys6xx2HJbfO8vO1vfV2HPU/BMqJGALk7bOiLutKiAvwxRLysh0A2rKTb2mGVUACB00NQX
8dbAXhSmD9B+e6JrSfe6jIkzkCB+EHukIPRggU4V2cjIp3i6fU7jx9d1RQ3toSsCq5wJmV629kFL
nFJ2t1mW2cpS5DNVYNNAINaU3sxuDifEf2w7AlMzIPz7pkXK/tf2myo8pvj618Es39/BvNMdsjVc
+ggHus7qVyc4qvQmSeB2Yk5zhv5yjHL71/UJ+iup/qRukyFY0560E5NYUbCwAb020rKYmSbnY9H1
3cujoGNgu9iewYA7wiVWpffZGJ6+NEZUn9cVKKC9OsnI+0lkuBWd1sOrTcb1Kp47IMTZHqPRT/go
y6KdCTneto82vuj1uz2nk2UsbDGyzY02ZvnB2hE5Nj/qjXuzRYZHvFTQhydbLjrYZliRV12PZCDz
T9eiEcrUL7H829KU4f2IiBXF/sn1cMuRk9XbaQq1YbIbL/yFc9NrxTM6jvw4nf2V571+LiuzjWeg
nbvmcB4vHUpTIXEnJpdlud/WFwE5rUqAAdxMwqlJp2T9x2/qzlzrGsDGlGsJ37XK6Hr1b9Run+Jl
JeoqM0GsPrYfFuu75r0L+14DFTUURGa67b6ZQsyphWHX8mos/aFoQycD2N2lP0LmWXva5UvV86qv
28vpD5Y2+6uZMwlmAb2vun611OXUPH+WQNek8jwbVob0mksX35vvGhN2YusyMAilNexa9obtNvNn
wEsqS0i93aDuGkYtSDLp1nm5Z5I9GiKRpg/Rg80zu9Rv0Yat7lF/7uotZPXka8RSr2p2Nd5U+W9i
ICWAJKC09ih0t0FVw6y7ony07cL+unvcIY901j0nrl4IONRQrt7BYJbZhRQWCdMxrw+8/1InxXSd
xwsSYszX0CF9uaHmkxSIdPrZYeOMUEuc9pN+Gu3HkyF6rzw5anAVEX0nDPfSlbC2MXsUXxAE2EbJ
Fvlscw+Izq4kVWrSnjALeAABpYLiMdWwsBc9kUAcqD4tT1uQ9nEX86vOzAoMCrV+c/578j4qVao9
EZdfAYzEmMfz7SoMA549GeRXKWeSmDicgXBpSLB/DX5pa7oWb8OVgs02Jf9q7tBxQP8BhCHaPArD
oYNi6cbInKdMx0MN9SA3qhP0R4tkuC8/crDQZoIZjlpKMpUmiuZXOeykA9xfvj3aUiLKMiZQmSTF
/Akau26I6PGNZ3QVBK3Rd7H2b9SpDC2MmsvRIL7iYu3lOsJgquR4kiNjxkgYT6BPlBVbfxjBWizG
Y6jb+MDk7/RHJ2tO+W0OXwi4HG0gGQDVrPMDYkO3yRL6aZ2EorHgok7cWeC7JudHKlz7hNl2M5MF
HZ7oQmX6c/kcqkB58xkRIkRyIR5p9F7imjNUNZc+nBg8eh+cQXxp7L+XtmtGfI31ONYXA/BjX4Mf
FIeDYPsUe21YI1mhw12rCLug3qDjrU77cLzjJAO3ajS0pBIoG4PsDVYdKWVQ/YygYx00X+AWxF7g
/SIAVUGOdmqijjIqjAa6O/Byj1ANoc64KAyDljVz+JKrthPCTWTIiyC5iiiInGdkxzGH9dMN4FsD
myZlQ8ZoGZPNiA2P4MhfSN5w1r1gSckNtW74sh361dOQdAFrCI27UWWBkxDHR3g3DnTSU4rqStNw
GG06tWza+RUf0aR7yOAMHd0B82OVGA1RNK1I+dTVZDW3VdV7jizMikehV6aadMRU2vyuRhe0xHmV
WLfjxzlx+1uPmXgAhfFr8fGKJnH+vRhMbIf+LuP7VankS3Yk0pBTHsnU/33XlJqFqrsNM7IbAs2r
2F4BVZJBTEURqOhEabl6BQxvgiNN8GxpNvdWMjC6S+aSanInAa3uk2MnA7Tgqsv8Z+LE1y+K8QMG
3VnrDkXWk+PRxcy3j+Ns9gng6QkVi3hwYUxjdgLLCuvKUKAtMUcZxiXubsAC9QdFpqUasQVcrqap
7Vow2YTn5Xe/YK2uVOVPskuDXJFwCCAPDMNazCGHbbX4SPONfRvvXp33pGPCj5Nc8WSri3yzeahb
qfv7yJiN0pyo+C3YXjnCmQJPi9ymo5ZMSPSv2ZVlTIppePpxQ5KrO8JrM/XlRlL/6BBAQyyGligV
IjpAClJKpzAbXTiSsbAwUcvaTy6A25QaGXS1DGPBqZweKbNpg/GuYMDA3CZleVg+pUT/DchlhfUl
KXRYZZUMT5bTeetoeX8qzHwQflM3imAJnxlGVWDxRtwZXZNJDfw+sI0pIO5thQ5NsKJF0wQh6YOw
xZZwfSNtWzYMuBiDxYQ6Ss93dD+ndemJA9VfMrI35UYtMm9e9vBdIA3oMsf/rHQyme6oZ80XfYsw
r3NACjUp+jERBfOWCeVRNKKufaklqOvLtCW/EoM57p+r0VPogQ1HS9E9WBGKvFBZiNLLqECYN1Le
5k5fO+Zv8c0rVNWJ3F0dtmUsX2CHj1NS9lqKn+gMt85UC0tzgBiHyqsuTcphjrFdnKT22rwBR6On
/a+33l2EVneSSJsNQxXnwhtmZD5x+okZym+6aGYWQRXqrv/Yg386IjnrqJTlHdBELhdXcLaAhli5
9XEHdhnUzBLwNpi9FccQGv4gmAlulkV8D4aOCklcjkokIVaP7trRm05tGi216uGxEaW3dj38Nw4E
CLsK3JrQRbSRxOzU2u3Hho4yLUV2blqfr01SWfq1KexRl/WXcti2cXhDsR+og3CernFtBdCBRscc
Z7xopgydJ6lxP83kxlaZDW1WEeK5wh77Zqb0bje6uX/rNYin6ZubpzgFrc0Y8WekBxvKg1nL9rZr
A6zgAGA+llWHR9h1eVC1urzJwqMX7/TYif6ynGWhpzCYe7PMloFT9NpZ53qJbooG+9hZYJcnKx0g
3wt6cuUPOSkIhhHrcgX5LCRQ1HbCiOprhiDHqAidyMid5xf2ybhyJzevMI9e9yoDcS8Vy22CPJ8O
7MyulCgycuLoTYO6zXDadl90R/y055ZG1kFXMfuq6RQU3yyq/3ZHV1f86NMjsXrI0bKT0Yabd63u
LqyUxDy6SAItlRi6vnE+oY/YnXHUK45Xey16W7+upklrC7NjDJXbHt99RC7umFoYOoZe2C+3nuGN
Creb0iZOMTnYM0mj3QYAEvll+ZK2ScBx3zNHbpEQShfXNEdQwiUK/QNFQCj+VrHXJNH97Tbq8t97
3AuNlV+T3Aq2HJBsFIh2cqku9k1nFNiTYX/B+kDXc1pcW/zBw+DZVX1DOhzwJlaNvE6wDsFpg/uJ
MBZA+VRHGIHlSuNki71z1C6B+qzTmSvtsHksjAQtaKyPQzssoykg+GfGIxiYidFPgORpoSuYz+MC
IA+LVZq17oa647dIHSbYAsf/PlqCFLTJgqPHY2oTqbFowF5IKl5IDwtRqwfrtJHZVkAUCEcXF9gQ
O0eLF0E0QVF2sBdCEgoc+a6kGAVgspYBVbOntEnLmLPvvcCrANNTtyIT0NivuQ8MIAyoVwqAH3BV
qWBgMVn0xWgpvhy3+fBwk48SClOBQZeB/OK629tXo6m0jcljcOUC22ff/tmhdLdkNgo8whWyS8RF
Dc83Ow27jCW+CyGxVtLxhYSd1WIwUIlcOFYMwOJF/6SW+qlSJwJr6A91ndUY8QoVbaF6uf6FcXPx
oqKY+rbGiGccGLb0qqPEDawJSajblbGE8ctBUSdR9h/F8uC0Fqz64O9br62XoB36vbrKO2DRNN+h
npxkxYRtA5VCrZHKCFdNtyxX+Ehg4MZPQzLjeJNB0PAYpkskFltL0YDrihSzw10uym8uG5dCTM0R
SjtLE+XzWFWFjnK2C0Z7ONZ6GO0lEWCkvn2NarjWPDPjxujC45nCtNYixKr6lHygVwkoiuC0ay8L
GXFG7YP8k02S6sR26hhDSjaO6QfUwERzV25+J8ozB61559+WmV2+2qbynFU8Ulp0gAGMod1ZlwG5
xyaEirlaPLetqDyk44yqRIqn6wa+4TLitMZJ9QxzozutgQNsZNBNo/wh0ATcK4C2dhDRT/8ojERl
jkTjc5Lkw56tL1BteHkhWt+9b0tbQMUeD0r7WhKMYRoszAiRFziaoEabAYFSnLQKzZYmdkrpwX+x
4vMjD1DfxQyKP/+h+RlUIt+jfN8DetSV6e11af7Efc6W5FlauVE5u3//aEilPD0uesccQU0OCK4S
u+coDHU6yOjGFYv6Ld3PuhD83MIG1kPFSRq+NwNQiBom09UhIeRgdE0k1q0ZI2y2ZiyxKN6KOKP0
TlodBDaGenqsFk0b1/eRpzukfiuXceE9TE5mY7lrX7MxRS00U5fxk8U0QYTLiIWQz9PoGhTiWTmk
ZD/PuiDgOSb7m42AQPfMRulXFD1G8XAwfmjTGg9TPAebNiauvoB6R+O5jP1DXZLJblnQz3Q8Kc4h
WQYZnZAtKJKdU0/wS0wivRKkd6QxMLaqBD+JNUkMJvF4q7tLPyvHtSOef/FsI9QGNvQG0140xF67
HuhQskaBq/8rYYGCjBC6KuYHaRSoIqFS86NMboWMbtX2v155p038/E732ForNeYP3ZAtXudDuOS8
t7xdsyzf1l9wyCTYpA25LsIllZ0b82HSDM4ZLCo4t5feIb5eUgJXEfMhbXJh0mqT/8N7X1tPzVHq
WWMrCUcFpJMRvva08QFUEBekXrmhVMCqjFl+/Ms7oCnCOP99KK10VgR416mwJ0b8NQzchQgPb26I
P1DwM+7auJXs3VE6s75xSmzi+i4mrfhG/pvNJNkkbhslsAPg8Ie5gLRh/4wtVq8lYYOzW0pDkHrL
1byvriiySIqH5OcoHkMVVTy0WemHqp4U9uMYDLy7kK/03rErQTKvoenYQy9/Bqx71RtcHiOoNQFn
J+lh5yniGfMxh/eTUAnZNU10xQC3PvneNdNq8sl+1QpuLj9cPkVylf/J0kmuLzDO9nztVOuoKIOE
QSiNIbsifx3gP93k0RVaiqGpkb7zwyesvRpZIRH+fB2HPmzAzqwKA5UuiniV6V+OdE4wBncWEBje
Zprb4aw+4pLv0a5dpv8KXBI1KQj+pJ/0Df4Jh0Strsxlu52Ji6E7lDKIoTgzRtvw+XqqVoggbg5/
h7zMS09n+MhO1ymPCmEdKGVgDMrNrr9kGp4kfJEqz1WXfgC/MmuYM72iOI4Ke8YJ/4G7NuRI7UnR
YDxkKSm/g1eR4v2wzr2/TFckgzJ6udcB1xPGiBoLX9WgGGl1tlOF+sForlK40eDdgRU6Z1w0rEjd
orcrX+VLP7dzRAlsIyoMrOm7mfcGLtp2RX5/z/bIvmM5BHIs7kFDqBxFW8fD0whc9CQNM3SbxNuS
5FGDPK4bPkCWbRiifwS8u3T9RzDlJOvssA0b7HQp2JoSGp4rGQIbOvELoWhANAv64jGlQ+ZvZx1N
cPNuTrLdA3HtnFplZ18khaSgc17sSoAmbqjJ+RRbbhigtmVKh8UY+A2J3hIWgfjwaAltj5AbvPOs
oMCWhm9s0RKJKWDVB/hUNwRSD6O9MKxxghPSBetlskgFeuEud4o6wLM3JWjxU0XjNAogKqd8Q0T1
1uVffadeIRUGRMXjmSybxEPPGYTiBPgZYKJ2gizrBNIM8de6dAxn41omz6+0O8cC5s97xd0n9WyZ
FudPJ9IP0z15nk0cEJLy2Kd2n3dwF/Q+1KadmZ5P9XWZg+CZf7pYvx0HBrZ1ZB6GjEvD/QXtc+IA
38DD1hVasFFQdVjFYxYGoFY5yEFh8lvczxdz4mj3ZjthrRTO/4nORpjjlGiZGEpA/9k7Aq+z6Qr1
RkMDClHuu0ZQtTct/M1iegUlIesxx8YNkYlMc0JzBVRM/Ex5OwsjOZAr0CjEL2Q6SUjDNGxr+8XR
GEJaWiNi7j7+usUK2GahZXSmN4xmmzk9chAMWHq/3qEOGd0lCwkCmLzIoRqc/mjdzBeXhCX0/9rm
QdMi73KtWxOacghIxkfn6l3jBk91MgjW1A8UXoyDwg92qrRtxTXpQ/j+2grjoLTT5k01FTsgYImC
XWhKIdWv6fAPFFiAxHBGxxsqmqqtxSz03TU4aBrORrNZdDxTYOoHxNHU3h/EZD0Rsztvc5LbDG3R
tpcNt1Dw+1wC3u5i5Hv5xg6Dl5WAYs56m0jr4PBreKgQ25SJq/wdzRMLs+OddhsCKnT9TSIKmIZr
bhfdWbHFVKwG3RSUv5zcwjzhR4qaS3vrstJ6pYYXvvDsTGt40zXS7cq6XMPU2WwtvjXqtok5o1RQ
Wz/V2tWFwLDj6vlase102M+Y6eFllpfu/eWoYH0/JTC/wyIEt81nfVLKo4ewRyKIrn8p66ppyKOz
MNsBmsT2hndQtDfDNEPRJKdZaMLLxmuxfOZcp4ggZUm240xXUDIM2XOrX+LUMZqHYBsB7kJJOL4X
CRgCEk4XOUx4g2AIDHvlHmG+GvSEAJqTVWL0dBVocqnQBdeM1+EvQ7VXxCaIiXDt+i6MjuOog7Kb
a/JWitqx9nKPwSU+ZxUcdASliRUrj5Jr7Rr4D4+OgFXzjLFYZE7AqIVi6g2I7IL/e6r7meyXL5Qr
bHhF/MWXzRERuu8EBQUNHrYtn/tQAd5UHEovY+uNVc+P5R1etE8I7w4v8EhuO9jvk4ZObJ5nOrnB
PP778Zkc5DyKlsSSR2FdluuNOVpkqzoyMjC7PqthIfWuOyWCOKMxJm99Yo4jfZpCqFXuvaZSOSLg
DulTi2rQLdm3PDVJfGivFCuuCR17X2FwbQeXAPe8fdIl4lUE5FlbmphAiZ+N9945O+aKXPczAoLn
Ks/8pVQhynOyspyJGOsrVS5VfAGg+AaTXFndxb6kDDeMJKmN/CSq6uSbqAHQSn4wwLqumWx06k/Q
Wo7FFyMTAeJBoUvD5fo72AXz6bsO0lg8lKD1qEoKq38c5Tsv8/PR+jpnfdvXGIYmI7JBd3T3jBGL
jvEzlxBxFG9n5olk9Fir0bJejQ7kbpSh4d6Lw6sZM/Imh7vzmfChR7KcK2FKur3Rch/H4lR3RG8P
I/mkIuQCXgxvRGqqEO3DP6X5RhaSl/D3WsKpZpatk3mnlbBfyZynM4NqQyxAzB+k7za6wJYvlR5Z
cZQDw8nbhjUGRR7m7n9e2g0lMQ54rR5yOF5Y3l26L4aKmGqXVeM9xtAaFZ8n9G1RRwfb2bCXidHI
1VShZAnopo9GH+PqJ2hSRF5fBkFtWTqaxhtoajuRt7L8uX386zSb8rkIFimotmayHcybSNGVUvKu
VapusYdyFOa3fSn5kAxJD4wXK2zkK63sYyoGkvhE4YkEWzNacgr/zjlWbSZMIuWBwailgM1dywv9
RrNWe6XvoLZ8ADE6TWZaXzyVcEtELfFkU+jmk4w4oFtRDwy7RHktgM7pr6Sy04H1/81+Hr2t01/i
DrKDejHNZgL0niro04zhRXIV+UXZ9OlCOmvosZkXMRD68ApxPv9PprFNz7ITJ6Bt0FiDnImdRLF5
AB8SEpS/b2pn/LLRjB2RVgbLg38TeTgSAMeSPXLiPNMrW5GDATGPtLQmsv824b0RHib9G6fuPvLI
XXLFTiC+xS7VUc1SiajZgGp2HWIIB5pSq7xs7hdW8feGY4s78YnWizXwk/knVzlPgY7zZ0otmf7y
r5LbIqRwJ2k4u+j/uWhWUnNNPCIjUyxP+P4WWCbQUgC9LBlIka0b0ce3VGe2ZiOUuxtp8tt9eyw0
dovxSczteZurYQ1R/Lu+sau+ChtMk+cW/VRcg9uaxWp/sBrJ/UQGRDSSUPFa3pLniztU3YjuC28m
WlKvUU+DLYChZbj8o7bMAp8uClp/uUydHGYVP5RuDdsoGY/Imt5IRKxIeYz4cOQe4haMOws+o6TD
ZR8H82MzzoJKSlBXeY1gOVAhB+d3CyaJdGFfypWqfdIvNRaalwSKEtKgiS3dJQ5oD4lqJpFsIvrQ
HKwdPWaQTpPCHa8dWw8gZBhBd5/fRpg/10hB6+BONtwVq+lcLvshuXm1IPPOZZiSTq5gqIJmkCUT
RyYjPO3t39SM+V4VnqBZGL5zO6B1ARPfjoSI0/r1HQaWT20EQm7hPFDVVkzMcfTJow1jbQis16Cb
KNykkkMzhSZmEhjnW1RdYI8XxhEXetspYiKfrj9LxNt7gmCNJNKY0FxPQD3BgMccYEkMA6g5+p0C
vSul6hsm65vz+KcOr/rTpbpfmG1sMo4skSB8X05dO108nhM7X3gYh9mLCzp171tvGj0+vJ7I+gKL
IdX2iH/jL1QQyAJquXS4TQd8oBvV+f61AwTQh0NKUN5Gx5i76zDZv6eEuxFvhw7AJkVBkRCXlYjP
67oEWXRBmByCRhFaJ+KD5HMgHMr0BFSEFzyAZSj3sJvG4xRGXJi0KapXeZByFWosl81pOrTbzKEC
AThEjnXmotB95Y8gHE7pSEDbjrpVNST7VjX1rp9l8BQds3uHjFEN2EaqTnUiOEl0xdri5t3OJx8M
cvlVMUA113bWcdNPs24aFKjyGEX2QY/CQz3aGEw8Z2Z3lvBCTtl076XlsCEaki1NUUwERx4koF/K
5CAWNJ4sRVybDK6cxcP4z0VXS9vBHW5wTYF2q71JM7TDJVnGLX3xeUeeHBl8xxtkm3/WR34jD3Pi
ooZeTNvNlvgvjst7ruJpWvEe9PfE51+cWCEfvKZ49A9wBD66EeMOgt0VVT5oTYE6Z81LDhZHfX8T
45OyGdENiWmC9qJdkAm6zbaV8vf/iSLpYH1ibwN6a1Q7GQgW0Z9oa7SD3XQNcdtVrENyYMhgUS7q
P8GEr9guS6LV9wD8Z15kacZ97ZQBIeQfWlfTNTwSvWRRG11SlJxR6TeybBHsX4hAWXuednaFniUQ
MWiN8OsoHrV7QCk+nQ71/78/6ovxR0dsDPIU4c9GPJ9U8aWqO26VjCiLkCGIT0C5BYDWWrArGF7M
ZaFSSOCNVdHYUNdqOikT3YJLIrYG6ho3nrY2Z3DOQJytLwFM0bp3L6/8fa5JEB1tdjfQVzn0GezE
TFLD6Kl9vAMwOxu2iSx1tdbH1H/T/OnIVc0ThxBYnEhEUwUMg2ucuSjixeqwaQdb+EsK92h4BnS2
CXqbdoxyub36zvMuGpmE1Nv6uwFk9rt7ICuwk/ctrjNwYaTexWoFvYsNN5s39ybG2RJeXb8uu4YI
DVmqSwo6zoSihipbqjZLWihyaorAxtKd8Rr9VqvjBwYev/Oh7dx1uavo0IMap9b3yIO5AHn9rxnM
Q4DiqQVU+A5H215Ooy4mscnv2QI503dIzPewsDEBR5/zMa1ip57S4WpBGxJ/hF03DXB+2/07A4ec
DKYBvyKcI96RusAOX+5nyNIBJ5dB4ZTf5vhGFVR7nR9WegWZDk+gg7luQvzqF3x1SER8NqTk0Zvz
Y0DguCp5uftHFaPNul8PXUOfRBqvZU1YWjHEJJc6/WHdsOy8gsuVISVe7H5NnBYJq/TSEFfyFMlv
JAtECPJ3tLZG3Vadc3WKZZb97oSW6ZATXcPosP4tfnvk0LN7df0VKXHKCfj25L8n1mYK320WB96G
jGoUDBMac47bpv6Tbwee7iusA2l3DNvFWXj5TXO6y9H77OKy3CAxx99mw3Q4APYqjb5IhGQIzMX7
3FS4K08ZKcNVgihOVQZiw30pGGPpq4IFFPdA3GDnsxvVnTdsYktFv/asDPVtn21P2zrwDj4U50d7
1QVBFQf5thQ2vK/D5Nfgqu8i1PKddfZFLfMJukF9rf8hTCxLJhEEqyfMk65PuPyFb8WXuwsDXXMx
S/UCaEuzgoqYNTrDznAiPBbnAiEmD+eY4vNX550BBl+g5XSweudbZf//7AvLdkhU6GiG4K+7v63y
9MHD62ELBYUos2thSqe5xFxdh09p1bvpLSfTd15MxP4mrmbjIYM7oRl0SRTCzR5WWM8cvQ/1r9WI
hISReIuQe2muOGDlzimIMvKidn7lFyYT/Gp1TquNFhBDnWjrQIZjkzJgEC9ZXCZG0HAb66DoFJ4P
B0FlhuIKN3KEQCGBuHer92W8DzQA0QNlSYjbs32eG2ud+6jXV0Lq82fTOWr6mA00UzecbsF2aniW
psJcZ6ONjJtINJTkXAzc+KXeOf+6XMmXHQCDSgYNIcY7eec98WPEms6PnWIVMkCQ88lRcQ1IofFv
wYJUdLtdMaavvgeJ2PzCtkJUeLahmK3TBNLaMxYkrD10V6y3t63uggBuuoYbVx7aARGsIHO7ugq4
I0YM9ZWXnyUMS/eyiKatk9K/98Ut4X8GH8/dHXVWGotIWTkdS7/CuV0PsbRQ1OOET7qgI4PbfPnt
l0GM7bKJQDABd3yAPCJUipldhzXN05MqsjZnd1yD8I5Tb6MdIEpjutGiKY51DZsc4ske8Lr/eHZE
pPVUz9hWRKFu0wEXtIEjabwvP4swCFWwqytZvoWVSAIw+T/qmRoUQ8fbay/DweEg/Xbbjh83p5Fl
yKo3po1+yE4Wk6LVJicOrmsE1vCjBvAQmWqZUtB5GyDlameA2k9M5EUDu+NUb+ygHH8dtG0dz/ZG
zpd7pId820tcHkg4xDdgfBVAhfbkFfk+i+RcqR/5P5nLP/aAr92lWjQGUS0/L3j6S0kyo1iS1/Fb
TnQtmlN1PfzXAGA+WBzBdixyVD4ogkENQcSTrBUVb195e8vC1+mnJif5rBTVQgyTWXRO5hvDQLFx
qt42KbZymeKkWoROy4E+zJHwQwW1Vr5WKT4xRIBYZccejMrs2DrlsAyovsb45t1OSOhkJul8rhfD
iHwMBq39DImflVCRZ0baw90ompSOks1GRBryfOndeJKyZl5bxXscR9ls7bF73yrNwK4t07yztiB1
nPp2IBv4yupD52VfKyTpt1rT0Jy18b4DSLsGl0PmtRHIt8nmvJ0eOL2mK/4CX/598mKJnZn5K6yb
gXgxwMAlkUlYIyXnOVeP7cKj7uLjCbLpou9y5iB9W/tSdIWXPkig32vY+ZRX8hVKVf3C/rJmEvhZ
SDjfiLVHjIt+lu+yIY4smlrt+3AHmu+9gIOzxcDMATTbbKdDCqgK7bzkzjonSZGyYJLy2FrpDW3v
nG20VE2/R3bOqnHb3iAP/GvC6xc5ykjJOouOj6RZxLTcB9TFqJswiM4B+E0rp+D6xLfuuRRt/+j1
/eYXPSnZAi0gETNZg7flDK8g9iCbQPwof0WIL7lKR60L5y9NOBo4eh8uSSeASiheTl6K/N8/l0p7
trOU6gqun2LqC4OjitFkqdFututTEEJtno63S8Pn5xAQmiuuPIDiHz5+W51kj3SyEGo1g3QxZMIB
PgNcTMs0cWRT91ZR0zrXmELnHQ7cKq4KLlcP8hk+hts6obbqID4PY+9R7dn12aQXmIu73NmSJ77W
kcW1UTmSHDcrILgeqdOrCpU0LqUq7/wKYhASJv7H3JSnIdSzVDeO3G/TzC4txRpooBlfgTF1a+FF
xNxb5F5Rx1d0n9KQU7MVzJC74900DAa63lIWPnhknkG/iObG8bpHeo7f3rFxN7weqvBtik1QZ3Od
scaykK5D8Hl6rcFmFQ5rjZOL+fLbGgAPwSzcdJohPBeg5RC1iBsWfe03xKlO3sYo5saFRzFLYuDj
rXFpekeK1/BT5WRaTkpet8tNusIA7wQz1sGxhEDpwX+/zPOvsLecOpj1JWrH3qXGBP5n9bvJKonl
9AceO8rqrjfNTbcJMP3KtSrn0aHarna4UvUVQd0veZH9elWVLk0ysDMm5FV6AOpCG5dejM0qiXXz
E7MRuZ0FSSAj1IM2vLA5XiANJaeVk1iuuUSfyEnQ3y2lqqof2hdE3si3cK4P/KblcH0Ya0PCPXGv
UKr6Ic2/gl50zNG2uGv1ND1TRnVdquHSTXCMbW5HMtvmSaaH2JCLx7W7GUUQX8SAXRp9StWSw9BL
+OXurZS8c4uxxyGEiEwOxSVn85DPCBLpiLKktK4SMN/4JVkNDOttUZ8Yux7OWqp56wumJUg5XSol
B5pBXbuTuWQqeXkKaTdmlAF0ZWce0qfl1pD1kt4ERH2LbBlCLkNp4O6nK4a3Cxey00c2yzWsgf/v
9FcUtYmUWjNiBWZXa53H5O9sZDRnyGNG3UXbdOtmxLVKVWBe2r8Ab8t8KXaqmNwlvGWYbfiPOIxV
fDnTOK0joxxoDEkuYHAgRUejqcjS++TG/JkXETAC73r0BRYaRyH2/S8J0JVzMKmDs6DHJTBOiC7K
HHiG2fAcNWig0hZ5HIwzlbGiHSFQQuHXuMGZ5ynKpBevDMleJEcoY+NKuw5CUpyArWIgCumuW+tR
+gu6EecluM80aHxcxaBbCP3uBQ2/Aa9JI/ezavWaLLD73t+NHKzu5NLBPE3lGZoqel4o54cyl8u2
xUeZwN+xKP0mUX9SPLEtVzX5j1FtOdAVi9fatQodRYtnWwg2w5HTh0VjAlfHJQKRTX9NXOE9EpJ4
aYyAp6J0l1+kMIt0P93ktqXaBS5Q7SmSgFZAavZgohHCw0AC4YVyEWV8QTIZFLs1m9J83WIBJ9iI
Oh+chY52IrakRCWD9hUXqQtV3h1+VXx69RbxNAQkCTHoW407y/NwuPNaepyp6SGKF1JtYhUsX0vV
N/tdqWAMm84RcEwmip0ef5jyR7bBe/9tvXMBETZZ07Wo56ylqdlUXkQrfknjxEX1jGd3gi2ZzZny
rlhjXkUnQHGsP1WoOMpv+h7kNeqg0AlP4FXNIuRiqZlPhVmAws50tc1m0UnLEixonhxx3qPVb296
FB8fR6ib0n1TiMYLQ6bP0jPD8vKUSShfcLNST+i2k4oVN4eYeNFfWrTwKoGBlbQrnnTkr+BM8hX7
FAr9Q1sPXbVETH+kvWtMGvPK5IyiDOXZcTvwm4shth0PdTjrx/12lxh5g1o/Fv2HFmL6zl2A/9LU
GZaalmBeKRbHnE7izNgoQaZwrpV+h96tRm3cUrTqD3C9k+JEX1TV8TSRTYM+w11uTkI1osgfetd5
TYUapBuyAEvPoIhBw4DptyPAt/KhQg8lC3R0J/g8p+w+MBCeNjXWbv5WYBHppxqcPvME+QT41Nkt
7Ue8tvTOOkH5q2oL5ciWdLjTbewmxGGtavcloK184I7SqBxmJTlYVHV0S/eNR4FXVK7E91x40jnt
xpij5WCPy8fe2GPB8WJOXVfKmXN7D58ThSNptWvpLD+lxlsXX43MyHzGnlpPFyqFw59clVM3EJ1S
fhsQc0TAACORS8fQZbjsly+essIrpQGgSAYSXeJGDRoB2nRjJ4JS+0rbrFcNc8bUSqxzEM2Kzgou
1iKmpbj9gUMPpCYQyLKzCz1mTGecfaACsdbUidJ5XJBqcis+Vck/7kURXwj0Tq5kJ+mJZsyfi4HW
AiheProT6QzQRlExBB+sg3PPEOGLFyPa5CBU9UyeVnwTpt/GzQYbtnVpGyEsXd5AjAYZa3hTX8oE
VaFvrQycS8R9R1mCpO8m34G3fMVfq9o9HwJkhV+qzYaOni5XK3H/XzIPGIGTd5LoA/097F3Q79mT
7nWAP2EWv76h4nNnSj4x0yWU3VlMVs+Zslcq/Xt/E1ObzGpdVARKlt1PbpbtXNVtjzzUEkBBX40O
1hMkWv01xUHQaGHNcC6zu4+nvVqFg/ou5UFwZtmVp17KGBeLbIHBdFRkA7lvI0IKmmWi6EWxwWiP
0ODrwdmgTjl9L5+TXSIiZs/Mwb5LT3G1tlqactGurgNCLLyfmwtFXYq/eczaGCkkWie4gPFyNQZP
eYT5miUbNWZOXNF1GayZSO/ewMANd7p8pNbX7CTome6L6JwySX8Ex3zSVMG16CzSci1w4NKfV3R3
zV0Wph7aBW8Wr83/eigzcFi4CBq9D9YM4nYsnMHEJk/vgYcP8SEYDc87Pw2V2YM6TCJmA8+PrImM
jIYH5oS5687L1zqhgbeNNjcaEbYOYSIqkIYSZZWSR7xXyllaba4mwbo/FbniPVUw4L0eSCXSVvzx
AgFyhCLTaHe4wp6zvSxwm7eSLPM1Ikgcou/VNj8Y7A/Bmo6+sUu3NjJKxkU5ZTByCCrIiy1OVuNd
SuzKwdypYQAK1PHV0eAvfjfHDtp9FeKiEdBPXBnV52js+pLq7ruNa6HDqzgVxiGeJPyPXXg+zUWD
P4xprmMTkI8QX15p+XLkj2NrxTgEmjZsHqsxVkDLiojm4bok8kufAN0UaWhP8rOj0Iy5k4orOXQn
IXNvgWnF4A0/xM+kVkKlNyRa3Fsuvv4OKpOAuppEuhc6Lm9DddgTioELGSIxqFJoaaBJtZ+2mR+6
inVx/W/nHuYgro1KUAHxxfMZf2PfH9mxEzVedFLzQVs/c3krAp/MKxfrOQ31fKkonmxbHt2ua2xs
uyW6E3JV1Paua4o+YQy1T8o5WXDcBWBLz5bU26C6k+BiCnJaG2P7bFUODvFV6pRGk3isSSJnfo1V
vGrbCkvIIjkr+4lBU9W11RqAujYRDuWfiK2PeCcyNZmXzgDFlHW2Yw7l5S1z37qESSFllxuP7iOD
G5+typrjWVsVMdbHtZRf/pm71hnWG4kfiD3Y40eMMqbboZZGoVIb2ToCzdnoJDW22/grUGLAvcGv
vLCaSK14T/u3iAqLQHGdFEvumoM5BoqYg1weeueT/BkbC6eqi5/b0PqzGalUs0Fm2aRvP52lx2Bj
/c3A9jgNyY+eObCxrFP0tQv2q+iCakgNe1V4booOzJqdLdixvV8UafKX+UA2Egb+KDE+jUqk2Una
oVQHK2wzqjWdbScU69STumFSu0tEZT/Uefh9K6U1A+HCzED3ecdzPCtij7JYsbgOeRHEImirNr3P
z14lGNqdndzvUegyb88v49r8xKhVHefSRwu7NZq14mb2yEJkjRSpkrinDCQHOEZXexVf5GT0aoF+
wX0lHyOqUakdGG2LJo+LoxU6V5hRF2yeN4eG++N80LOHgcVjWcU+bUI7ErVyDGpMO4uqU3HnI7i6
207cw831+55xcFsH5IvtU78b9OoNuIxnx75+iundK+avTrnA2/fhhcLbBE8JARJN4Og+CUOuQDbm
ao+9j0enDaFI+rtCyDjJ6skjcwMI4VvNnn3x2tSKCLHs3uwI0d19o+vH6AXpi0vIJ/wuQcFxJOV3
HKHshdUJWjJ98LJdjaTNkZ4fXpgueHjF+AF/nmc6vNwSkSqs4eMJB3B0WVMe45nEEblRRJFqtTuU
xdzLxJaBICu7+ar3glAkx5/1lAo1Ss2RhY2NaiWUQeJh4ehPffxeOeQg9HqbajqvwtDQybtWz8D/
z+/FC8C6nEgN2f2RYm+Gj5WPj65enyYCtZBjfxaAnvg2pKvVh+UsUO29Wj4ZJUl9aF9nvfN19dh+
a402uJgrKGkmj0qUKXNZiD7dt54CzkogLmCAzbeLTUj2QQV55mUWBR5SERvnqXx0uC4kF5DoBDr/
k9Q4hwA68fWnkdfhwP1emgjLHCTUUo9B6SiUfvb3Qb3Sadj0IMFuAxYTPrk5F9krjMzxaDCcnNhq
hAntsVe+t4pgQV3ASutF76gRXzjuVpOx8rd3Qb653F3bdHaD9xTYtEorho3FiOijYaIiD57JtIlE
CYejHcOYVuFvT1hNAaiUCo9W4TmsUWWgpFksUzVj1/G9wxHSiOgOug6Wu4sg58OL9LsmNnavTEsr
An1fnNn98DeZZybOKaZcNCxbjrUhqbpJ1P7QdLj0nnhFZoSjtVH3InC+y0upQAYRvvmbVccv0On4
4QrHDxSHPVkrYVCmGT9Ar4mfNVlzqdP3kbCLc5jM3o3jIDpijTDxV6b8jOTfFlS7XAfi3W+KX+ln
gUAk95PUw7FEOEI0uJsx6hh2jiG6VErRWI8khq/qQ6Ser0r5FpDLrosoFW0ZUeru6NViWF944IG/
tQS98wNiS9ESvQIuhgbL8N8z9M79F2MLwjCvAZbbiBqI/TnMTGV3nvbqTy6idZHZb78nBR5CqKTq
u1rYL0GRAHfeoejPpdgfUlb7f5aM9AeEb/SLq1OwN/xZUn9/pVz9prwQpu4nQOa9zD0je2qgPnuf
uekDqrRGJlKUcZlmA6p1S1Ue+gbMFMrAthjMZ/Yjv4ahXo1IiFlKpUe/1z2XiCxkgO3kUvmnGhbA
WJvO6WeR/C6yLpR8Tg+6UrPkwsrQPtFuIToL6NMMWUCIkjt6BBhD6TThItNhhnb+LqwFKFFcjxVV
UmBA5th2lP7yy0FEDczyf3rP27mZpc+pFRKV+7zyPNL9AcsKKK/iqGbIR7hX92WA3AmhSS69QhkQ
WqVQdsisXO7CN5kEJsS1CGX5SWLJQRl7cXE3VDyp46D0/HMPtOjSGMUXRNsv+wox6gZm/A9AH+m2
HuWPcgAVTPluL1YUVRQaQN9yVdTsCwaq3OkMVslt6pawfBbve1Kyru+DHcAgE/7IaEjM7nWul3Au
vWYq2yCEIbnEnt53ipn13vafph+vFUFv6M/P1RVo+CNpmaIsLHh8qRZFHrZrZopT8m0Q9Pisqops
K0lRhx8Gr1weGN2sSW3+O9/YIYYNFzkTyu98McdoWWQ1qe7cxHkK4zy0JdvWchf/ZKfXL9l8U7Iv
j1I4Skgs73vvfu1qxpOlyOBpogFek9cISUtkjZWdcrTOEQzpZaxUZFTuViK/ubQzkh7EVNNdNke4
31vPuwNPmD/SbA6wx7ogKg1/e8ShAbhzK9DK6/oCDAuF5pXm8K/OgDa82CoQ0cEamtQR8WnUwSOE
6OGi6889FBYUXFiJgJPmf0mHgax8NghleBoy8m0anXUSIEhTqZVbLqJJOfSH4lf7JW06KILkgbT0
FxiXALeeMf/nHN5d4THPkPb3L53K+yUf5wk5brsLR8YhWI7OAE/nZWuSmZX3B1rRi3YNyxsly4BU
j8uRhghRSFw+5dIaEaYAzYZnkkqs24elyO5pK/uRXMrPvlwIu20PfJYmruFq6w9lyK/itNI2MRsd
N0zaoy5gQH1E+lWqGLIUjr1W7LWeHoxAt4q2iCLhB3LAhmxNFQsSiapmfzVYFMxyWH5Dnfb/HNsM
inW0MJyKU6FIot8777wxPidUN/13b8wDe7klMiukQv6g655ELz7UlFpsErHlrDPbRv5NQE/7dk+/
iZCykNji7CTAbfhGxFdCmBeCogOlz2YtAlxDNuNMIsRQ1ou7aoHLaXE32BcghUSwyzVFhfDLfTms
u7xVZWicifVZVt1DPXaZrrelRXqGSyGg6+j9Oa0xQi2i2SiPYqCC/U8CDnoJNTQKTIGWnhWO7oHo
iMFbfCSi7nLlrgsMFImGe+/UTFHH/sZbTw+WD3OQbtv4Q5ZU2/UqIhjJBMM/Ub2iBsojQypIlM10
DByJQNNECr3lle8sM3upzvmLIIQ/5FukC7kxUQn7C6r6GigAVrcN0B/4mUDozcrf5mMsl9h9hXzf
zckBQ8+uo+qMHTA5i+YoTrUSh5d9taLNbL0lgE6UU1bEMmOsJwWT8OTKZpEKOn5yFRdgv5MGtQRN
cRdnRnVCuqOYXX2Zu3hFc5CtdwXly25ngLCLeYSocb8v6eLJuUx4ictROu3rSZMwI5qsXJxnSsnq
Z+3leLBd+6nGMzFNTGEzxTevzeUNHaYPRfgoYDIN57mI1RPjxTuHwafMrrWw5iBxxvpsYa/jqyhn
WzZbBcedqW2zPdw5Tg328VgRiCiSK3p3CyM2NDQpJn5ny5wG1oSPaxPz8lhmarEXgMY1+ClhawDf
oeqgxrRWjyhAEOpOYhvVrqLW+iV0MdrWySXDRxMg2JzRQ4+sehgDXYIktPukuk701H5lGBX1ZvdE
9z5H5bKTK7N2zRuCH726H+DX8O/4x5Hdp39svaX8z4lXk9FTOr2J+jTScQ2TDIHdgrtgXywiidox
tWcEvPZ0u967Shi0MalErSYvLIRmgR/u33pSGzk02V9AziCPcl1eRytbPvH5kO6awdIaBd2CpVuU
vaj1a/MgcHbAVtNcb5jxOMTXFHdGEgj/szi3Ht/BBj65juFDv7oqKXGHhM0Tk8dX0hDVUhSP/rSI
lSdhtCrPDZcCuZCcKLbMWCiKrYtSqYwNB7Gjefk543/z1ISmmcDkVHfM46QYOO6lGmnQ7DpOMeig
MDsm1nfVRVYGCS9RmVy9t51wFGEkXiDk6FrXrXKo7EVXTWle0nmLxJUXR6jkQGsMNF9yWk7Y08u6
hQOToKzf5t/Su7PLUPFW55S1bnOUXM+SgKAMoZ1RcC01QQduYztsAMSGqM9083SB5SdkpiPddx/f
g4kjUgoZvmhfYJ0jCyVmU1vLqyDf6HSC6G/KWO1bjOhpAq9aV8FVgZeUYQAQnxfJXjmXiLhTDETi
qWITotMHX3FexkeEojhi2iKDtPAQIs4ZJyDmUEQ+YLw9y4G2/BXjvCIPOt3kHYl+tvbzveyP0gil
fHZMP3jHCj0pbWN8eCQMzNOr8yEBeCgEwZ3oxFg84Rd+p+HcbNyR0vrPdZHw9QdnBf3KkJtRfuYY
HjyyeV4ivYPPqXABFOIsFYjLXSw03LS067Xg4ZIsPgK3hbP2KT4hU559oWyH2CEPaUor0G/s05oP
h1qrkpNq3m57o5HL4tppYRKPJSjkvhdTQJpM9ePaooEKCEb4gRwVtinEwrYQCM0kaGrFdIt7pzBy
wmDLddUd/28CsJT3bpLuD39CyJjJFpyQgEMlfkB2E+jRPvq7UOt6ckdVN7l4GAlrOPd3gC2mL4zB
Esnn81qElxIMieuwtkoYY0nF7uY2pq4QaQAWlYqHvaj1h8tCrAcZCyMVK9R6W8T9eTijqPv3ThG8
wkrgxc/jWKq5IaFXbk786BhrVzNtXN/BpAJMARhKmjbMMoCMZ1qDdmEFxTrRxxTq+pFqURz6Lp1p
fVBX8ufjhVAEM9LlHLl8JBNm0BLPdglfayG3BtK8d5I1/BKQPGL1w+PWkHU7OZeOuWkmwBkRu/bv
9vo+NLcWi4uZVjLhB9fXruvjs4bGbloMhJhA875Ry52eEIxt/Z1zjlQpjln2QkzCqBmAkFFdEhaS
5oecsCEWgBs+SWbJsOWRSrW+tEb0R3fRnV0/KzeUfLFaKJgCBCOTCfl0RmxcbiODtn4Ck2qhyyHr
bn/hvvNIeVBDEX+zRM7+irdDSWH7PIQNNbtg80c+63eG5OAfWJm88TOD61QKRMmdogWpKyq8AUzE
lTB96HHEvXcp9sTYpN1w+lFBgHAd3QX9Vum0cbXvFxJb84ieYMTUj5t5Xc9oA1Hv1CdbcPEZ+i4q
63bWBTCm/5YGeQ1hsp8hQbV7WoCe903Q1DJtYJxSN4OtjCvwAGmxLtanuptIDVViguilvDADq5bH
iFxiUUzwVQtpMi4yprTH0PDv1Jaz5gyPYClNo+GSvGMDVKleM+jZ5v7N7CdlDcHZvhxb2/ABJUNW
5G8omdSo9DZNrpfEbxmurWqsfD+884YToGm8o03Lztnpzuj4CttPIG0qV/Y4FxhLrNyQ92i/PDbJ
AyPI9NKE3kOXP4nXlhfw+P2eTDQ5P4Uie2Dwlksf2UDCBF949bgj30InPKb66GeJgqAU1ld8o/Sj
nmzjT7HmLwxHhW6Bo1Ou/6RlQ0feryewlJRwPlG+LbxFoMF41EsgpNvbF5xwEboXO2S/g2dK40pi
jgkcIN3Z5UQuG7SQUMR3iAmLKmCb60GHirAUueOdEzV/JNKC4MkGVTCRfpyaWlVakuQYmOh1eAqd
XiHo6p4jaiW7lrXybrEiazIgqgs7OAsgiTB+82MJjd7c7Ci8Md7/RHJsNwN8lVkjpsxn7UmNNJwT
ZG9yp9J9a1gCmdkQZlujn4QYz/I/jQL//Kl9shhQIqDAdGaA44OZ0betzTwqd31AfVv6IstgUL9B
BD7n6M2mvyCRa6SeCVURWZYKOYhAFBkwz0/ERE+J9H5QDRCHI2Z/BBcrgMGVA805/nQazZOJ1usC
E5He63iw54ugSlWwOPq7dJXpa/4RAaMOjpmUTNl0owKVoJUss/QrUNhRfd8HKlKH+V1qxw4ZJM+s
yuG24C4FUVpK9KGPjWa02BorAsetVJ12C0m8RTo94So+wYtzCKA1BCAffc4bHvhJ+KAzxYwD2+4S
/plscmRCpCFmQ2t/6pQW5rmDblmF5FCyg6qifZkAdoxZ/mM7QpvLGbF4E+u4e1N2nugJRP0d/kJG
dGF0Lj9TQGb3SLbyepXzSwJFPq+j/0PuBHdHZgH9I7hqF88n4reH9qJgO9heJRVZEeZeDfpNjvIC
2nLPeiB0GDZHHBO+Z4+SES6aiVV8xtMJ+rr92IavYwAq3jcVzajl0LdzTBft/4PVOcuM7JTXCeQd
DfH00W6U5JgoZZgQ1ulJL35cmvN6HS2VGfq1+nR8RTuaffY3cnXUqBPFuKas7BilPuTrfP6syy0N
I+/Je6hBHgs6NlkXtIEgeFg9IgT/nfjBrmWllPg/RDT1/eMHl51ueSevC2r2Wh6EnnRd0/d+y9cn
w1v6S5DZfxJwgKgil79ZzcDCkmVwnqapPcuhqIguI3WoH12DabJrZMje3Z8F/cghYu1TfZMcbYYF
6j9F9ty4sLHUDhlMdCkdAEpmh7h7E/bwqxhvfvXF1gPOOGu9gZlGlJ4JmDYfcMOZ/DwFEb86qFLH
B6aegiGY42zmIuiM34FCm6iKSLeGipddta8r3mbloH1Y0vAMDTotPFdunH1ry93FmMWvdo0sXljE
OjjGGdavSFoeJIlFRDSl+hR+sBR6HtkTdmI/LVw2mFuEVdd8s1aycYKScXBokgMv3fBHT2VWBw2z
ASuZFGNU5D3G5OqwI06MF6hfn7oR0shh7EPqYpIKDBTwC8C0Q1xw2SPsY6U7P4esDHxrEX5JOMYB
N+TYOQT0NvkHCWGKyuX+l3GrFZkhJRVVNhTN6Fjq9Q9ytYoyKgRvA5H5Wfd93ORWz3rEvFjcvUP9
zLG3Hbc/dQKYAmmtPuSzYoI0jlMQp3SZSoNdUTX+REyRKbXPH6ThloFWj6dS972eCPg4WLB5sJC5
s60Rbt6BmuRDSPKq9rJfqD6MssJxhK7L4l/zcggBYpGz7ywRQ4rk0FUiAM7UJSqmzaDDMa2yMjJe
U0Ncblva8KCvQPLeT5TsV+0efb5BANq3mBTeWg+F6vtZlluR0YVgnMDgzcTtRMY69j1W/T7UIKlt
GCdq0kSiM6yfQhgSp3FNeLM4FvQY0fLqf39GSpr6tm5nCaSo/goXxXLXouOOn3a3vvl/t/NRx95J
miioQDBRS3nQlkKDNs/bQLpdQuxMrX6U3zIMzg+ZW1yaYpHFjcrZuNEA030b+sGSUB9DTbWy43DP
zjgBOPdC8Z1UXWKWY/ZjU7kJrs8S3BMOLsV2LpESXao9sAbmNURo7+E/aJN0jXW5XaIarkSJAUHD
Q4+9V8a7tvAedJYZ3ooBJju8/OBMSrld7HBeaBsr6vNuA8BcOpG0IzUo4d2fXL8nI/fJxGmBxGn3
zm1lmR6Vvkzg1sJEx0p4DrNiyP3Ysk7OS9OPFESYPxoEAwBNTwkeHS40nl0KHLEjT6EJ0OruZGLw
fiubY3VhiAxG52HMSzNjTWNec/NmxUgqX7O4yNK8Dsx10phPdkk2jYIpWQz3Rh4Tgs5aqLpKHK5m
dy7BiFjz+WnB/CPpwfhfux+Bwpl5Dojk0F2OiGaDBBqUFkKjYSPB7mw/wOF7c5sJuzRUFQ0/3Oto
2aeDocegZXqAa+k98ayvermYDqtmWUHlUUPjxfotzGnKtrfcQoupovoDIO0TOeFI9nOdUAUSJuhz
YKmJaN/awpMhlR+xhtJCGWDUaAU6GDMnc42npwRuoL9iOaHHcVeptwWsGo3F6klswvLXI4DluXvz
pPPZGlngaNcPifDu0gaqHdARpLjvskcs5RAI5D3zdu+68cgyAnXletU9VvCUkDGcXyV38SuWnCk7
bsu/FO0F9n44H0x1IZ2YTMs/UhDAvYBuIFqYcNEOC39wG8htUxmfztgoVVWQJh9cuIqgh6AI5+pr
BPUrbRmjasX2UuXIX/zOILGDQ5c3HKsG7/9JT3ljpxgr3BpT7ht9eg3cehs3wVndP9iUaFgi6aP4
qyZ0k0njbB96E3LrvnS/g9HrLv45sIkg+GtAFAp4iPPY08/xKCJ4v5V3JUAsnf8SGDx3lmp3oY2a
m7QUYUxSQeEp8VjeLWFroJmzBpZ/X4EO+deNQs6jrvprQTJQOLMDp/iwx56fHqu4TthNxqrDVH8m
hL253ThWvrpG+lkYtZ+i4mx2RGoXaJmsMX8KZz1ZtSYN/y2YALSF2uGKduTSwQo5RGorvZ77FND4
e8XsCaoDv4OaQgI1AJDBiDnNjUNQVSAvP/drqxnNkJd8XRynuzw/JzzNT1VWq6uYf7R0c1E025uD
7tnNcUXuC0TxV8HoWWHZAVc/Rzw8jzGz4AIw821WRCYqg9dkzyLqIl9250fzP7EvFyo8vnovafWp
/CdYXov5Twh0mEegwJGAGXN29dOSp7mGfWySetoX/oL4pgL/OfBYf0+5cwgQcdXb+HDBxbaXM/I0
rpzB/4nX+CeGy4DyriFolFErOTKJJaW230qc0a6VOtS7IASRyYlBzeZLqbCYoUTd3OYQKO+WN89W
hkdo9wPP9Mr1XosRzWf+oVjPC3n8sBuhlzfpp0ci79jtoBxsuDX6Be1fdlObKBlRvNLklePkDAOv
fzkSJSN/rKOLLsk8ehr8ZLHU2t37O2fHmF/LKWH0pWXAKSESd39VzrwF/7I1swAY/JBlUSwfVyHW
YYIQwPnoJAvpqbcFPTwOYchEQQIpmPyMuuJjMRGlP33cbUI6oOg92Sj6ZUEdx+zKyZwbC3k+/jVp
hq9GcxMd7IGqDOpgKCNPj9cLC+N7gNk7AQJkQmxyBJMf/CswgH0HXMiFJwsy+ONiy8mMpCPlaBY7
SAH4xZrPy+4FNv6vB5Ic0ZoWTyB187gtWSFQd13iybF/TpwCwAOSWVXeR4oSjEj73AJtZEEs4yUf
/nPimUGjWD84ex97CK2NHT8fy2QwiOtwnNgQD96g8R0mh0/bFOIpdHuGLSvNL4cbYxPa6FNM3qVO
hqANDzVN9CQ23Y1a6yJoWx8LZYAsc6QhpiGum8rcLGfWKM0pwntzq456pXqgg3Jj6cAKOhpMSI6v
dynK08qOg7yX6Vwq7JL3anWVeBwBnMhqYH6mcpp/1+N9n3uiUmJ+WmVAkr9LnZcg170f9q98N9Ft
CwZtx5CIXk2HtxNdK8dd9y5g75OzdzqBKym+0FEWHJX3k7EX4Aykl4PKRYB+1jUePy4tbSatvM5U
Lu1JBFEcVu8L3Xk+t+IyHF3diquGigPrDJ1BSmjau9UXLy3myMja5M6p8eJzg+fnNH1pmcVts/Ee
7vx8J25VyrClsqjh9uGjSnCCdOO58SmLF96ySzcOuAQwegW3swIPTIZSIknNDs5lkGnbZp3FDXr3
wMV1ETGWIMsJT36aSYVQHzORjLHTNw0y0IyPJ6EGhPVNmyXegiNFEcSHCWGp0aN3F0nTsMj6HrO5
xMrGCZeuUtwlQPNpbQ6FZLsq1MBs67wAAz7OOORg0nwF4L4Z5/p2zOaPa0FqNrM1L2jzHe9CLCxY
a+YUooHCHJVm9E+zd2udPjlPb+KAblv02aQ9ngBItFOj7mH5dJ25i5BMXnIwOJsxiqlJDTNrWPsB
ImO4nLcvEBE1CBANcBhRumaKyuRgo+m5JVZUYok9wJ9XZTyzASfLgpWpWDvpNoIhXIWklnY1JPzD
B9jYxFOlF+zxFgvyqEBP7G86UsaBfGKchqGH7Wmkomde7OFzcIgFYk7Qzttd9Yetf5cUHGm7sbdH
EIgMqR46yQuKV5mIXdqmHgX/Tymn2jHLrUTeIPztdffjk75OKhVtMS0T9jGKXoZOYDqJQkJNBezl
eafziqDPOnbn+D5ZPjm7Jz3Wb2yGXhqFrTU8VXKsuXil1EPkBblk8GH58hIFnKZGwyjzbCC2ONYE
+5jACVn4p8+AnmXRGzK+bvs83EdUvy9ya/lVFPjKrYhzIXZvFTmMU6BOY7iMb4Lj1wjBoheSowE/
K5jwpOIpj7GO5Qzff1eH6EMDPDg+qq+ZHgxJzfq8WiMfZAAfJuYzSDJG8Wf+20lauB/xMkNvSJ3Z
GvfQnvC7ovHxqfwE8WHQ4WQChHALSpE0b8Xt0XETjuyR8hl+ynhG7kC4URyaF8uYn416mvVaFxs3
RAqaUnDDnsOb/G0Vx9by6tEVnS7uYX1YFNFgAIxW+VmxThR2lmop+yUYIjW0R3tLDJU3MeXWtRR0
bEbo37BFQR+FIUbQOJCc7a3vQ2/Gzgnv9ENE2NLPg/X+thCgPYaII1d8nhHA1yXgiiiS2RKy1Ks8
HSuly+cMZilgO0aOdOGOaTWpbJXp5HIz8A6XoB/I0zVmBUsSH7LiCuuO2qzb7KiL86JNc/99JqPJ
MDh8lkOPfe7qGiltylw7yUQdEbGWh/toKE2sCKB0+ZbhIHrnXjzWSprTZ5sFQbNQsXHcF4el3kr5
24M2X4AnLhJmqOs33Wq2+k5GvIGt4TpytATdgU8HZktH5jL6M0x0ta7FNLBY/qXZ9iZJ6O6ywVkt
knuRE/h3Cn2lW5HGP3yU9/RP9bUO6fVFauQxPrEzVvOwDe4voZZKIuOLSkzmGQf1XAC9oIW3LeFn
9BrVG4b8hKf5feBXr1PFMNHtRs+ZcM8WGaMvsvOHjuoOYRGNyOcsrvGY0hk6C8oLrEXs3s2ZrvT3
WcNMav/0SsXdq/YnwJ45gUY0ZWxoae4xd70T4mn8uKf6EACk9hbr5KlndCjQZU8iNepheyLc1TKG
rF8UAihH3Y2S167mX3vsRQeZu/X2WpW1EHe/9ikJc69eRUC7Iiex2vX+OVMUSZ2aBs0rk7Flin+G
gW3wfgAcWtArYAECSKmc68mQSjvnGfsPKYzR23bNcmVgmus06SqZDNj3eDwrbgp1uwBMf2CaTLt9
vLkBKHrbq6SMZTVB84OcVq7DmauX1magM2wlJDHHOm9/cAqfeOSr/CD8rqR+F6BPWih9SzlLmIbV
dtlUgQWNJr9oRJ6HmegbqNPDlGNZa5lmNUKT6H/uxZXrdmTpIaN6Cez7z0/jkUqSOfZN+UQBhRO/
peUmBxqJa0fvuPB0MbzTHWlaM/RaY+GPm9jhB8EWwH5DGjITyaGKNxoArbnaaoG+tvxp3/QG7DvW
kUdyrQaFkC/LheD+fLuvHQx6hcKmySHzExIIIZ1IIRLtN/mZbhcROhF+dJGHmFfHmKWwY5+2+R3X
U9Ydk4k4YPo4o55nOpUxL1/TvJbNCYbCvnLbhdzS4uIYXHB1gFIiK7ZDmeXcnvJZIHnrVHLUenaJ
s6kBom2pgNIj4Kuapb9fcKNiAg8TdZdWJq2HswEDbuvM2b5C48rLy4WuEpcApoId7oT7V75Em0AN
KzF3QGevyusM02jPmCBUI4TNhtWOGQ5fKiJnrviPjrzTPwgs70o1onqnJ3Z86Vj01eN2qe7X/mTl
O+Zf5nwh8t5WeY5wCIl1HOaVejBBYsIaxF73ycr6GHVH0eDFQ0o15IzwLMxY08lvpX2fGO8crmvJ
UAgeO5YaEuTVkyY/MOyjrrc+iXSTlYiT5XEvs8FrGuw6gX8oLgvQXzbXg8fPhp4qxaOdVKpQ8NlL
f1WOcxJyMbY1+hiTFttVhraz88ghxFcmcJF4kkrsn3VxKztT1A/2L2ZMLk0fd+Vc9W8ZrIe1LGKE
ME/G+va+jY2RgdnxgEK0Ztdlt9Y9ossxqz43fHxJGQXjJBYBOyYTS9Q1LqjUAV8is2C8GLbsgo99
1sF4XzFyFMiB+HcuXXNayCOWz0teHLp6DG9W6FFwihd4m2B5N0S86zYZ2V8l4RfcYWVErWMEfWOT
FPT5Z4HAvwxt0UterAEaiNybWJyFBichjAN+tvD1BU3MRgTr8V32vAtGJc1Rdyva1T8rTGpncZJl
zPLKv/+fWmo6AVYkvldwYO90pDIaIqtaIKa8E328Csdi6svtgMyi6NgM8ZsfyUOSir0PBx+Vom+r
wWgrXceCukM/s7F9No6SK8J9FYJL8/kZer96bKfJgpKk0uYyg2k691kNm/tF6g60bY4BMjE9+5JB
ggA3Mr9cAWKujKqbgZ9RQAFvAx5gkzy8naEW4U2yEJao+CAzC1ZEHlFdcm7kWZK0Oc2UI+98wR5Z
OHc08F/s2QeWZECifMDf5GmKfr6f4QjJ+VLAh0P3x0P0Z+yoVpVlK8l379GG3aHIqdz7uQYFeS4a
KWZSC2p5zo8KmsbdMX4hmkFJATpJRctIT/Jpfxln2P4NHyqrRYL7NyoHrhCU8oYwxv625LxuEdlL
5mTaMsRf/LWq3/rtnVjE5jZ85Xc11ctqv2Hw7lG5jMtJo+GziY5j/sR/Wj0g5Yt1T6PrapIMLzxL
AV/VkoCSr/P1PooJ5qzTRo0WmwFnoK0HIRdV82+drkfeRxz1DbHeYBEXMihiSexIM4Q82dvUNPsp
P6R2/2QZg7diz81w3H9NpCa+AaS0kGYOwbhvOIgox5qpmK6Jq9PpiFn8pvn1o6ijvWZNRVbPZOvw
x64oXLRXGrg5PELbei0uSHD4iwkFLyWxsUUe6FsZz3+o9c7jj7VeKGAMqJJjOWOX+hlT2Vzq7YHu
xeSEur1TKXuMlVKk2iyhUahn7bI2hw/X6loh7Elj7TjfY0779caOl4XirYdvmpMGGRvxnKX3mv97
yhWV1rA5DRgHtd/JmULd5G8StY6KVrIi9gP+GYTkQFKuknw6rUGARjuh+XIJtL0WDbSoEuVvU6jl
xiymJ6KgCxTvEa4dE+aw/Jevf8n9GObRh1GPxNpZLXyZ9RVx/Ho/zrSWW9wJK+DbCjiOU8u/85Xb
AvbqvGyVbW24xICxSyqIh0S1YxGrihm+gyyR/gpR34YESmwsip0m72XHNVNaWLhhWXT8ciVDpi7U
VIdpu0kJyXVBwDE6HgfJCtxDeGBnyps/ebBYcb2FbWocGXKcCUOTabcFSzcKjVDmWEo55TM31MQZ
a9qLXTu7qLOMPs06OG8rR1L7ZfMssVbPyq8fY5USHNqad4eP+i5nDabF5X3i/r/9fGuYXP7kUUiI
J6Vjk2calmAladPN7MlT5Xlpaj2JN2o9huLkoPiKe+4oGflPlcC65fv/72CxqtguwgV7V1BfJLX/
aQ85ZYW/a21Eo853eP/ix/QwHKxj1bkqkZ7YoPY2qfP0e28kAFSbBmJ9HkdKf3IdUOJxNPUBKMz9
4KpNvz/YIEJcUCPGJqoYFYkpNQkkQnBFyS4CYcOsr/Rh43rRTaZqGFzLo3YGjCTuMpScHXNUS6VF
XRyKGaXh8beItrJm71Fi8ui4L52UA93R7TtmCMBBqkiQ4As+2qgOjKPcnluY/scskm13UKtC+QN8
Bb31+OPeKruL2ndI4grHP09Ww4rOmRDbXUrD+n4aSXkHDwpY+RFVbLzyKairUIPyggAN8WhKWzPx
kg+B2qJ5Emn9yAU3hYUua8Pgs2tmSALkJKyR9GrmDX/DYG9360izOQAVnrvrrdtmZHN/AOdMX8oH
11eOhepV5kzYX/cTShr4Esgi1TSvLv4+hpJfiwZ1AnmK5vkWc0cIeGZGnQt/vvq9M1fDzamvS95y
EvWMZ0UcKlehiYm/svsJMRwibIQG6fISc1/9CwnCWbnGtY+P8v8FUJXqfshDSAZGPNK3YlYBe7qG
mwIINkXyeztVWRPI1GscTDrgaculOeQ229oTwCfs861LY4g0/oTgua/NLS2Qw1DqAMwikFhdD4rY
fd865DeVBv4P+ysppMi6CCwvCmKLKIZ0lFv5sfpqIKHEhzYXPSsfDl36xGnsea72CtJ6pz8bZvFd
aqkQySsMwUhwUO/tktcWDmXQs3fSGq2A85V0aZy3oXsE85K8yFQHtnikc6YoDFYIHpLys4N0uzTP
bAC3NA+qSI65Rpk5WBonT7KJFzv5ESSyBdT374llc35nNB+vuGMHltyQwboLD7FtYMw1uGJa7+U0
MDeJAd4w+O5K4B+eQYAwNK44esJYpvpnAJsT2ZNqverC5TDNxYM/oU1FPy0Z+PAM+LTGJizj7nlk
UT6e6glUC/ppoj3pQsUiLhJiw9lBIVtzTFDN5Q/2/uf3P1o6YNkHNQtsUkD0puFcecZRyDGVFdww
0oVq5X5GP7hIv4d9SSpqNRq5etfc4Ig7WO6lSrcQqGgPbsqCLT8MuAkh1GugmVScLgf2eX+038RP
jRnQJLt1JCrLZnMlmd9g7kQRdrPQIXGu5grqyJHJairKQncTf5z9IgTJUIAnSLcanLWfp8+XZE5W
QVkwfGU07RsDTCRpaSJ8kKbIU+zHeG/UQpI6ROtygIBcgHEFTSJKVQsn4C33XqUuONZzPBFPHR7Y
mDVz3dk8rZ3qCnX0BWKq2unRwEVUw0sHCqJvEB/jczQCkfoqDXoCKxzoSZa9r35YUoRsfGt+ROQL
vOvji2I2sAr/ujRRpQcGsRcvl+UF04XX58m8NNcYUK8RVmizPicOUBOruIn6LUikeXl5lgd9lSKx
fL2UxXwvojpAFq7PQ6IKtLGMWGiTBbIaSP5Uvu98Xnfxl+i5kNKS0T7/ZIXYpYXZeRFOJHeddB2w
fhYgbGLhsoW+FI2jnI389l2qhskI9gLFNxCS1YQY1FBEVILfJHjsKnh8SXNYoCptuz4C8pVw0f+p
zC27+3cPUhoVqGwvidnzycD+zhav1T/J1VU2YZE78nuZgtqXel27KZtGECw4ujSI3DKad+JAOw6j
lCizXWFqltrZzR5QcsBB0/cZrZKsjLy0AaOCDNVG9cclouEFm7vLgenmYH6nzb0QIsKy8rg0MsX5
rn7D2zXLCNucxaC+JP1BzWU8JjOXuQ+szVxCl5BJp/stazxorfGEIZgXhx3iuSjs5EKfVtrTf3vf
S3EWKco+oqng42Tl5+3aEfdMOevsWvMb4PPVrtxE5iJcmp3puUheOXgSdiVVy5dwOHoARSQ0FgMz
zCdqBzAzWj5RLSynqHzdsgCKUL+Sc2X1sk8xox+kaVA+MCYpbbZSYAQ0oRIgZb+c+O+MnjEpHo0f
aBTVt49PqB4KxKs0VnPrxSw+QoI4RD+7oFcrC4FsDVi/LdRNzOkwWUrSksESt3dJpX7VaETv2mTr
CTkx3nmaie3pDhnTUtDaqU6kok9T0Y+XkjH+EtIY/Y/TuJAjfNKEreXla+8cef4FI788nbYg+Dxa
8HDyRnyzRcyKazSlppRwpGmmchu1KYO9I+zbRtUDJv3yXMv/CiJ7AiNr4p4vDxcJwDqci7JBN1xf
aLGZ0r2uO4MalqjLVsb+OJThHAGal+J7FKVlCH1TAdUIumkmL+ezSeQb8BwmmG+74J2rJ0AZJ4FL
23JJS/IQbO97de5YGPvtl1I/Qo//zC6iPNs+TcVdfSP09DVxaHtinTBOUSRRFB1gOdEGapnvfgxL
0pPbczOPDMhImgCrBXdTxcGo++wrYOxwFQilAWBLVhGRS1l1wWkkCVRJ5SUahbVG/+CXDHVBmS9n
fEpE8KWwhfxk8XDAJiCo7ecImG8iVdh8bG5ZBNJZaPBtp0bUGFjnwNnp5FNXOeYn1EKeqey04o/b
1vhatOgOEtm4DkRCUp3f5Vj6KEyUolIUafreDntLf/+SScrDHUsmE9Rr6D11UkpXiJFFIprIrczG
3HXFtTS3vq/fjt0zn8v5pMXl4LV912ewmraOC1bN1OGaYUSO0ixL0u4do/hpZ6uX1Cm54BpgLmhd
+HHOfVrsJloTZWJmSiw3N8DudNmxt0YfTpfr/1jkzB6SjNCwFJ6AHhIHaahfDu0hmX8NmzSF17f+
vitrHfclW+X1/Y49Bo6cxBcBhX7duUkGcFs7dMQp8f4QzsmQU+103WcxbCdftVzi/5F+X45PSUJw
vvqgRh7sLP6oCXMXP2Bkz8M60J730Rr+xIFPlJqUAZXAEh39S87pDCABKZf576CtLt3gzE1DNxUh
QNCgQbRcJrTR6Xo040FI9li91B0NyX8BWQ+V1I+QnH0wWpRd5A/YPvIqtJn/lmGh+GcTwQZHjcgz
j14nqM6s37lGkZG0Cgj+NV5C4qt+0Zx78asYXXCVlQmhmZJwArqj37n+1iJhLIe2o4mmmW19zLOd
2dnsQhQ4SkD69YL14rVQVsa2nqPABQDVrjmzmcy3gCFxlZSno8quwwX84HV0SNktRAQn2ENkkDQK
MD29XMiHeW2U67AeBUVBesaRI5QjHAeGoxp3fcpFqHBsp8mw4IG8hUiQtZ7ll2PispAcuvhdgdw9
2Nq0DVpiVNPUJAdb1cLdt0t/bFxOSn7QmfaS7XEf5+MR84DHKBzOoauLC6D3/a/HqMf0G8zLUeSZ
XJfIOEdVf4ch70C7ZruiZFddsSVfibFJ/4fgye7r9OklpMd27gbpCCrYijGB4FK3+TtLw3rTV07p
JG165ThlkYjyOaspHqTDOVH7PfsgS9XoGs4jGTj5mxjWLv+zeDcSXJ8nhW9MKxZ2avXRUy9Q70ol
sF/ZKiFbeDEC/PtgGjDJVNo4oNpwPUePQraSJbMX+zFHF3DWGGrp0iCsLehLUaXv5O5NzSzFu7ky
81rpNcWzD2tYboIlc1CXTL5Qx2NWO7/gqTKmKttIznfA5dnm7NcKBA+2FOCcl+C9c3bWSep1+r0W
GDW7u65SeWXzb6xwErzFR1XGNDnnbwpmnWBWFwS565MtX9ybrmImSZw82Rb72zaCz6LFm5WQlnc+
YiUHQgFxrDrVskrP3qU2l4QtjtVAUoRUdq+xSxm3B0fZY5/uH4sqciNdpCpQvaF2Yup3hdNvHfxX
O5RY6bKOqFqudHaDnzgP4dF3BUeEoRwKgyeKv95IsMu0YwxSibcbxlsuPvTXJ1odoP3CtgVdUruw
atFPcFu+JTdp050FV4RacewtVJjXg7E7nYty3HlCT+VnMGOuDLnZkWrwkzm07mFLpetNJ8VHeg4k
R9Vj9TQqcE4b7unMVmjebLAhFAPiXUYZnNhe/Km4OI0DS28Vwuo5GEIw9SqmEWIymqG3EoOp/Ffq
1hQ0VjjUk/aUoWy1AVBzPfli/9MnKzk/x28MTYaUCduScT3moMl4o/ZSqVSh24JvtmDgztCQ9KQh
FtX0DU6iwhpeo1rcJC6wsS1oyXKQpRsSEzkgJTmaBc0SDip5g3WPEZ8zUIvB9BGgpj8mEsWU9J/p
yf6tXAacPKC6R/U4I/f/Slvt7NIClaHYVzhze3wPmtdO1O5qApGD2XbrsgDBdrrTN9C1oWT7nXy8
KBEbHrtrcGXwd5oJRgeD398MXvmu9x0Po1vuqAMB9pz/VroPjeGVTNF09qXD6bREsX/HD20yiIq9
SgLrVxUbjPoiigb+qo2AEVxnjns9n57vxCA9HDCqZRfv8XuvpogTS/nREH8FIzqsmKdhs9afkYA5
YkM2In3ipqZvIUwgdzIam7hprccN/EkOK0APbMfYBM1SsOaNCuh7UQU8A0roxF9WsX65JmeCvaNS
dZNf4OqSNc6TsnaaPOxrxaasOatdT6YTkng7pLRxJmbcjE/+5bps0kLeO1R5WgFSsspPMPb7WvcV
csCIqSTtlLNMNQMgw6io7WmjgbYhdoL85b1Hx55/cxm4DUiEbxZY4dk0FZI3VSUU4VHfrZP0bR9O
gYtNWnZgAvxpt8Epzesh5rQoGrMgo8oGRNKV5m11dnwtCbot8p+fXuB/CMtp3KY1/8D3eQaLmPrB
FhOg/Oe9SuK8J8TdC8ld6/9BIurUbsLAaLKJX2pGtBAtFpKkDOp0mrJgXIoQ+qYEdX/dOT9jKBHK
UZMby4hqaQkNcIWuc1NYJSjD+5OanmcPIoShryVZGWVH48Owc7tRc343b/IgbxfyW9wf3uhV3XLK
rL5W6tP/iBseh2mOWnUwpvWrEpEjKwmoS83gEcic91Cuyf5KmtIoyn8xC6fedTbKfYjAOFlRDLh9
Im0IQmb9indN/YDbYIppIR7lqlNeyrCOj+6uzs4XN2oj6Bs8YXAlfX+XyKPXSCniXw/BXUCZ5zqL
XaEBQuPUqQskpvUYluK/fSp1U2YYrTTPzzCCNyuf2D0AG2sb+YG+orOaoga/ajHqDecnQB6vPSF1
d2GHWSoeufANHFGr9WXtxoJNn6M9PV2uBaRDEeO0VQN0L+QqdXUCyQO40U11lA1C3IwF190XN6W/
qh/lsoCXcXf9bSHcllhqT1ffNGRABs3dkoY5PvuF8O9sWUNOz26hJT5VJmOAIHYjB8dYrd7kXC/l
79htpGCoRlnUd1d2NrgPNq9L4uloHkiIEpntvVKaNdSczzwjKyUySY47Dqw9yXLoRzZ6Y/vyTdyh
n0gXc+tUGn2XzuXsbpgm9Ye5TUDH+IeVzjFN92gi+2GTYaMID4RoDXpFl5+n/D2qGgzZvvNDGbC1
cMzb7BFwr4ecPiJFQnCTw4F5Cb0GLGmg1bJORjL1NiNU4BNqsLJL+O6ue8EILxk2y1ecAs/Ghma8
oAFjnCVipGV2XGRPUcLWjv3XQAjIIBn6FvhTTxW/Vw5rCIsQkLC/6lBemC2KvpDMT0QFIJXIVi29
JmfAkwxslIxsgWXCdLbHyteNWv4CFurnOEXbMQDr3MCqsJMAJfxDzf6QeCmKGbOR9bmpLsGxZ3i3
XhdMfgf3xvbTQIqVywVYJv+8bGh9Z1JULGY9Ghj7jY/aNwLnE5xcpnVjxiVq6aVDNEPYw4Iw9ux7
JTJw/vlkB6rDD8MD9mFDYu0Eqvxy9J9f4u227uWBIUX0hyR/n0RUFkHHJMIGaq0oRevmPoMPMVjn
ZhJYN8MJqnKYYqli72NlsdZllAh88gdWcxnuXv4GIZ+ObYI/oUBK+J9JW7hTH2Ct4I/1RsbG7Z2+
THwsCBbtQIgK33T22vnxQ9Z9J23AGABrs6peV4Ks87a2hNaY7WEO71Ua8oER00tlR/UPQ5CLwaYP
+dy3O9ndUR/l0TXZDA+ytviBj9E9Tyg0kwzsMpyG/p7DhsUp7RNNBmB5R4ODsMILWVyuPb5T3I/u
YcTxO3WNcnIYQDpVzXKdu8iIboYrzXFu6x/7m0NUnsoHTS6lbvWiezhMqY9Z1PXxmZirShXPv/x4
w6EIHi6xJ3+CSG31j2SVeMcxqPSG2GFC1h1Dz++MM/uj+cOfk+LbVDzmcL6aCgRCYIMUw0u8YVxm
twzSS6af2YnGk5NatPDkO2PtymniRb/xmi1GNqQrXL4YoG2ho0E5Zlb88o9ekwA05jCw1MuIHXZd
cpB6VRl3WgMVdKKcuOBWbPBnW3xYfXoZ5SHGdzL3w2wj5yanlWP1dKPPTfzCcH8pijxMoUwao1Y7
mXcwJ5OtWywF3BANwY0yLUQfpbntAyot9V7hkStabgV+u+QgSRMC8uaprUd30lPh5Dv+/f7mDzt+
WFI9p2EaZZLT35YPEIMcFqwZ41D11FCXrZAyL6ebyKT3AfAisAZJfysNyDzo+yQEiVXElMNqO13Z
e3RvytXkW8Zjymxwhk3ZPWiW2S5UeqXM5ha1qbDSnM8jz3DBCcYBpVfqJnLyMQHuXO+e7R2zxAFE
A5fZ+5o5OIYSHQy4dU7IcKXeGegz1dkjmGjlydjJ+kiXCiRB6f16Od7CIffwPBTLzOnwz8xwO+pb
O40rCIMuBQr5RQR0UUa8KtafTO6m/hzKsWq3zAKcGPFVGmnU5QigxeO61irwWZ7lDMuxGGAbmfzg
mIuCG8zXRgNE55WPiMMhlL5dPWEzEafTQZ3XEX7g46hiS16qM3/iunfvjzLj6Mqw2V2IqgEsVkfH
pgts9nJOranaIz993eKxEOqnqiXwjdi/qblKbbIs6ZZ/Wq/WiYFO2Oy0WGzga2dkU435XJww1uhP
e+3XNASDetk0rSGf+ROj1RGb3E3u4uF7gvJPKunzzuQVZuwJ9cNty0ifN0cZeiHfkZLV2lpd1Uxn
byArQ+Njpd2DJgjG0FZ9jsItge3pVH4yNSQXXXr/7kwypgO+bK/R+7ch1PlkwAs7CbDvkk3hIaia
g39Z82hDLGveXdHMBhPYZ5D7IFFtg+/sUqNzSUFcz/VMolCnSXexGEARsJvYqCN325q6fS3sJWpB
YMpTFQYs7TyT5OSnYnmcorgi26QlPuAaJNSsXlkXS7cpsjvIv6rI1t53A5KTWyKzAGcMQavqljnl
cShkFcMaqMTmuYXFVqBWklcrkaYVNQzPFjz920IfNS/2lzVNr/bkgVk8WbCNRZzZQt9PD70mWoJ8
OPIMiRyzqq/QnCrarijDEkzxVNEGh9gYukKCwK0xqwTQkyGphPgenm4HQpk7x3J9cS1yya9c2oiE
hnTs5+hYTdna7GX7cg+0+vesZmN3zMdbwuM2i3N7K0c7yMVxcUm0IE8WSlxYFGJVPGAT+wN2pv+s
G05fLyaaCIK3o4u2u3tasbNe6hsbhwiMGLsZxlE9qUniFtRZo7DOrGAZPSKOyQUa134SoN96RjIb
wj+HBleRQoY7HO+WnFTC741Ovh42nA+v2gk+sbFvQAZaNqrk9jjsfYzFqsDLQu4ZozsTLODknrjI
p8RebtiSkFpS6tEve+kvPGTP2UOSJERoCPIFu2cUwCX0KImYY1C+TbNdDqgcHk6q0ejoq0LU7IEd
oNx9oW5hY9arNSO/xdrvNjlUaVqvqcIoXNFlAdmT8puUdreK1kiIq2vtVdd4CP4m+CfzDpL11l+T
r7IXPGoLvC50cxK6q6XDBe5/3nGxC78m3RZ6xUk6tcViTn0HxbyCxDAyJsusM4bNkkV7oaTHaQka
VNRVjrs/e/08BSORLjsNZSt23alA5FeDZBvwsxlRo9EclRA/+3vOC+7vzNHEz/EaEHCyGHlSy05V
BEaRMhTc3qXb2wujzYa8x127xItvYdB9Dle9mwm3r6zPW/80QvHM4PNJP+Ksxsq8PDcEIw9kOxU2
2imkClkGSuGwqb9Q1D+nw4GB/lA3bruPCE6rZySV/fMZ4zHOm/48RoQfeKxj+wUkTXwn6sjlkMvy
NlXCPeJP77+AzwUWNwuUmdZGjDT2wPz9jiJxmxhgSF4gv07gL0WKx2bIy0j8ofqNmKfw6CJBYFv1
STMtHaPPsprrDFJKQheULVP2c3Tw9T9F9aGSeFr9AlPOIhQ4BzVVCHbbsch73anCc7knKnJ6L2Dk
vxcI1MYrdnsAG2HTcpBG3+E+QwVWNN7sZnoeQJxQtjdol8oYUq2NZXnx6v0CJmtyvYXwc1JWT63Y
F4Lf1j5s+KNUHRIIpazJ6TBQWzLoLw807Dfh4al+FCpwiAL9tk4s9GhFgAKBdKiop+vyMS0QAEYN
R2kf/8lEoKRN72bq4Y/w7DjRS/VWai3j9xz+IEjG+Aacbqu/7JPAi5G5M4fJ0YVQWWyWrxNPw9zM
X6ugwXM26IzrKpRnUdK7xaKcJB/xwqdDBuKb5UndeWw3BBx2VNgsFbKPZUp1oOeBay1CmkEb30V+
ZRBw+9AsbEW6fv9jxgYjvHTsmf1DI/cak05DHZlPp8rU2Mt3ql5bf9ZHtCCUWf+KGrhe1K1lrw05
qLLHGeJWQSplzSAHoO+ezZqdKFTWPiiCsbzjB73jyx6f6HfpiU8mweSWm+sRQBL0Td64c3cE251d
T3vI5XhZ9C41U6sy9syKrfyDFM5yIULkvvSP5uCGVjWKVHmA1r8qpo7BxSloBv0lxwfTdxs9B4p5
9unPm4ehW0Z9cxNAPDr7rLYuZ7GWj5IH3av0gdTNtUdo2samoOkR16IkDUIv0jujy5iwoNCsXsgS
BaAtkICsxXFFl5GpJoFwTT34vu2cmstYw70dZwgq2Uf4WMHfY0KEbyO+xQJW0uuV6AZTQ3pbUlYt
6FcwAVYMQZNGw1hdhKsrVTi0yu7LX+8RPsw19SBH9WbOo/BHDpKzAR+CeA3Z52RMViRPvQtlxJsp
5cZ7YQFH2rVr2HJNr4+S6DySSSTbgSbEyrPCgOOzNpTIO+N0ItjQQb9IXqrR9GkKRXQDLw8tQfRM
mPESG0cIRHxF4sFXVhg/riMR3PtD1le4JB2TVI+twV1D+n5oTqdiAgUEi2fOxdRli6zcx1XgCZ6E
wRmd1zCaOfP1g1dQX349v4ObMd0BYtTu1tngEZJ3MZpkp/V6UTRsBUursC+In/R+nowy2c93pi14
JepA3HtItkQmMngO1KvhScFCxopt09SMAtfkddyiOhvv7Pl1buSLp1s+3urVCQH5mc1nQlhUqGwf
7Bk9/1Q0luPoG9thfnujuA748yFMhSuWvbkYm1pZpHUVNfVZ8fTtVlMBBglgeFiGFhbm/1eQemra
rLUQPaxEjsV7f0aMJrejx7jdyiMM0fZtvWPBPKQrH2fekj8qBf1bWTz/FmhoZPqgnsjDsyFE/tj9
1XTzcQzoH9VC0bFPCCvy8ZQ517m335oFQGwGRApX9E2LoYjQi+5d/tNeERswLwqxuHkULjTIC+Ra
0AVbdIwuzt+F55jY4deJeKreGS+HIjdBOYhIQJeLPF5oVAHmdjc0rZFDX0htxx4Wp8GsfSWbNNEM
GlgcrsqoKcuOZzUuMqriDsZKd68uPDSEJxYMNwdjMtiA/4B7+o7BnFEuBh3Vnk+Sj41V2BsketeT
L5e4ODOIPYE0zMwX+bKK4PuFI85ccUyDYVl+mXtmynApuKWJVofpm7jUxpA4fi/6Ea6xRTiu8RTj
T9Pe0cwHDZ4b4OZUUiLV3GlpIWEIS1R6uOt6xbfm9HoYEHCJRv64+7LP55/cqjZXJlNhe8wIjbFl
gfELmLXibTz+SupkRgcgsgmkGiBOxJw3iMlilTcQ0B88SJZ6MjmzhMuZlUgeqYxN840qvy1r2IHw
IFI6Z1nNirzdxGxDTFNK6Bp4Md84sqr7pawN84Aa97X9nDwnA3ZtRIA2lZeG81hYOChkDpD1hElD
cfp3ziiiS/MDo69ZZjUkEsGPUofOg9bXoHBjYx5MGg7toIqsH8uMfxy+b6TAyhd4tdnp0oxOwYg6
EGG603DOUIwrZdVrMt8jhCQmfhGZNsrC+iXZrcj1hB3lGnZUGaAVlBPL56zrYLAFueugLoYIdbrU
TjIPAK2WsF4gbvO8V1UeKtbUBRQkCefv7+XKSaNDEwuWAFgBncKTNag2y/jgDPrSFX0k1icJRwot
uguiw/hqk//ToGqc1zlpbREZQj/upTKd0+mh/LVTBEU8zdHfUUlYJUO2bzVSbQvfwyFNsT/XyDhf
G571dAq9mOb/yfpmLzamJ6CFRCLQ5Uurh2ZXNzwHPcp4fczxDAVoTsHK65OlA78JXXJl/tU8fNcW
bgSay9L0JyxPcFGpwbhUKCFJrSmjBWYFGCGUMI2PeICqBwriKkVJID+p1njAjn1hTzSQwrztrFQY
cOK2luLhG7XfI0d3Qa6v+ySFfjp3tV2D7e3XKPnv8n40UU3qgHpieuuZnlNfMcQ6qIo3lSJcAnzQ
Rq1b550wtFPv7RPF2w5wPPZhVBl8NZR+dRU53A3KOWpy6pX4C01wrnQalco9HMhuVzbPHBk9t2Jy
p2zoD0HzRBvOH/0LhCOAl25LyvhQXCJkzAJqNLY4/8o5V1B95B6xgkL6xMylhNSaJ6t4ObNkEhRr
iUa0ZPVQt4t0y4XTOuk1KAmucpQce4DDOT96g9zaDNtDuof66ApC3rw+njsmGthj6hOgTraZHQax
By5jgjXs3GBxApjpZIZb0OVW6yqPr1TY1f6Bxc47CN+MsUvqCmpuPw2VRL8ErwPUitD65VVt4vqU
O2d9Hmzj3FvMJt7LvdnpdPpt4bRtkDkqsbEsd+3jtmgl7ZcKVAmqKSKed7ObxMoT1uhkTtBYm4Tc
pANiJCoZmSGeCayZ01pX3mLugK60vLSi2bPNAjm73gQI8J9/a+N5tWQ+Xq0lF7/yNW+a7eR3yBqJ
L0ipULoGI2L0qxXdzmyQzVxVD9gDIxuXoHk6ZLiaZibz/T0SNjHyx2fCiT5gNkMARyuAMJHFT5Dr
Ovz/zJ7r7zXwml5YIkXPvSAGKPJjAbuU5Jf2SdHzcoAzQzhlTFgG+nWKaTDJXU9jUZDTCLPBptXI
7sckrUMpbvObk6A3QqeLvkk0zc4Q9EZw3WQvfpKtLdp7scyNx7cfo1zSDcOQ8qqgPuJy9NByhIYp
VW1PLRHljfcmcogG9oOJYziPkaXvfjkjW/58RirRQowCMyCsuv4Zr+iyDBUy57AFZIgljrzODxcZ
qmWJ6nMkpUB3y1rap1d0DgYL5ySBe6x9KZ5QzMGkGG9i0ZUxIzlog3gcWQU8IPDR1+5I3fG9HxXQ
kZBd9ZeStQwi3RekbrURjjkzumjjfZA9/ttH9DSx/XCsoi2vfLOcwNmxsYMKHQt1L+tzPS8pxxka
LWHm8Ipe4DTf8e35nGQKwHQzDkE8mc8EzEP7USkfFtYY/yD+7msqtvImgllM7zk37GJcple8s0xi
HYfy5bc8QVvo8nVI7zt1QH4YRjtz5dz1BJYYNgXOC2gpHgMYT72oqyoen3PeDftMreAi4cpxYRJA
9j9eCAevfXDpyjI7I9izLE0O2ywGNHIEoF/1s3zoJriemiHFuAIh79ZrwoSzcenjoJR5VtvYHd8v
g/XfzNSfBnIfWXer+r/yRD2lsADPFvzjehP3nuijj84gxLk5EUpsu01mqvywqVV28WITOBcsdGa+
vkSeiytP+QJAiYONMD0dv6duaF2c7xgxA9mJkLHwsGhvFi8Mj/0LMun28+sPpXhAnoOLfG1TX642
V5MkvJw5wzk4SGLi8PzXmE0mwxocMjDbUeD2pup5TdD7GBZq0h2vEiqFC/vCsVo2YnTC0l8Y4Bm4
aiWzkemlLssQCtHYXD1bPHlZRM8NrpF1KOm79K8zsKMhKiWwhyMN8NlJpH9mAIGo8C2cX9eDyy5Z
p4dpjl5mJCEY0vZ7I6TIduPWrIU+oROQRGllU6npjRC5i7RnD+H2fTdumGzeY0xhbmFPyoj0OOzV
3Eep/nkwl67tYc0GuGb0hzpa+1Ax4IGC/8oMfQl0fZKNvoGeeCUo58XYdsHkSsMfDY9Y/tHRRUlK
KJCMPw7YPnjtdqZxmj+4tdOtPMfkrwINbg3NCd6J3FkGrTNuvyQpImbc4zaypBoIlc6XQMv7AS6V
LvUwOIbH7huAhfe4p0Zud2Z4rD1rKd6/gnFFVJr1spts/VgGjlKztlLVRTrcfMFcoDuCtSfyxniN
OVIDNtQb9KjbW6sOq/zQY2WbDrxjefkasLwphaVOqqWGeNgHt2RlC0V+8UAgvUnDw8NrozKpNEPp
lwup2JNHc4jkiQz/JezjjZHqgz7jS0fNRQIymiGFPpkN9wKwBPiUfCyk5D7SGwxpla6yNJY5AKtc
+Ujq6umQn34dXhhDDR5lVHkY05lVvxX48nvtXsmfBC0COsODfnIsPOWS41DMwxQlwg5CKZZGeKcu
nANChNCjJ5Rv1rd51kkAfvzU8bo3B5NnWk/7/BGsBczhCQzjbN81ZTgox0OY7uzdhjHb8xGveyUn
Fir9hJdL2NicQ27D/3sPHSaLwUHH4GY52lqQeqWLXHpA0oPW0I4VsduNR6znxbHwZw5Wt0WUyPcW
Oa4wQp0du3fNhoN6EPoN4YEftyhz3bdnlS0Jfby2SPUi2yrvZQhSIDAVCpxKWn2Wqs6H9IfqA1u2
H0NVwmjzcf/f4Sw1cugi0BZ0HKZ7tGijEApyrUe2E02duVpdnLTqJAZAwQFngoFXdnJnR7Nwj/+N
AH47rBrpbEWTWLyH34yQtwL+oPi5NMtp+hhWrLzm90Q1vMtyzS57qW3kiuAtVpRv5g85wSc6ZRtp
/c1GfYMbvN9jhtatyf9n1mo62tY4QwWm6RIyENixKotCmMAoH1+BGoYhLqAyCcQlKMRYngtjj0gO
wh1oYFFQMVWP/9amMguMr5fle7liAkYqwu63QwtTC+RQm5Nl2hPSl+f0kVw1LmXQXZfnfK9hvZIw
CmhCM+IuKO8Li4Auzoc8eo3TjwgUSOk7bwUWu3hkxrAFg30t7UJYq4ChH0jEx+wyXjXwkk33M3Y1
CCC/mhSRw9JGCe8Cd2hu70Zhk/3ydc7yq8u10OoAwHKjjLNj/2eTo6u75out9uZ8b+9J9XDa/Z5I
TBa3PhARaBnLM7dttZy4CfoqwuogHRgofHesKf2Sl31DB4WGz9CJbj3jK89XPkPb79loGI0YSG0q
qzb2OAPZpKvqw+GZ1LW5sZA+NCPnSu44nF5MLxHvSVhAmAku+KwOzPXdgZ6thmpMwtXXpuvc2/QW
XzZU1Vh7zDJwJSLW06tnySAilB1GMp4r+sB9mCTGYmGlqnlRroqAkMNS8JiIOJx9uLNvxNotICnM
cRGOZhuxtyOa+HjUV6wQBXzF+VwHefCaD2u8Nb88Y4FSyF0HWMnlgLRLGWZGPB4TwoRvmMZJvUpi
GcKZl2c9nnWKcePnL83wjteKh65B+V2EdTbgaIFenSRH7V2Yvd8CUr2XMxt6I1HDa519cDFE6kND
r/FT8d8bhInjmPZ6CBXP3bu7xmXWCrl+LYKkYQD/fwBPkXI+vbo+0Goplv2hwoyuveEPyL1kqDM/
x5p3kgbZzNhZNetE3egHir8bwmKsL3lsEs8Yq70Hj3dSUkJiYTelZT1fe9MK7ocLriJxgVsmq789
2nNMZc9SRk16F0y8DDbEZntQAYEM4uhFCUXZFxSgceKkQdiOL09zIxOT12fzHFykM1mZUtyCjs+0
APo3CluCVP2IjqiLbB0uX6c7/xW3MCo906Mp2/A90lTGt5mgDsE/pPRWYdRclwmPv/KHyvzDwsDl
VEF5ZhpZXKgQD5E+iT0Y6rfntcrnpZivV8b7nQ4NYUzxrHZ3qyY/iOx57iDSEOBihpywl1swQ5FV
evUs4EKoG08ZwAGqGrRpfMBKYejglkvcIKlJ/plkKkoyiuZ5RIIU8Y6vnzKAD794wggQs3ERXlbt
KhPCqWzmGYcXCf4AVHacBdGFI6P6MqVRSDOioXo6EDBZlW8DUSazlFmorFNq9Z0ZloJ3pY1kgb5f
C9uf4YrbKObQtcq21doiKqKoTCOqSqgQoA2+xZnKuZfUbwZZ5T5Y9JrFb0IADEDkTU0iQtszJQHG
qasiU7wV78tz+pIVyiojyWAeCf3C1dOZbjCvtB9hyEmVNvivD3ioS9j4G+nJ38UTWlbTvaWkHiqR
WvI6vItB7tx2nd2CLbpsdmRWGFQNB+epO91sRcoSsk4NyB5K/Gvhtuv75pSW0Bf1+9CbHrJT6RxB
nOV9AdN8NtdDQzDT+cQn9x3bbvEZyj7b7IBDoW+CzrCWh1NesHDSWfaHqE5T/6BCgjqnOTnApQ2D
bzd6BQXRd0M/2bve23mvhXpsnr8XhRRkhzsXsXyCdCNS7K1XVwQqHd9+tiZ+fMvIiAAyLFxmp2IJ
2dSAPAGMMgcgFQUH9PXUvw7J+XqHyXUgDls6YPa/ytL7SV0uf5byGbuLhoQHFX5ZdsQRgAHR/t9A
wmCmaLE6b0adWMOMOa5h+zNvMUAS5UPA9S8QAF+xOo5ZyCqEIvFPV6vG8o297+wgeF8QCcZgiUtM
50oZI1pUedlaqPdUzbK2y6t8kW2YRDCtqg4BCHKtwpRfaRSAQcpKcpqtWbZlaeMf1tb+yeE01xBn
OVKpdD72l9jq+F7um0LSIgrP9mX8PJF1kTFgdZ7T+FP50FXBDQu5HwhfXDnzlOWPCeZQcXMCQYga
Gf5XoStEOUeQgfBIeJSux6FFUjC4LFuNWdhGKapnRh58JDzCutnAwR+2rliq59t8n/kDnk8+OOk9
FZZX3kEJYfoI0+RMRXyhVgX4uAuYJKAFeA4rXsQHUHObji6QNPPy9t51L39N1UKeR+I2LHUyUQTz
fxNZi9O/CRuJwsv1WYnXbo1XX9wSBIiDt0nLBt9h+3EBFJt22s0a4JjVQJRNEFYNPju3rAJK7C8x
M17KFRMhb4Ia3E6ZG1zltp/yfriFHqgDbYNCEu21a/aksG1h7sEHTFIDTZn3VkLzfqOuVRRb6j8d
T0ivUm1TGd2DRYEHKZJ6lHSUEHZE+l/B/h8Kwmkh+dIK/avz5Rl/3hxzcy3mNo6ZjzFqcYHIMHIB
eHb48sS6DgMXYtFd0KcueyKlHkjUUm3RhnZiwdOt43D696GNn9ESNa1uOaMtrJCAGEruNp1aJQ/a
QzZifaghrXzZfuPLW9S+Oi0ZuTVultqVDLjqvNzdHw+cLL5qDvbLa3brJp/WtiUdReijhUZoNaGh
Wxa/3JKiyq8VzruYOR9vgTXMYx5/bpg+iQ5m5FkCztLFFa8l/PnT5/3jNVlxdCEazUxVotwfITxr
pdN7cGOgWMkr7L51G1FOaXhdaytjBWn+N6TGZrQvJHCb6yf2u8R6MYRNXj0jEv9cg4ssL9Wlia8g
B13OgQkQWXG/rbfByuLz1Lxw4HJZw/2KZYflvh5jya+e/00Wg4euIFNGbPr907QAC3YSNctV4TWC
VtQqhiLyW+L33MnMCE4/3EN3J5bEOWBrfkRJQZd3TlNht1+Segt4m2jOCw+o7IisaCknbG5NrDDX
12r30jD4XVuhxJ4FWXR/PmZySNGn5wZE+mkK4nASNQ3QHQ1/zdmihOHmrfJe4WD3R2sjGJooVgWn
ca85YufpbpiJKiOJRlQ0oS61V0QeuJdQfQSnK/9jVtk6zCe3Lwn8cfIAO19SqNjdTv3ZNNhee+ll
q5dvr8l/TuyluKrMMH9ik3NemQa2ME5+2t4nFzTdPhRn3D2H+WXSDHWW39jRlEStMOeXdld53BOx
xzzq6iJ8AmNgHObZCPJPOdOoy/kYc4HXks7V52TRBW8wBdvl11uYT/IS8rNedirhmFGye0NI25Xu
c5RTiaQ2vXluIE2osQGNraJ4jvA9gnGAMTxxtMbiHUTkKDrM81iBB0L31z4TX3azvceb7dhVICNL
v7+5lZk4+S4ATqBpxiLL+OUK/8RK2LLnDwBUlliXb/0WtJ/eAD0/aj5x4QFGgGWXj50KpGzZ3eK2
b27mlmWJzbE6cYV9AMiLy1SKScLs/Se5VfY7IgLhLIVsSBZbxgI+qjdpwnieBSkCGs4rlccsyngZ
5FRX1y9icec9pDgTCpKcHa4rsZUfVDeLOMIKZrzve7W2iBa9tNzU5+MDgH+jxuX2L+RPmLLiU2oc
xOrtm0TFsTsbDiU90ZR3umhLsYuBZs5GgON2bEnLTD/nmkVdA34rRk3jqeFNrKwVYb15pK9EBb73
I1SpJvDiZVX1t6u9j0gyfSs1SjLIYNLp+qGIZixW0hlQwOQ+ZphKN8qS8aXMjljp8CPmNK4sFuTz
XG6wZAqREejFBmqEtwD+qGpuHYjmKuDU6RC5XhOY51Tk+HvHR8B/62gSY7ueA40PwgiBWes4l2Hk
8zh18t/FSxWPNCL7SCECZc8hm0MV2rJAaROBfh2RoAcHmMjIz8UDcOL5zs3vy4lecJuNIo2+/Gxj
wgKN6F9nXQGCVfJ8W5F4rSoc+/DsWLl8bF0DzbOXyUlZJNwVm7SXztYgat1PNLmJXz/Jq+t3SWzR
z2qNGpUZYdhoRjEZ3+NjjdNOlCE/cgUR5nPy8HsUFcEtxn/ihBayXr+h8Z1MDjVN1/iWkMpWz53m
G3d63RkxKHh14qUGBvmSf6QHd3C8PQ4M40NdyFhcFp0ZmnDJyO4SJsxbaIeMj5HANRdZjngLjFzW
E3ZYH2plgIpG3CnthV5dKDjyJhUse8nEAR8g+SDamRzjQ6Y9uEpbwxhZRj1exp/BM7beiapkjlEw
75ZnjZn0VriJLf3Le/FQEXAbWbSAiQ+JVlr8cN9xO/TnpsCR6w49QVwcjA6Qcc0vsQZBJBCsq55a
9Bj7oX4ut8i3XOgNw+Wbb6wx7oGo+tA1Uz8Ae8e99yK0HAWU2Q5W97+ZmmGAKKBKXus2YIRVVxys
FILIgozNO7DxdDQF4Sc5lRDxn8StYff9ctcIzqIAjeR/WpCqGA+xjLIWRk6LwwxaW71UTGvyXiCn
eTmOthbVyZnwamosIKXkg3DQJxkNvW9v6GIbMrccuSeVqsuuIClidQLfVMe4PHuntKOmOW5bo4tu
6PzW0UkNFxJaaTwnu9bm5LAW8HSmjRPH4bjSEDGNL9RYMfmWRYEDWlC9yzi2KHG8HHlw/ZtMYWEH
k1b39r1IBmCJnTGFtdoZOdNrcEVU1sHk/+S6ZAK0RFQuAT+PxmHYyk+naaiX5UZuzxFEJvHSPT2J
TJQtHSBr5rZy5FG/eiYL0mp7LDXyXMy5uF0dkhMWyb2UNVeDCoyJ7h/XI92Np04gXM9WmiRZ3gES
frIOFiTSO1fspPFkKm0h6trY6DOIz/5Uw59kbwDLttv+V6RhkCi9Fe6R5cVAmqJpgoBJg0rSVxTn
inkCemhGJ0rM4htjYMvCyBIEXjET7G4Z5R9malMsfPBEJKymns5jmDsqapT8/g5sXg470CbQWzA0
HZ+e7LF/0S6tXpVRVJF9wwgqtkBf9RsnidKHZKye5Sg956+82O7UBtrux9cr/GW/8oAVwtgAr6s4
Ohxnkjjpds7UzW10qBkKk+/YTD1YOCp2Pju1Gu8GswEwyNOr0HOkRR3SPXxyywd9i7P1EfC3fHUC
RktaE0s93pw8G4BmnT6ee+vwXAGQkjZ/P5whTghJmg0p173kZilLBZgt5m9UVQzrbei2rOSXeB94
puvOjEdM+hU5Y+El6k/jQmwQGsPcbQynQgKXb56K+ss3Gqv12pGNaVymC7wUgDI3lL+Ys5g2aAuQ
Srf/v+HauUxitq+vIavuOJp//met17s9Z55pqfzjRiPUHFMf986eE+/XHG7cbh34DW02COgUDhnh
0C5qWtDGag02pjQgVHo5LqKxhOZ7ydokkG4JzRbFOP/1qzBQCKY+/b4bjxn483Mefd//jorbXFL5
ugerzpmeXU818nZXypl7FT4WVs1f50tPEa4XohnYzR1MabA6DEeDjKl6Nla6txB2C93AnhGBLABL
RzHukyqtMGSYyiQSmv1r2aoD9uB2tuV6k/ujtIIvo1Sz2zFpHSztgc8oSrgZrbrQ3lVbW1c5V5LP
CxV4YMD+zmrOxsdGwZOWeyq8U8zJLAHFHH46kLqrE0B6tJXTXDkN77aaN0Nbe+76SI6/X/UZ7YVi
Ecm/1i+h4RHtz6cM8WG4jy99Sk/lJW2heCFfyRgnGtyAPlGD5UGiPJ1/6rmgDq6vkYajP22gTO4W
BfrF6uubutqm/5J3juBbgfrT4ePaWb777tC+zieJkclezM3wMqfKs+fmBlFMGacfrsGdNHu+bE42
5PFGciSkCwXG74CfvlcYuHBCBYi2qHE8PNAnw6Oyw0dszVJinIMauqVu/rN2Y45ReqwRcteiHT/k
M3nXkd7a+xPj1wtgWN141TZbnZV8QT8K3Tnmqyb9+5GnCQatLBBLQ8vaNqxcyWkaM48Dmizo8Co9
qNg+SN+l1Yx0GpiFjlHDLAg7Gf5wfTr8J/a2T0xo3zy47Q2ywu7BrMzlIJaShlpjtsq7mgNdeq22
I7mLVNEyPdXAUIfKWlZe8UiZQ+Ga+Gi09ybUHY2AKfkPkEHQQ9dUxXg4j/yfE0kVrJDSKcei1Chj
jN/Dp5ulZ1y7i8Hc1g3OOSJM8Kd15vjXmVfn24PXHYxGq128UA3CaZA1tAygCesNHzfgpZsnElCH
CdQio+D8y9aRRMAZKeousJollVT6GKBmqQr77fNvKXcQ3KOHdXYYsN0kfe0CO0jCuXCZaLaYgL/4
DChlcJqhV9p0pxrd/qNq/2zgOZqJCMoS53eFMPEdRNSMpzqtBiJq+aGvBGXtrcKhxa4dxq7miksy
7Z0R8r0dQeUE3xD06pCBpth69rmHNDtDu+pRUH4kLtWuRkCbMFJ+820mxc1AI90fk44Y37NWuYWG
XBQiRvNzi2S8f6sik4GTfkYEtMm4RI4i3x682rp+F0pv3MaVBf3RXTwh7BcbJ/u3mUIBW1/mphbk
L5UB/7/Sxw1Q01lQEr8vfjLAGFaep204pJUKs6gUA+g2oCGJ2Nic9TuHV+DwM1dIsCyZ+YEvbouC
GhmGp8zBFVxGMKbErX0wNpd2oywE7b6optNFQKof4AJ2KO5MlkEzwuoF3ugJQgdK8MBEIfurbGL3
JVIqi75NwEu1KXaCexpBS66dd/I2S4AijZ/F5RikyDRmV5y9pXBxEvufZ3E6ZpVobE6+DIevTag6
zz40TC88mYUUQAKYWlgw+E/kWskVsQjMfL9udgqV+5LGLo/9n+SNvPWIYhdJiwOYYAKYn3FJeoPn
m7amYzo/f7B/6G5MEeRiHx7jwrwDyXjdaNX+99T1mMZqvSxXLqXPEJoi/rHMf1BpDkFQRrD2y8E3
8elVLAaZCPBZlpNJ2r36pJtOk6uCPyn37uD6qvIOnUGfd79/RdXPWmpnGRScxHYhDG57NqpQ7JsN
l3QajHaAYogPxTk/flbcLxBzmWpqawZlLDcRaoJfb7L1PytA269OOu2Fw7XShPRbQDG8ESfwZhM7
GO3Cca1lzZgia3ucmgek3lP5DVcxMl+4+SlUwI7D6blZ9ZUSCb3SMFk2vVHRmOTDiBhSLHYezrjL
s7FRdOFkDbxltEt5D1A+kYcl+COVLm3/Vm1JiN8XeRmB6gMsC1MAxFwgHDh+agXkDZpMb4le2uQY
e0lg5CJ4eeDfjagnzSIVe72eJjvLEMrIvsYfmDVpLgxG6U6+G0v5xtiBJizzJXW6i4VuAYhTJ2MV
ED66X61Wxn7M3+cX3XFzKuiocIpwDIaEk2DwvtqlHq2qa39neHmXOFktLgmblBbEdezQzhYP2ZET
K21AZHIUd6GRrUOr/Sp/lFTGlF56D61d30Xf8FMxHtlE3y0ZsNRjqevuKgvGjMVs1slKFCtKtmDr
RSpMNHdpftmYCbM/HMrY926Yzfr4dFZao/QG1iFick9zHMcQ7hW2f4xwf5+DQ6R97fxs767t3qW+
zYOkRgWZQgFfKkboGu91ZchuB2wF/G7xCd6YevMIoz4OZBH42MqnTWtB2KmIx/5WqgudVj1Dxhd9
L6Q3UdSHKIdGTNC3gJuAaj9e6on1kfaBmQUgYUWEERD2Oo3Feij1FlcqBqVHbcwRnEmRLPPaNEX3
JC4YpmrhkRl1kcriiGYVihrT7GB0wTymIzLvm0xFwUsCHErf386HaKsJX/s74YAR9BjdJcRNJFG0
ZUy5uw46bZWaNOhQTr/IVQGeIj5iTiUoFgE5jvHjdoHsW67Fmu00hGys4RopdQgBYHhHZxE7GkNm
0Drn/JDbfmnUo59GshH27SwNSOs0Qs8q8aWpnMgFnAQx3BD1hogKCgE1BWlcWsQFh2hBnhtRlVSM
OPvB5WFXvORlhLRBY7Uqca0PzwH7p6KZCXyWk+htJmZusKuZotXij7TC9PheVVOTALdltWtOljgk
3Rjunv5/tSsU5cMzQ85czgWiNRewSSqM+75LQ1l8Xpd0dIm2c8x9M6LE01H3PLaKYixpotlcjwG8
iDqE/JFVY3CTMcbcAqML9O7yMhiwJzzh7/nYe6D8sB9XTfKayjE8k5KGcvnx7O5jxzN9LIzdVb2Z
cMH//iVIkrujHllGTzbMi130/JqTgw1ijd+4s7Ncb5bjvotxd/g0U7KW7/bDhVHMLFTFYlxmZD39
xNEAAm+pyBqsS2YFdQMHt1lDq5dO/nb8kh/vQvOGut9BxFDhqK1dO/wUizVf/MRtgGB+saICULRF
cxcyMp1wpOsq+/7TgqwjJyuFIzW1zzyp7CQ3l2VyIRUSYU/B5m+MKeZW9699G2CxaFTPJZjTpOzu
mCyqfCFTdbp7/wbSs+H7e8N2+L5L+4AwCQbyH3EYCB7uEE26gG782EdlCtwUGwLssP3Zfp8hENjF
3hkgKbbX8MLdQGyNtmqEeWtXWrQsaiKZa0IsiVTgxJr4tx0kKnlmC+kqjTXAwY3e42srW49Dum8s
ni3+rKTGWSb+hVTTVwR9nQB5DUZKYnHhhGJOYcPZc/tAFZsfJE3PoLICXSYjuli0Rj38cFwU4em2
bT2q+7wugz8MIcWXoTfBytU//UL+fgPJqzSqTblu0PXxrFxpNU/tU125dRvNpZ6bpGZGVtbr4ddb
QsBmZ/MNIUEA5GEtNgb0da2xROu4nZDt1svnhXpRawTZcXW8/x0HYLOttj5IqTAm2jBwPzwLEYdW
i8hXV9bRjGn7LduiGzIAQvKZBquEtH2PrO7HwljxZPgyTkbuef773E3ubjH9yawKxKlDQbI7RwXm
YV5cYnH0EtL/2ZYrCyaYNPxi168FXA9ll6IjWptU9BL/+C8iEEAb7Qw0ES4O+9DYnYqko9V/pjs+
w3wo9yLam/kNvYDIKnzKnrKFoPvPSscdWPkO6DOKQMhGUmnj//rErJFKHmd3FkXarVp3jhCKKT95
Z8Hx/0cNNvkDhN3JG9mlXuyCTF3yFr6BGUCVeHBa3VKtDcozS9ILkQpgJVLVPCnkM0nGRF7y8TNT
PsdHUWIz8WVjBVbwTmW+cnSHzUY7rdbdDMY81WuiLspGdRlEXtO41+/e2E2KZhPk6YV0S2JVI/Gu
wD56p5DbwOWLg7VZSyn0nI0Lh/faoyLz7Gcj2uIpNGQDi0kpsz8AlZ0xo3YMXDoFSNSfjBEpwECD
y9BuBaAsz2SugDJNvip7RXLcGnqVm4B3bloyJ7ulhoQc8lrKuRQAjRtN6o4BB/FH+dEuI1q2SxRr
K9KglT83Jv5HM4POz6jd0M1PiJ9EgiCnoXuSUTxfmDiDNbK+5xLSu1Zg+p31oMnRsykwJY+Z1Ad/
CcPiDBpCxN+AfXOKrvFFQfeF0Y+5o8xzA+g5AXgP87bJVI99QGnfaFDL6u6pTVkX77cUsIdk/GHX
yxV+q1QC7rEcmCUudgtRNUhXy5LQck2h+KRtOozVD79NeqFL2WYaEsFnCdwMOB0I/UgJc8gj8HS7
3AYDdWhO75V04SNYNxFzl92BMcEiuYAPMNf22AS60068DNO6JXoUz4BLXoimXvCRMnpg9YnajaLT
OB+iMUsiPwKOIo8MgvV6wdPoT1KbKpi+HJIWanE2UtHoFonwjxzzrl4/F/1kOHg0t7YC5nBXrvsg
xHWfnuFjbn5woCHka6Q72QA7OE3Uwg9v1veruQKBxyxuEKhk3tfpTQ8J3rnFfs5ZWEUAl4/8O4bu
ng5/0TKDfbCQ9Zf0j0ORIGvnVGDbmTzMRLLQmpuEpAzmseBkCmeUmeZ4CU0FT6/RzhaxRganZAd7
MXnVgnUSvsBufihvnyJCwDBj50vUSb1EByTbp1ffc9kQOExAtEticfSa9fuGp1mI2sGHgIdh5QyO
nuAHtNyFKro3PesJjLjrtQTwM/XuTkEG/Kib3vuD+3WbZEt7XDK1imbuSf+MMqu3ylgoETb/ouVw
rEDC/1ZDwLpbPbfKNFRXFE335oNrPUHzoueKyB+m6sEaFp8bAAafaeA98GdNA9nkHwF0wV9OEPJx
IxHiF6eCKyXMfik++Ys6+J+PrxojzbMTHsE6Btba7MluxrOh40DTFA4mZ58tvFMyjmfs5tNUC91i
QPhTEEazKgkzg4kmcpvJ7H3VZGSwYYrnHwjvbs6cZxxvjuHiMMMNEC/75Xhq7HWzsxezHZSiia6O
4NXarRmW1lo+mmP1c5kJX4OQ1oKQ28Bw66pS/Fu2uw17UJpnA5m8Utr/cdgLKn3HXabQAKg2EcsB
DthpJYucUfm24LPZZveiEmmH/St4PswVIgAis08Dy7rX+AjuhVA0KZ8i6fqetdt6fZ+cyvzbrx8e
QFX0acu/ukOHJ5Q23tP45xdEln+C0vWw6jdFkqqTH00PhuQQgriHrViMxf3pMp2sayghztBfaqSR
0bRYduovvxuWlrg9TQW3KXKhNtMafg3F/CsEWtM/loNVE01Spt9+IFi3H7LDojfNh8yokF9cz5xf
T54Tuj/opp8g7QB0LQq5VKa9CB3ZZG2emuhMzX8ucosp4TA2KkU4sR+XvJuNI3lIf8k9ScmEGInE
H3nEudEXO+i5tG4biFk6ODWl87u0PwMQYZZw2s9hI5Uk/BMpv7ppQ2wjgw6o1MNbv+vparxmKQ6j
7qi//o0hzBYTYJk7tdHifkNgiXfkJbdaEt5CuP8WJH7EWjStdE8ylB0YbFLbRuImJ0ne8SFJzhtf
8y/15ju/6TRQsyzd+1if25+Sh18leRUA1pS49yASShDGYE6lVYX8RIOlb7j0pW0Q0zqwiVjxbNEe
tp/PkJt6nuo9RuLdmpca9djq3xV+RIZJRZOgvzh3sWHw0qKV8P1yhtWZhPQRICrgkPZzU0Pu6Zpy
dcnV5S3tllYONN58U86PMzyTLr4r2qcI3hbH1xIXRElNfxM/nzEJlP95DNv0B3Xg8BAbk+IPeFt3
D9z1ZfvDWF+IaZDPEdvszE51/O8iQT8Wf6l2gI/twgcedOak3Kn1y8QbfyAigVfnBJWcsVDgurWH
/jV5fupLu+WuaYj3y4aYoJkyXGKL4RJKbzDUl0/QOZKbhY76YvmJvNdeX+TWI7n+WN8mlO9QUZo4
E5dLDnRWtylo90XBsj7AHaAXSdZ6Zsc8F8IVv1BKjbEvQ8idmx56H20mAPgbqrz0V5ve9wMa6TTi
crg3oLbqGuEzXQA5dyKBzl2ldgih+yejkj17LrPzrQ4JzN0OQryO8qlx0/n+ga8BLdNw0SmxBhem
iwAZGXI7HuPyeYRYy9tqVT3n8DV8+zk3OkQjaLR4tIcNBN0WvGCPdJ3dFY3tqpzOvqEyuTru50xe
Zp1dXvpcabl4m0O61IRI4opGXzQG4aRALAkmhsWqfZz3iWgf8KurS7HzRHeggUAo0+6dcdLYEEZm
HzuS+Wx1ruHSKcO4AC3GI3CNHJwCsdMZdO5S4ROn1ZJ5zC72Vm5e5dRTGtUJpPZqklEBAXGDTQ1S
hIvezJKcsB+SFTUD9scLHuzbcDnmGte+LE1JXYZ8A7soGYCz6I4xXPctrVFqgEwh4PxU6k3CcDDr
ihy8v8iWh9vAlDZM05ODatbmsKBNcFtOvRVZgloVUgYaEFYWfy8E5Y7mE3MMiF8SNAUhMCLXeJgb
Alz584mTYk4lN21aqFJWWgvONUn2bseyumQpDk5kTPl2Si5i82cxbUF6V504Fr2ZonGxpqCw4Ija
As3gdJXTVlqh1Pos+P/UVCjFNqNe50N6QnaACsGZ3hPXZ4UDmCvE13e0gzg5bQUlx6POeMSfniOG
vDEaEx39sDbm+Y29tXG5UsUiHSfAIw/ugv0RpiUV76dX39YBb1Vmoo/abbJsf/OTGIDEv4lpAAL8
kLVcKJaQsCxMa/9a0Il5POjB9gsG6GtuxiddppbV0IvFlqd5uNuyUNSwxsGorODIi8Sw93JLixPO
PW7Uym+zTFGG+9WZV4GjaY3Z/xO9WqP3wETjQuYDdhLcD9jAv6e0XnHSrjRbYaaYjooOV52g1csD
O2AJGa8CAb7qcQQmQWTExZeiQT0lPcoXDdNgphFFvlFeJdNbs8IgRp6M6GRreApI2L1mAhLKZG8e
L1uf2TqdO/akZi4usqn1j+vfSz7llPAh9Uh+UtB3KWXRol3Eg2LWjcP9jk4GLl6wbxfK4dZCfQ24
/a/lDIkNkKL9yqFML1mGv+2NWx6i/ZhSwHayM3FZWizzcT4avkpWbd+ObD3IaibQWpsWdEkPjSXi
istDVt8BmUBBmYL53sGg/D5662WRgyMdpeQsrIBp8YbfXFIolEBve85cXOMVO5kyv9BBwaNRN6I7
VDbDA5h4VtYOJwfuFqT7+6g/31ZI8FHYi6SVOwBh8lA0jeCamnLOAHZkat2yQeaCNsUz0Y9Ee13n
Q+Gj/j9eentd+DLxG68vCjNLH5hVpZMs1+MrdrD/Z3283VAM2hADL5qkBGfYzQ2hWHQ8rPrMOqE6
GjtqM4mOBxfUIGA7gL3RWE2tnaxUvra1yX2tVyalZtYogHQeCIxMBeMw6/eWpn+r6/hHHOpg59q8
b4MNDW4ntki+bgdXIB9dQT9ENmsEMUhomuply3SOqEIpyRQlNLrNVxSwZvo8LnfpU/yFwoCcWeNq
fb9w60aR16w3E9PpR+R6D1xnBeHSsu2uUYGLY2OVvStTHRJmQcITzZ9OZTwnl91UoJ7MAx1bOHVS
83UeYSvNn3HxcGxTo+miU9jEW3vE82clhuHnHbDHvUQmwlITozjO1KKWygUeRmDPsNtkn1Go922s
nlXptqIiRN3JXcG4Sc0TCPZ5clLrX5lb44aJPhyTjf88W13KyZUu0d1W8+TfGwZhflROH3kr2Oao
Oda35DLtZACAyFW+QDuSDapwr0ba2zCQxbSRr1iHjQrQxeBraS6btFHKT29/7UcixRFDC1JXlCCV
PXmCJaBcGDXPgeEuxReEIcuTrSL4qPbfk1D8A3dLQ0ClytKHntoK+vVMa7rLtdVannK+WSWOrPWx
JS5W6rHZ2it/Vpamctgf3VUPbFfc1abN0RzhKrIta0WS6H9Wq+qRfEsGJJjbesqqjHtNR2H7MPjF
qt+V/Xb9+XwV26F75gejUULXraVdISwjttl4EvuMiY2kH8xnq2+kM3r6XkWhE7M+qc1PPzURd+lo
s1S3pac4DuoJZUGytSmIAV/9v3pYc0GjUgJpiXDhmovI/WYwKIrXYJNj9bFXOGpBRVusOzwnShey
X3ZOqQpi102rqQkPQfmMnIMTsB4Hc+G7ymLKs1ADhPNNdtOaFgNxKmLlYgN1Saoa+sOUqqiWJO3I
LjgY8XqC9gdst1cCaI6CSfR2l144GnGM7NxNSoip8Zr4HeV+YMWUZahFDVw5YfPrpo/TVYMUz/wz
ptZ1PU+72OK0duPn33Q64OnY0EnSxysT8wLAJ3wNrMhWXRco9G9GKYaI8qK8wDaj3khZyI+UF3/w
2kfzZ7Y9t9o4YvXxO7qw6npfDtaGN4FUp37Y5WKtHdXVyuSt+saW/GfwstNq62Df6HBfWa4YCFsc
rzTgmR/GEt5lce0ankFc5QBT6qTwzbU8O9Z5knX5VvgxQ5Zouyx1NDnBwRcqpELVLl6jn26UGMqE
6KoGsM4lBb6JXwS4nh/r64jnQ9oZeJIY+TpAVSmb6o4SAShUfue1YXfbDLQbLOIdY3AmveYIT7Wy
00dm2wC3UjRJcJ3mQmkcyDNv+AAigeDIdGTjAxKgEwDGcA4SxG5qkHugJ1YtlxIr9DEnTECJ5t4A
y4tILs9GtBrB2pxEfj9E7fPQ2mtAU0K3EzIDbEccz63j5VBzY6SaXpmHC6ViHKb2/lOuEtLkrhhP
f/k3tWIcdIMkzb48lAFBw1cChBenIqbxkTLojaVbfGj8SrG+zKL/NzTmbI5BlP9lLva0Ow+Jjniu
6jQRNlcOm1kQ6yLXcuXlJ7t+wGjkp7LzRS7Osu+L310HDwYPL1gsGGvpp5fb5wb5XuS9rUNDa1xw
kYkoYL+A8rfLl6QNOzrUOBvlYXd00pRTAdSv6ZPXK9OxzyVS/UofX0ABfNnWTBY+QF+1CO18LHbR
qobfo48+KFm0+1iFqQUM/7N32tuh8frismCDMtfmv834o2+VlXtCD7r0J31wY1S1Crd7+ExZZvFu
ZiozbuftF+3iZrINjrSgZcC1BYKSWLmYTjnrrVpdpXLhds3KhYlkVqRijKvmf3SV5mdkS4VaxcDF
Hc12Z19medqCM6Zcd6YHhA3RsUNhAbBrH2sF0qTWSAnp2WJWQD/6rjIrYu2DirtmRRBsPm5mPIt/
WWeyOtk7PL9PRAOgoQhOVbWIPG8sRNRqXTQ6yftkNhIyHYOqPo5wmaQROowSfviU/u7RKHjY50yI
2m4YeijyOtYCyAkwROo254xw1YMDyypS19IZYmTcJszBDHRqeTgFBH0oqUXQA0RXNv0QuTTNrX6k
eJqcG9ycNwOFvHmDG2EA5JCGa5u7fakSWbw8/r8bSUiNJ/l+H3LEyZBl7vN4mlCBFg2O1hrB1o+O
4oDgWyw+kBLzP59P9iMbt2c/LS4Us7/pclymeKNC2UTi1REZzoWUnF2uPJBD40IjmdPRDkx5N4tn
shDMZsdNvOrvygrQRsb/0khBeUmc89EUUXMlUNIuljcUk88hFDC/f1a4IINHZssTo2WPNqZV8moG
z5vFSwBWFd850AUpehIEuYO6iBylHERDYXa7htzXsbos6ghLxBI3IfcgUIUwtW88oHidmToX+Hbt
kQnSH4yPzwqX6upna8Z9fNZNwA776at1EvYWpUSsvvLj3rYFccWBFKJ5dOIAZjYeKmZrDqtSCywF
vlHbkg2IcG0RFyWg8euK+rPz5uTCDauP3ypCyeTiNQICPXTn3EQJe1ht0IrswdS/QxNyYpRel7Mh
7m/Fn414i+Y1cfdmK0QqLWtzESlClENr1NF/8Tl0ekkLRN9FtXI3B5v3T0hocoGN0ghZkIL7PO1W
SJ07x137nbAT/rwi9G3WNFaAlk4K5bSU/2dprvCGyULF5uuBstoy+EHYmFYY5tv/H9rvfUAPqrfZ
F1B8nxS7POuLEBnBPfrZPghVg5VfDYsu0NoMHcv8F8kXDPsDjAeA0D16wfgm2Xo7GJ/TqEYAxpCS
fax5BSydn87pXyUcDGPRUugL+bw/y7KZz51AgZNgqpnDHI40o9OvMLgODaScvNo4h8UG8bFWHmsd
TMOsEWcFEzUFUPhzmUHJkAJXY4lfFHku025khLnGuBZ3JtEp6x6n9WbGk1Wwn+RGiPksPx9sRBjw
ZndQwa08/NcAL2XC95b8vo9wFXaB7Axl2GceZg+23//f4mdsaX6cq7Cv+FDQVvhUFS/TASVf3AsH
oq86Nz4SLaiSHHGA8F2QUUfxMMz3A0iVRcM7T+u0WFgea0ciz9U03+lrZOnqSunLCkqrLw5x1PXu
7cN8taYVIGL++K49EaWlsAODFrETxVkrTq8yZXiej6Kn6R8e9fYOIGLPgES3Ks21ZJxIzbNNuRGm
Rr4HvELLhY2D6P/syWsQTS4KFh4XYKMDLMFL9HEBtF93++A1IY0Ju6tdea6uh/yKKq6fSRml3ECH
HTWi+htutMBs3LDvm5WiGDIt1lON34yd2zNG6cIaPpPXHOtiesD4S5MDBitVSZgjbRoKWhZ+ReVh
R+UniCRmzAUg+DtTnxPPFnIJ/pY+3AeDS4AxelqabRT6Uw/dyRSx49DIAQlnvDR2web/npyjpy/T
SB9RxQMGevtRkjDRnxtPhmMalI8KCxYUiiWBA8K/ugglQL1IbL6lBr2HMd7RWcKFbpX6LMdXgwrD
N+7rwh+YjSOUOq1//6nt/yIwYtKxMP9EAhpaw1eex1k7S5qFsxTO9rFaH3QF9/64rKhBoOAehFH+
nFYzZxD9hk9BxwB5BoIUcWFp2itQyJ7H1Nr00e6kBB+pJZtvQQswXjhG/fhKmzg+byQBZPHi3YDR
2lrsb49nLb7EC8oJ/072ghMgc0anburCyaJ6mzPh4pUxF/Knm+3OvTPrLKpdG5DpX9srexjqE27w
HhEB/8LF1M7ljYU8x1UvTYJ8C0M34VEiaMCq4a6Ug1wpiunLwZv6BrMLC/d21i15opFZrj5UTPbM
hCM/AV/OzDAN705dDJY8uGoYxD7z/+jyaRDwOUIjJabrOUkimZKXtNpLYnWrleI8CsCIXe8igKOy
L2Jg38lg98wDka1jFHrBfhzzK4BLcsz7l6MOBheW3wzGsGn5K6Glt0lAUFmwODfNAp2APi36d9nM
r4plm/vKV6hDFh+p1gz4UohZGbGKvdGIFal80+ZoEzv0N3Ft9SdTQDYdBnJ9Wge2XvJlwIUwK5/F
1mAfkwLLfaPoTly4QPnqeHkh9SeNPw2Z7MGgrBwahucGLIcTP8UL/pl4PWefi7H3BZ1sNfFNN1vv
6dNwJHXK0PTPCkS7ATQD5ogXZ2mj/7qtr9p06+B9Kzp3dsMBJA0IszuFqmdn0yyUI0vXTQazgGz5
cljJhh+RDesXlhd9FRDA3cV8DjNOAV0CtS8rSloMRplXgCL3WnBsRNTj6AzTF29NByOWSGLlVzAs
wJEjIHrMz4XKsTH3M+P/NhoI3HCpCwb/bK0MO+Th+t83CX0JFhKTOPALQlT91NQx6/vtzxPUx9sg
5i2y8kRE7zSSCeSXVag6cLOALTqEZJM3N4iuErqCL8Pagpj7bmZuIPQAGlP8j4w9MQb0yzArwNcD
d2OL/wbxlwlXFvjmB+ElA0Lr3GMYHEWaRW1eHMxh0KsfZzL33PYU4m+/Ig1egYPqNdZAVON/ji90
mWRNwe+SoXVXca16KHlKJAHeydPktnjugQ46yo9biecTS2PnWYkpUKhc0OgJVvvTG30+VthF6dL5
siaFL3mi+MLx4/b5/KjDFbmQ1EcpiTQ30GUnVyZw7ornzatpYg+rA7HqinfaJMnMMbtc84F64a2Y
YnH4AUv5BiB0iRtkX+w0SEH6pfeQZXvnMwdq2/jfhECPqWaHITXnpPII+MU4sZa6cAApqRR9hgXt
ATacF/wgYy2Sgi3SaE6lifFR9GBR3tY16mIJfyb3DHmjjjBHfq6HD+kd8Ke/EamaGiO1Im6OtGaL
3WIkuscoXRfBm1QvPhPWQ6nrVRO0IjbA1N1HL1z7KGi8Ita373fz66eqLRGjOhGNW4+hCMrM71aD
TGaTNoLjbbmRX8dtXRg5TPcukGYJ5i8GwtZdvE8NdfLzGmHaMlcqlmq4YWGdzpalGGMn20rG/5+n
zyVH9ocb82WwYuP2PxEjDPn5eZkcaTRZFJQwTmRgNr3R+twZklbY/d2dDJT0M1q9TQwuIykUUlPB
dv2jb3OFrtGEtPKtLbnMW1/0Gp+42zIUYYwB0uFjLvp91xsuZqvB+fUCvyQiaS1JVqevqXOri3Cf
lpDD6LBqC6fTTAap7GgYgf6EhtbQmSoFiB0tZX5pnDy0jXgjuGzRcbBlA3Dks5uQ8hn0LUsy2YTw
YfYTOzkn5FdaGkFG0luU7GfwEeJJBaH1h4avCyeNg+8BM3wVBbAdiYC+0K3zpsPvHR8wVUstxglO
YLbzhIvwKa1eC5bMQLC0G8Er13ASmumQbJAtWvI+af+OdBESlvOIL/gcfjQhwOzSJr0GlOUVydmm
JBccgbuSEzoQzE9n6nFbNlsi7URjSi0ik00med0NO5/L481V4kRJc7vqyLphzjHkPCScPg2PAfkL
9O7+Lk+3IUt9oxm0vSMqU1N82wMnlM+T6/dXHJD93gRhmDeEdqemY4L5gnGZsLLk/o4ZQnfddj5B
+ST2A3V8Mwe1NECMWBemuxoD7ZkegQTFEFaBRMhcaZazZ8F8v38W4cznQTOt3m2uisz11EV26zUr
M3S9OEL5pUQU14n1s2mziJoU/eWcUEmyW01KrRClHdh+aSIhMmcX4FexrmeV1WiKV7OiWYd/PX12
OzWvoK1xuqC9aQm7TgRR+2O6CIFb6fFPP+Hp3ygTUIzx/k/SN0I7rw4RcjMD86V9RLRYj7fyTgI+
Z9NVRCHbVbLJTVmLAav9XlLSVOxNYnV5F1KwiJ00hKrTLjqrJ1J7SXW7NwqmIzfYeTBsQMcr/g4/
en+XMUVAbyGWFOYo07rN/MrTHp7kM0e2iXhpG3ZNx98jEwuyuaSPWUdAwtfYXoKV/NAhtHF1ICYF
yTk1wIEGPCVaJxSPqGZU0sJJduVm5FwJeK/8X3Ztqa2q5pG7EFZy4afW5eXxKBrDgNK+mnbOZn0q
Pf0mI0OLV0F0RXm4STK3SEt3BpH2GmuCtVBfJQUjSqQrtOqWYGWa5GnJMnEy8dsn8yiXchIs48jD
mcJxiHQrbfz8FWJe5JKPGfE1BdM0ilbVsXm1bF8tuNUNQRD5s50750NBoeCtGeYpUiVZC9uXdJ4v
1GOafuHHnrwbX1NCZ6pkxf31hYgnefcWiqjEK1oNOrys6fgJg9VQeoRyUKW/iHyVevPTFj+JUY/F
PPpvVGb/eEgE7db6DA7bqYASn1QF1B5JzdJcfhtZGQo1Sru5NODHhLtGss29GDRnAfEZYkUbI97w
A3xTgTHJQiplpAXKCs9vUkW9gwpBPzD0spcIHgE8xPYm6r4Fg/0/+dXpMduaMZVDTv27xaNk1K4F
GMOnSUUw6Pd+MIuPpL3SzH+L5XpIwOmPLaMFkpsqDO2V/9cIpGLxZ7i1pULjzXdUk3/YjUTJ1wtP
kkIYwZUsfQhRejlLX/9N6hS6cKU5kKCodzaV0CtswdXRO0u1ZtCWAregfGCZ27razHPnrVaT0Nfn
0JQNyVgD85Etj6GE7Jvm7Ap9tPkBDx3HNy4stWNUdPmuAceRkyYjRe5sY3M+LpxdsjbJ85oFvR8R
DOtJkFSrDIBKheO6Zo1W+jRjTs71c3BYx3/xjtJxcfJdhqWUer/CI1mFOvaVMLv4YBw9jmbQsBMF
Uofh8jFEputoDqT8jFaBQ50IoByy9oH2DShfrJshMLHJB2so0lH7lXYTHL1Fh+zG07YE/z9N4VK3
9ivmCs0LqOSmmHJ0YvNjvdfjs+rTd2sDN0edsdlcwH+dkJ3qzvWlq5tWz2wxQwlPrgcM8n9WYKIs
j8xW6NWo5jgoucRsgyzw49xDTxEaYVc9Xri5IvijJsGWoZWiFrBR9Wz9FVoaGyD2Gp6Csgql6zzP
1AbN8hhVw7N/elONtgwtasELELX88TRd5EhuZrRbooArsCkU2gWZdFzopqV/nFXfucGAa8es8NA7
w+Jax9gDPEshpSRv34pF8j5kzm0Gd4TrvuqcC7kMiR87JI7bur4PF8YAq+43WKUCVLbLjBQgmwe8
5SUD+R7eoL8wLe4FVoGBW1mMHwBP7+u8qCdr4X5Agvm8hASZKQbGESXnJp+4L1mXk38S6IWGf3Xg
azCLwlvZp12bx7Og9g/rzBNcafnO2gWTOxl/HbEOcZ7EuX0EgydGhn2zkTQeEeqYzlro25UBEyU9
b6mI/fKm8ASP42gtKUPppBpneSvJNvTOU3E1dPrCY2VzBLDSGX8GwAdTQ9FM0nWKGa7HLs2sQE5K
FAiOUJNi51l9H7/5dgw5EsKh/PSrDlNXZfNIHSaySxwkRw7Xb7j5RwpYpwwR/vJ6ALYEFzauR9VS
uaOVFzOYOpJ+xTEyYx0n4MKFqmno9fNNjUMQ0YxmXsupa4zOGazg9l0GknbEUcRETJBDrbWRzRuI
jM0kLA5nqpdYsxBkxiwZkvmfwC+dNfc4u1Isr1GxCgkPSZcvVakFPyDFmzDKWt0ODiqiOLpLlFOE
rWfU3z754/ZKJjt9IMFTxR9/pFi5TbZ0AElXmdtCaT/5ZBsqyYZfCAkfG3Ztdw9P57eh/gxWapgB
fCAE3cPH4NEhyRla51mB6F3n/UJlPitTa9MvIys7x5Cqz1r6U4NVyc8TnXzNPTa5br21Ifwwrfgr
Rl5gr0HeJRYmMfItTEnjgptEuDGfApPijBzrgeMYCJTJ7Dul1qQJS6YSrpzZjseL+pzSO4VpQbon
zfqoZjGp2aO83HqmR20J9Su0viwVun6J7n7W09yvyk2dwNybbfaavePykUpXKgEBGMKZOJ9LCJvP
oWb0No1B//eV/WhpbtDh+wNRejgl3CRGCqdODP9Bbuycn1BtVIvoFpOZz1cxh1pf1Ls16CkXo8jP
RKDKzknKUPqWx5OE9bAdy0s42LcI8McIX/lU2BVXl9yzM70+06+E9Z1e8aAFXMZ6Phg9ERJZOLGJ
akmkYwpGunMrQrBjgLoEMUaJ8OeW00thOCVLoDG10Ke3acYvhdzBkNg3UsLDqzrlUM2dk59pEkUH
ZPKjQDC3mmrgJJhGOAatJaPgz0YsX/8tbECK/CqWwSsPwHMUW+1lveYQFRRWrAa2K7i5VjU05qd8
6Zt8yMGzqWarv8zXBVBid7PgFGYzhWVNKsUU6Eu1TqJvThjGhA3WpZzbkgZyB68i9/Z1+u6lAijH
LyaWDiKclX9tFpJBSXLGyAK8BtOlDw40Ydkv2pTbqNiZRc6E+cmJuNPq6y2LsyUla9zpTzGaq9Kg
KRCHTi+G+ATyazkKDyqeG9vpjlJvrBdCdALXt6Z16dmaQzJnbJ2+CR5v80q0+ObpdABmouv9Xjol
OuDxw3cJoGahWAH5FGvOAjF9dc7IG4RWV0ZIc7DPtr/tUx4TQFRM7odjtgYoOgKBBEwnuwAZP+rP
evSR67cxV5u6CofyKIARzEBr/9LYiVSonGsbLsZGagRHiOxJmaTATq/gmwLMKyWQDkwfidsgH/ly
4hLRE3GTtzebLs/9nFxOBWQzNd/5uVM1KdE0Ao5fgZHNSVrMfJHJt8Baxr5VUrfoF5bqZU+dusgv
eQrC5m/tHMT8n4BLO6B+ckJsGUxlRKNzb7s4eC4aJvQrI9zCKEEohFHV/XKDENRHmb7TZxLT1qas
n2Ekqp5oZOCWASQq03ofXzK40ZJtuBh1n7WTglkepw6Bucz/1mg6pbQT4GFjoc5s0N9cm5XKGa0U
wjLY98iRMe0EL5GZgRaSFT4L78s2B31H9gsZ0blzb+I5NxvpPNu3KqsS0qCqPMtBjZ7XuCKdLwoq
vAwFKVXryw7HMWOEfFvSTka8dS9Py0CgKWsc7gR3OHrtIT3gS+LD1giychd9R1LNhQzGLVFodKVE
VjWlQx/CoLCNqP27dx0CB8U/JE+kbzLiVjDpSWyzidnmUR5BiU9PrBZOQ38nNfqADQCE/Wmw3RZd
v/rtKoxS6Do5IMdqeZ5ZjigUaI7DDByZSM3OO9TY1igwnzbssOylEoV9hRbwMXYOf6G4i2JER3f1
S0Qo6W+H6O8i+GClwrFcGsyosP+nZUjIfl2yhBBhg0vyc2J5dgnXqpNm/+G2Frp7CpmUSI7rdtjY
XX1/ceZxGwnP4gkConhs1rLjrLvEOzhAWTnN+rIu40LkBwytEussXr+Lsua696lmocEodoDntnft
OSSTlEhAZQfHq1JJrxmcCC7tgPcoAL6kfCG3oDSMx7ZNOHu754e7wUmCw+/0r0Kwulq5YnmmMyQg
HF6xGk0ohX1AqQ3iRhMzIirWdjNdvGs4FdsZDJAwDcEoKbBzMU+G3NmhI2XPRX9wBweaqpbIxtnk
rCuOvMGZ2HPjdxv/7NAE4iXNb6VtenQ59YBFbY0FUCFOXzlQvfQp7vxdabwrqD5z465UGyGjq7Uz
O14Ty2kWrMBJBk55Wc/C5UTw/q7jgmI5VSMVg9XLumR5CXuJfwRyE36dYS/KDD0Eyez1MmMwvGca
DxQp6IvU3fDmm12ad68iz9FTamDY+IBVTR659Bx4KBC9FA+swPaufzFEZhOzTekK3fEdrtuyyR5c
Ns+TajK2OzYQ1iU2aGZzZM/Q5M+vp5Ww1N3owv8Kuqh2ijBuMn3DhF5t2tGDAh/94uukg82Lohml
sh9f4McrMqUUX0SjRuFlz+3sDIOU5emR/uxGu4Gp1KLu8FC4bJlIoia2rc6053CvljrhCobGhpQL
vRBn4Hgbe1ahHKACOoPVaj/O8ZKNjNlGguh54LrwY6+bjB6MyuM3sups2Wa+5du20EhoAOiFhd0t
etSt0dYXWVfkD88qi+hd0ibdxBNEEIGo/PEGZUcjAa+EH2R7Qio8dKVWroqO2UTH6p4XviHC+YeC
5xiStTHJJFAa7IYUUDGv7gSklLrw417So5IuA2UxkgyoyDZig5RqSQ5tLrSjCYTFugz/0NFJjG8l
RiohLMXTk159RU1BRadAXOid3SYFmRKgYwSYotBGX/zA4hPN6SaheaTURAaKOnUODZNPP/TxGwTZ
Ns25lcWGooWYZxCP3vIQWfNPREYkIHF+uCIRwa6p9oyGVrbP9xCdZ1XqIHMN0yK8V1BvIgsepRuo
WHlUempf/xzhwyTNLLHAB/UCsxhvwBrWM6Ze40jBJ14/vVc9XM4bnC33XNxpsbQ1Efv/dtrb+xr3
KhH+xs7SdAJtY0iE/w9kihKo42YkisJYoMrhi+9db9LBp3f408Cpq1Far/PRqv2q0AMpGwUS+jrL
Qlqj84TPk+J6QDBpaSyT5CtunAgbjxcQfkZgBG3xj0/OI0CkQbjo7IKWTaLsW7ziLIlXbDjtRgtU
RR59isdTMg8u0mlNYPYt1XZiV3eWgR5dfm2Kp6l6UP4s8/rVDNzph3PvWVm+W5qJOfEKu8WPKLd8
g/r+iPiXSg9+wtnqjVaXcwL/5lTLSuB5mGTYLAEBelrmMeaf1rpjXxJF89FKlE6Qr7JYuePprxtf
nqJoURLRaNZHlTcf0JYd4ZOo/kA0sc0Hj7CpvYuOoPIZIiIp+yh43FMvAKM/Ni8YGgasNqRe/cI2
1Wb3w93empZ8Vv0+x/x9Ybj5W6DSpdIwMQqjZrDU9WarQvlqGQ2NPOtau8HToPCcoE2WVwSgobfk
M2hnVUGuvWtXIh4pyuUo7sIUbaeOPO+ns9f4rdorz82KZ1MK4AC3ftZb26UvtV1iptvObKQ0joGG
bJXFp0XF/AN1941HgDlJBuKukvUyZ5oG+y9HG+WocPKawEWsBK7qmjmVHquVyNhamwf0D9Ds1N9p
XI4v170Asm3mxJIodo5zPEOhtpuJ5ZMfyfo3+s9DJabEdpd91GRetKqqlxHeTxP2SahqVLCnz/VP
m4B/c7T6bOLRCCib140cHF045OfL9TEjpOAq8OgXmoKq6Gy9l5NhSt5FTyaIwubHmP87ZAIm0jcJ
BAS66wTZ3oPFYqTjWu6SHQBXf5lS/Vhmq7xGE/13zImmDG1MVmt530lRmb0Dw2AlxZzbVYfOfzMC
RAfmuEKJa2S7EvdUa79LoFbnRKParW9vgO/m8+8TySzCNHtz71Way8xPEk7hqPikubiQqJJ5Zlet
OinxxmXu4yEnLaLe1+kgvLXuJSeszIJQsg3AIWd+Yj447NtHbUqLNXuuRb5ru5lOjRhUFXKqthJ/
sPs1RJBAThjedF9I7ixVyOBR+zGnj/8qdH02yo5sh3wUysI7E4za/MU2PwYHMEHCJNkajMk1HpF4
PpfzuTQU7K9U5LehoQiRHhOpxmR/A62ItSI/w5NRDOG+fiu+jWAEPunJGlcw0n2yT9eBVltbCTxC
MRr6BzcG9k7+ydOG7YyKr+QqiTiZZBcF7lj3LB7j/b8AfCKIl2IpmOSqD7S5bkX1vawEVh7U4bWX
01ZEIlkMKocevFZJE/H1eJr2uJdvJfFCXrX1GJWq2hiRf2rQfUPoDpPydRQBuQj3LZgJwWTr2uqR
ZKjuD4ERPeOzu56ZaB1Fzs+2/T50ZFbl7dp0fTjoVL+Uw+cZErqASOQa3BXmjooFqcvrv2RQvwEZ
LuBeunxlN8WuW/EyKHXj6aiZoIMxPjDYyJdYj7q0g9/PSWCipWTIzxjf3X3LlBFUASLfNt8pDI2/
slxeGu0UhBJ9OLfk9EofAoUuMHxFnro9JcdwHf0ub7x+ZDIKzT/vo3MfOlHy2W3LVFNiPFTOZqax
+NbXazjEe3hyNXKypax9JAY8wv0CW5mNRDNA05oT7AilFYP6R2tFpwwHWDdPsn5i9VsVX1kB41z+
CcQbtr9zvgJz4J0anSBUF5CXRwUq7xbpI9rMX0vqSIMQFwM2Ggcu3AXUL4IjsiGzalUaQN73J8j4
G/kTrRzZ20XX/YhoVv7B4ZdPKzQAGzZp/ItiAzgQ6x8VBAuZKKi1cXaqc037YV51IBR1NYFLvUTS
XYrNR0MSpjQKXq2tNhvjOGrdNmxmN7kDbTb4G8Oaw/u0RxY10EnF8OC5zv0uh7QKLlvJg1mtDNfh
BvWI8HdGB6gckl18X2KlDnEIpmFB6xVwNc2F2r5m7pTDnZw+lM1QpJ+9cmCubqlLKfQQULBmImxL
T2jcpssFlwgjsIYV3dMvuM94AtjhhLJgQezLvmaVaGqhyO2lKuUgqbEDTn9hLUR/XSc46nZdwxLb
2AO4rBKnaLFhvtlHlbZgELcwFs9R8S4hbJbknggxrpXUGdNeFrMvRUvBoRRvQx+Z4LT+CDcelI5w
x28K9nODqBYYKYNqJZT12ZSYaLkBzOZ9ntF3U4YhoSb06Sx4NN9JqTYQiZar51GMuX6fCNdSZH2M
aIEu6zNbDaV1z9hJDeslSEqtfgvqNJLj7UmS/fqDGT6+ebtPYx1A8Lt6+WwwdI7dDRnclI7b1Lyb
1xoKgqyQ8q6i3Z0ITrCYvw+CgKTaxQ/B+G2q6eDCTFrIrdWlxlWqqnkGOrrsi5OlXXeMaHaw3jax
vfSkJRaqvo4y7d7Ocx9r0uKXnq8nXhD1j0kuYXPOixw9rAURX4VLxT4lZiMo4uM7SyN/HzUDId0k
j/7j52gMv2InJPxzir9zfI9FMvPWWWmfyMgoutM7nmwGh3SKcckesmXF8NshCzS41exA3U7x2MLj
A332ld//gVCy39uBcctro0KQd+zOpqSBBpKJEHy9Ew5LSbhgIYh8H3Q6ZVZIdo/qN4f4RtZJbDdI
aUuWJSS2fxXjbrk+MOmeGXQef6C0/pwB1odWc7zYbl+gSw2kk85VCF/YHikNQpwbtmZObxVTQ+dM
GIaqdV7nev+xlq0X9omZUxKzziZbOnkeQs6cNVavGhXZgSEyLgr5IL48wAPdZg3LpM/Ul/aP1Idj
t9bU6K/p1NTFGLqyxuD08rXpSYLpkbVw7ES69c7PO/c/N3cOVRJ+mYL/32KcXZQ1ISl1a+WdBw5W
ReZdzjV2XrsB9kDRJ1Z5bdScqt2OiDJ0JaU+181wu1Y+nR+NNzEcGd+8KOumXNCQ3PgJomqa5Vst
7OmMb/5ZFLrPP6Uw9a0tm1rxiIzcayDAYsOjJWlj4CRs8d8OOTTJogyntXDvAnfbT1OiFZKyGGYP
hZQdSoNmnjbRg47ycGU7XuPVgTAmxOa1tf6bDKMj2rfzRhrfZ24/i8GfYkiwbzTUI79wPwhOlma6
e1z3owdA9tg7CrkxMYjXBp+Y1PkHsR2jJH9YCom5mJFL6ro3sLYrio24sG79y9AF/CCjnQnFAQxi
BXtAr6C1VhFwIxO6KP+QzMGz7sCb43Upn2uMelEZ6P88edNcrD2NjthZHa6aFYfpRWy1fyEEkwLf
8g0mqBYrlkJyMYsD462IptWLDDNoHZCkhtJpuP3VBvyd33Ln4gBdxqN6svF+JnmALSjh05qF6JRO
uzfPI9mf7ikS4rBMBZz1oaypwnTfiZCyhYzj/9QYgS22TA0gp5kwkmTfBblPS17CpPIEJdNO475F
a2i1ogHt3LXi8JMsU030Z00UxGwdbE89+8pCuMFHIHZ6QL3bRuAxTjtpRSItmhOkhstQ2onA6sid
oS7bod+VkpV9c5NLdzouEQ+0ThwgYeEvHLUrcIk5nSzdX30jvPhMJPWFKU9XICt8ylH21GDR56RN
zfxpnvREQzYo9Lk/pUVmcEl9vhuM7SyyBwtToJyUcs8RxvzXq30eET0AQngIuSW9PaIMsQGKRRXM
aEMrfOmlIYEtFGqR24o+aI0ywTFb7OStgvMhCEOxA0AbGuo+Ywr8y5Fv2p4gFOk+ExgRc+CHLXxk
8EGy+h4mDdKqMyJKdhvYkD3r4EQVHJz6AIa7rCJzq/Y5FCgdsQwilCzoSm007b8ORGQ38ah4GGkw
ZRWvhLoltuBleinGU5f77HibviHYduQTD3r89Rqq6yckk90knULRJkeHd/xtsx5vTymIRSlqxb6k
0JLfG/3OklaMtLVzUdZecR0B1VeKGGQW+zz2jYJMXLHGc3I2nEuFPnT5XoLKH1p7f6syyymxw2kn
/2yoww0T3biaLN4QVDcseDkQ7GuIQcLSkAVBCSr4F+1xuzEcUklK4uphX7Lhm3n4oCyW+FEqHttj
rYg+YHE1gGp4onOXjPHVrReCXNPNe9wtIOTTvZ+A5R+tGJQ3mXH2zDb7OM7PcBP833Abqz9daYIo
9CpzZR6ghuHjV6VhxO/+Y0saRCfFXMzZizrpca5fI+JRBgyop0PebR4jUaevN73JNQyq90sT4udf
9yZzGIRWzn7I4/VTRVCaJrxaZsnaxC/B9BU9dL69Ccs4rhK/sTAKSg+UTn9t2oYDPsKAe/mWBMtb
vTpogl7nrnwhn1fodMWQmtCd8UclsB9FHBjoOF0gcOgFlGHTGMZDq5OWWmTq1Fdy6qtz9S/2fBG4
2sRPACVpNmRl48NFe6socpZoG5UTYfRIejAKqbVUQgV6mnY86Y4kiJ1HC4/KMKLIn9kn8PxYgT0y
0tLZ1+cLvtr/RM9HKxytSu7nE0Z4V78dWkqzwCLKdQBNACipODLd/ZnFqcu3W4+wcYEsuQtBFhb3
CpPb5wPxxLA3QCPiISQwkQet9eTfm+rNL5v17pvRJQnkpDtu7vZYTzpeC3pEiWgfvIG7HjDrMyKE
iQLz0SDXjngG5CVg9/h38uc24C8pQc0M9CR/vlg8NRHVYVUU2XM56y0zdeTMUfNiQMdSXe1Ep2uS
HabFzUeBWw4thDzWZKqBwEAxlBkh/4zQPLCM3BjKVpdRBF71BBNlJQlpGG5QbgUqrMbNCpWykKSP
jvhNIOCSCgWXTRgUfh+pnFyorjR0Yyg7OZopfuM6BrajIZBRxteBo+UbVmrhiKGf0rArYA5X6FD2
wJ/DjQfqFCnH2lnnhjAIedhSrUCPVbEEnMB9BcG1T3wtVodHKA859bONdDfX1hB82BcRrUjeVTZk
DinuzRckowNs2dTM/2a3CE0sPBJYKnyB7DDwXqKXY1kD/4OamtZkeLMXgTyfiEAQwfXxXrK+V07W
A7fKKeMsN23QqAs5P/0/S/J85ClfWbHUXmpVrgJmWTwMlFrQjUUdgvEGLOBeS3vrXuaDiyFaodhA
2SRvBqIkaX7HSKj4o7BHaaqQ3A5DM2ZMNGSpSn3ERMVlzN+CUU05lZGDibZUYU50uxvAsVhCBR0W
81i6PeRig7rYPTZNralaWOX79k6SXRC+wiDOlbm+8FeJe+R2+OlF0pc4JTlIqMpHXkH2HdKYm/OF
Niq1VtqzhVzbiD/Ix0IQJzyhw2BNT3hgWiItcvZecbJtcl8Drh4KhbFX5pdB+Hd9iiF1Ad1hpPJL
t8PU94aLL+IoffE4ok+twMBIqu7mTHT9mI+c8i0vQNSHf6GtHlZbwd/mcOmGOHrrOt5wuY4ErP9O
Wt7tfWxCk1ipSEshCaRWhkZT98b1HoZQ1fYTNaCy+Jnsyl9/G9nMh4wFlk9UPe3DE4rU7n8j13oL
wF7YVcsSpwO/nyHYMbNgnI3LspBeTSG9vFFYQHMWmlljfQi9WVqle4HnCyDcR/cLNTQWH76BAvEU
lmnlp4GeYNokPLxg5rKaK0/0sJht08b77/V72ELIcc3gOdVhSx2loBeKtLv4zb1mqOPoHsOqWKzm
DNEgUmcjXbccFqjxTylc/UPqSr9oRvgtjQ/ahK6jhwvxS1mjbN4NbvtRbqVivmk4FE81qKOnKw9B
H/GzpmJuULb/+WuTITKMW/LzPpV98J2PSPJ+d77Cia2N6eVEzSwlPpmwzASX6UsTcRgiHsEoiGSW
IEB/ju/Yp1Iw9wnWTt4Ke7ieSLqLi3znwFeQNDshxlCaedJbUQkYkucM0Kwj8H7ouu8AcV2+8AQG
N8LNk/WiT41xfYJ48zQ0rQSDZjoZMZcs0UifY9Z5TJlfD6zTySKeCebVHcfpcqTT6CxIwOHxOv4B
AL6VMj2cvPKhf4ngv1ZDXXNlUWQYk55U/Mke0+YH297t82SpmyfdWH1CsqA1GKtYXKMjIPrajeOI
ndFtuceBGwFCuV8oTCG2VajW8wt3XBdJLE8HNvupc6A8ptozi3SS/UTBh7GAzc/xBFnKerigokm4
R6+mRhiposTupshtT9JdkyEI6e4IjwcqtU8I1DCO7bYu9QuK4s+Zi4u2peG+UGLy+YMOswUSTJwi
MkZOzedAJW1+WgXRLWKFvgrOhILAR8UuQnt6SR6pUlpuZVv0kFDEwWOOEmdcYT5Ni9tW1DXgLeHg
KCoC/OazJpSI3HqqOptHCBBEBq07dOoH+JVrBRApZhW/k2Ixu2qUfRNQEZPst75yIqrlwgKxX2AW
/k3HzDDDipkbKbjz93n0gfHwM49fA5ROUCkfhAU12Y32abUiKFOA1gLi4ky3oBXdY7edbkkQQVbt
Isy1v9AsKYLETS6lfTEL7w4zNjOPDgC0W0pLZqTI0Gt+1FjDuR/2bkZWXamSG3cAEMfp/1tvL6sT
YPnzVqBFJnw2NbhbqxzmcOTBR9q49JnZ5xepNxV7hP0AKKiRPyMU0HZUhC2qUn8TlOGh1XAKrsh/
GEz502ii2Yow6ts3AK2c6fHpH35zTJANHZFiCnQ/XO9AzdTUNCs27BdyVirP5+V8aCPd3Fp8S9OO
6n7NlRKR84tAgPNu+mqMMdwJy97b7i8xq+Agxx0dxPcZnasOInpt6nJqGY7lq71wHMstQLC/I3/w
cLHH1bT0bQOnQuf7K998AKsh0igJPoThw91zNsZ8/WvnDHr2r42qM4ens6rfyJqcSpnX1bgK8L/1
Lm2o+iE8mI1hRjSksDuQbtybcgdqcBkQ5S5KWvahD3WVma7t/8iN2rNwtqGVMt0oPgzrPwCK7a6D
bSJpXF1LP2Kkuyje3hHgB0pCFGzMn3Y8zFJSoK2BICedIcu9uScjUb6vDdYEkGYg7dOM4a/rKfgi
C0mkges8i3MbTEMsW/tosd+TB5f6mHybObIbIQ6swoJXkq8gfiIqhQ2CUlYKx0/JrnlGHh9OzYAd
DvKVwXBXHmY3F4eyuSyBLv2p9Edeugtoy8P6hCB3b5xlRqM68e0qfi0AtU1Zl/+9IEC9nQsRAl+Z
tY7S6medK743NfQfsCBMiUu36hWmbEVPYqlwyVHNpK9QWY1AQ1bLHLGg9r1W1fm750IMK9xSlO/h
qUA8gQs2pmGT92/dGVH8ENeGhBKN8P4uREqle7x6vSpu++1XL03SzfUzY6vwIdhoQzQoy8uOPL83
TCXcQwYCzcmy/W0SYuYCoEwrmhI3vvpWuPF+j/4uuaYevJ6GNsBVuAbuxB/KnyglT/9bERe1R2O5
nhkpNXlLahVvY6q3Zk5Z3KpBDrFIKpKo/bQvRx4hDRjrS79M/8iZ4QFDbr8g1612NGlgP5MdFFyZ
IgHQWZsfrUy2dUiwsE1Ytho0WRiFkIxpTkCnOIWCd0OvJ5omXKz87fnYbEQVz2Jcg6HNMzrA+8et
+15HMmyST0qWIMlyBFVDtHspz25Z1TtzBU3yCFGr4ODxA5sZu5d/BeZ4HPY2EEAL4tkQ7mB8jKN3
xi+bu8Mph7K1mXqG4YFTUFGb1R+ckp7p25+OXFIUoMu8Csdo7ILrcZz1OQhKVtJrBKU+7vgHt0kx
VSCwo6Q8f1/2/m3TgOrUkXmv0DKTey65QnQDp8VBN85DEjtaWcZ1PE7SQU5037wLeOPjC61JNech
WcyLcHDl/4CBEZ1YALt3tb/DW+MhZ8OhjguT5l96+SnMCAaMqrKOoFxpVJeV0HFdK4WN02gBX+zR
lsVvjs2XAeXdUHAb2OMBoBqY1q/Gd6OyjXF+Qh54eePCstmwTUp0vTijy8xDmLzOw07VH1Ktiy8O
CnQrsjY2AglvB/+x9TyqhRmHAqaWBokdJaGsI09FDkrXtlrX9tpPfSwO/RKx+wpcKWUk2VJgv9pm
Nj+YXYeWCHYmwkkfWqhUxINrHBTjv/wQrQWB50Yf2jDqwPpH9DxaHnffCbryYf1g544gxIdH2L/L
8EsMmCoEEi1/dtOVf99NZUeIw31teeEX2bqwuUxwMuA8cFFjiODaU5GdPn35jVSxxrQ68KapsX9J
TRkglv3Bpa3a6/nAC8vK8SknFx3b4Dw5bLbf55Dq3E3G/cqMVupsxjoW33pqnK8QnKTX6Cbs+QeF
QENWqE7Q5sfkagNZDeWJBU1/zxntmFvV4tyUoCfjkF96HNmng74eWThFHN0YhRxeV5R2Y37cP4Wl
8ki2z1CnPoQyqhCjmFKpH4eP+BUFTpRAxUfwweJxnfppbMvG5eCB+jT0Xelmw1L/jjOzSmO1o8wI
xU6rWOHm2Py7sNugZzUeQZ7BDG7y/4Q5miSrecvarICo5EfXTo07RXZ3m1vhavMcGsJu7ImE5wzc
wIQs0KZPrwCQ21UbMpYNgdVI69/t6E8vAVHUHb0LNFyEbpJ01oGcGo6fLw62t+5b7XX1ejrxLMo2
kIaZziJZXL5PcMRMYd9as+V1rDPyS2saGj1pXnjBRQE2z5VDGMy6/Q5zlF3RJ4UIJzSmlAeqYBJX
ypIATXMcxKF43aCzBdbxMage+fMkcBTAMFvK0ceTMP0x0HOfwb+S/pr5ENTP7X2hAZDPQ5QsJsr4
OQNuc3LuMaGEnP1n6xJfRMsLH1s+GYNvuhKDMt6Q86coPa2Csoc0LRwVmo2YhwYhOwWH0AtIqsF/
M+APkxJu9QcmR5rNER4G4YENaR9Zl4Led0RUQ6CasQQE4HE/Y2oVgiC5BkUbaylCCQb6j2S2k2nL
BYPXfTUmYwyGl4aOu2k1ngfXaqkusI7TbIQyf6MxRjxF+HWZ90+BcAf3GWhpFtn8mF3vw/VfkJ50
AqMo+bgTLqBe6LveQsuoRGOkm5NY3KUv66zmFOIiXxWKSaww9qOUTy9f99C36/OHkMEK+D+EeiM9
f0AXBQh85uBFwdeSvBxioBnnOjSTav77X0MWrLa0joK3BHdAFdx4BWpUUajO7B4R/QXm3plCZOHt
pYFkq/sIxNsyPwh4PMSW/adLFk3zOj0KyAkD19NsT2hVafn+laKwimzot8PvqCEUXKd7p2VXgkh5
LSMkKU66IBF1AXRvW7K9CSIEzPmSoU2QJttJTY+mqatFgFzMEv2BpbsMUwJK59vXkngtcrbEtRCJ
z8dDKrzPU3Cv8L4VwMqVlOUufDWbwLac1Gd57TpMAS5yJe2yWJMh4bkUX0T6gft7kHLm6UrkwMIM
VTWfUGjXDUzxv+lXOnHEV2tdpYABc9+yl339/bD4e2unmG5fBiVOGxTNH8INkfBisVTgux1ZDhZc
aCbhQO2/p3wGAyzx98+4+WvbS1+VLVUvJ8TOxKfmY+Tuo1Ozcest1Y2Wpj72XX3+gNdT6AlwWooh
bVkRQeij3i7StGf5nT2KseRRePdFD955FLS5c8kbiM6KGA648GZ+vR/LXGfFKeqZxmpG9gHEUw4F
MhAO/BrkXhBDekFZryLXKZ4fQuPfYv2713wpv/H8oegC3nWJ4DbdiYDaTrWf3Dme4tYVla11Z1Lj
cxvuAZFo+TFYWvS8DnHrQJEa2M6D6I6tRd2helA0PZT5JtaoFnAApl+99Cnydf5Uw9Oe3WmQT0o9
y6hAXTiymR/hZYrkQhnDrGEc20tntv48MZ6ITHNd9ac//TaDxgBn+adgKJ20ilwCbq8VPRiFmLCZ
mTk0nXRKBB40w4UDSctQ/xbZ7rtMpw2OTGrNEWFdgMCEfJBYkEppvzrtrlCZl4RdO+nt66ibv1UX
VLBVIwc+2yFod0EGCLICSc9FdPnpI8YgqzBMwjSEh5TinEGYTB3VaNcs+MrN0ZRCG6cbaya2TXJ7
KZEtQX/PTxbFSpd4ngF5UpUVtpeb44Bjo2jy8zWVEYsVpLY0HOvpIDCAQpO8saEovQWCfXLWw6VG
vaw+UJq4MUPp2a8vHfc4h0mlQ44BnC7+STcPIp9/DQuJRzM7C6ShJgawndLtET5szFsEnK1P7N0R
OVHugQZKhDeHNeLejPvQ07lPuci0oT3DRlpG7ggS2zK25yEbE0ZXsKNJSOeKnm4379baiftWSfMR
2+LifN4E4pbBShQlgLlctWG/ptMvg1Nme4l/4IYha/4w7rPsr2sQzpQnBoxS5nsezJZ/6g5i55yR
y/rmI8/yIFg64uVpA3AH1lfjgo3KzKbZXa8mbOP/YRb4TA+TZXGN8wRgzxRgdPYN/frAhQDH2bMh
Rz/0vmCnMtO73A2/SrKrFsLcFVlX1K8zrMgMF5PT3gYYWxm4QV4OmErJjg+a8fFOq4AOGa8iTl+u
4V15yyb7HHJete5A9aqcSKZNWSoRlvOWcfbm8uCcZ2SpKYBPjT0Vry43nxiNkaHuZZcEqGbhoEVh
gxpw1jt9druIaiiyLMOyIyuSlie2dEsh/ft5pRIErqt+K7zyf1oWtNPnp2d62jQUAjuFLPz+5anC
J3Z/YclrTYo0iGbT/jeSOalOhZ8MjwRZa91Psc0m96Xrpn1t+ZuOJj9XAnino91PaPzqs+uED2MQ
qPIXfFZQNhaYGRle1mqZ0NS6ok1T3r+DioIbid1/2Jqrwd+uru3gh9/QXSh8bbqBJj8iVMtw5Tqf
QzgtHXOpm2OsEnGMjtfxgYOE/LhAtXMDm1lzr8ZPN7Q2XDu522/oPteIdhzVW5sqm1A6y6/U1yBq
1CtYfWacdRqFOBfkCspASIwtBxCQKrQYh0N+TBL2Ln56Lq7fToxF0Mc/kKAIRr32ad6d5CIz6R+X
m9U7acs7NK8xqqaf7Bn0QIU6JXlzPWCUzHtj2tG3fp2YQXTOfqFcBgnguEBTfWuTZD2DzSSEjGZX
coHhI5PmjArD8IRMm9cU/vC/ie/VqXAeGJnuSrRVLu8VnXE2AC3myKub2GETRpsEpTUbv07Wuau6
5emcRk9RBKpVazTt80b9+/Wyu8J+Lib2+WudnLcIXtY/Rd6PFJffhcid82A5Er6GJjbOIcC0BSGQ
39Ka6diQTvgsXm5VdVGRLv98yrm0it2F//jeSIKbjV/3gq0odNo60RCAi2MeaVYkpEUQq95FgGhR
zE/FuylNeIJ/chB8xEAaQXdf2gKGnVX/SA9LKEAv0V18oYS/v4RQYSDjuqHjbFt24R29+jWNASzf
XdPP2D43X4Yxy3Okj9PboEQMJmpr3ad2gfUHpgbzf2cmk9nUUZHLFHPLdNmvCwtCDNgLwPSZ5Rsd
38FmaQc9+h4iidGxkAjUXo9RVmjSdunYuPls4Yi8VTjO0xRVaHSADPZqLWKLCfFpZ9cO4LE2dFqn
0R1G3+4F/j+vcM+x5VlSQ+KA9lNrXElonFExE8eRolZmCUpVKQDX1kguufDYEGG9Blol1eDuKm5V
zMbylfb4g7GAjWzgAa9BHhPEZpRaYPRSVhR5WUIcv6JHp62YgZNpuwhq/d0AVHA8RMtcVZfa8qP2
Dv0gaRAjbBS26YjDwKVgCmibnooghtFTqbXdpfHtzytPssaF/9w0lOSBgMEbXDc2irQ9IwmfUokl
4spGoJHhBAHHInBAWmLEVvoTVpaK5wgnDMlmCpo+ZCU4w3Svtz6ae2wnG0WO8Q/6N97G4sfp9/f7
qhMnpqOmp6/rE3RWU9AwBb0rKLHkAJUM9MdZlne8JrGrlqbjeFtX92QppM61a+5S2ZGiX88xyQ+D
zn1VbKbf1N3uZH/m0ZDcSBgS11ALexiaAoznlWIpjVOefrGC+cpi9/GES9U80BG8Sh0sjMjxrwfg
tqg3tM3x8GB/xfqVNYE+jwmjLw0kr044hqktJuplOGRjHD2YFnSms4qjeAbyaSszRBZjUdksJkyN
TbwWomjQvaDM/58ABEQhT5Pnf1Eq/4ffY/8hYt0et7S3GsgpADplcEmMp7emzn+1RMlq1u2LpGkh
xR7r3E2mrPNew+Z9zByYu5zJFuvZe7pvOzchpJK0rtyiUWBiei7S1JGCWo1O8cC2WjzIRJaiokGU
bM3rlCWoGkTnEhDF3KWcMiZgpJrgym2L0c86QDGI2wYeQDG1C84V2rlrbAW+WUoKlTKIacjdhpp2
S352u3sG4YsE1BNvatoGgTZsX/Frvgi+6mr+jtcSoySSZqD9grzCeF+NvP5w8MOQ6RxADF30O8Vu
9V1FdwunhDFxcP04s0tQfFoRElxhGVm6b0G5Gj9njeCo1wgHPPOvPvFfAoBkHgddk7l6uTkNTUqt
qRcC6MXb74LAdWtq16csNnjf8XinZMjI/c0NnNjQuIZ57JEs7kD1+3bCM19Oe3pYCScOYdG21fr4
mN/aXPWgN6POH6spaiivK4zkja64rNmXcuw71gTf4Bg6i0MXs3yvKJ6yKMqg7dP/+gqYoOiwnxs7
6a8C9UypZPhRsB3KLJOlIDcHZqx2IZRcjoD9fUUNKJelnU6Pc5KWfTflKspQR+D87NjZbhAHXYF8
IrhkMxiHXRVGB2/P5XEeH1grElfRYzwQKZQ7JUVoYBeI86DnvbCX+GszZZgv4CSkaE3i0yjUei9s
L41uSsp1EghLWz56qMiTTacSnPNbdzZx4xqCX2AV+sRIILTFIYgmvDWQb5UnzdAuE7A0ZY8HHEus
Z37LGseV9nQ1dzAviTqqeFlWrpAFaBrpgFovUrkU7BkuGo9j04LJQrVQGm5pAsaA1gxMArXYOH0E
kTTFgBDd+MKHi48wtf/mC1hikZVpnGZIMf/dVAmH6SAiHhuxj8hD3Dgi3nUvY1OKTDSVL4h0hDen
8tuTmmPPMJ1clL186I2VdRro6C/AujlSNRyBzGRho6SBXunctXKNOsyIq/5VZJu0F6A9pf3f5kCC
BrhqwG6GupmWncz/nn2vq++4abxYXhseq76ol0B8pZ2ss6Hrvn03I2adxolkgdvnqCN5K1gLN+iX
FCI4jLFQJ5bB/bQ2qh1EJaKJNt3TiUdgDLAnCk7rKpWrnACgWfOWtdIFCT6rNazeJlhnA+7B6fn1
wdFlr2EgE8AuUKF/UnJSwt9+2k2utoyK1lzRU2MyKuce1JZH2jRCKXlJBXVb+jo/Tefj5owtMYYP
qu/TfA5GE9SREP7NZptlJfHMxMYC9tHJxLFhuTfvUD8qnVO+bcufL9UI820YispMl2l6CEeUIC+E
6Cf/OnFjkWgbsphD1eW9/FkyVGsMZO4TI8v4sKpEM2L2gbzaDcKowBbY7EH1B8BRRRRutwpM0SoK
cY1te6pbh+9SjqZ4qC61fitiigqPch4M17Q6Kn/uFvx7RDgahT0J/GvITUz60v0789Mo+lZvO93r
0J44RibJ+xwC3ayQsxw67AAJvLJ5sDs5hqgoshqC5P4RgS3Mv58WHkVuB/hcXGhr0UkmZb/WDkO8
ucE4AHQt5PwUYG3CQuSIZYvO2COSDRqlsziaH3a6UcrxEAgI7W9fMI3xMd+qbuTEY/3FP28EXZiT
5bIVr+uq1xTU8Kk6VpPGqto9+0wAW6Fu6BZzXf8z7rMjzV8/6qmGi/kOFFeb8JgYps2aLejLrsRl
/1/1r9Xx2bdnfRYFx4ie1WNFunsTTBc/EtX4WqZIjyoT/Bz4LyWX8VoQGIOXiiMIpj+TJTXz1kC+
iNhQUps3/lMDP0asiFDdgsuMGdiNUlIaNLhBuznC8POZeW5Amg70X9T/pEJACKsOQPvTr/vFnadL
HU2buwlyjx2uqtllc7cxRdVvzoLwRRXboerXN+ce95Q9pkk1nz/jVtorZNfOUdOxJLJYvHMjyWeL
/vkLMNb3Y8WCbhfwoqW5K2kw1/fwW/wyX9bPFq+OhDnVFuvCDZWeOVX+o6y/zVAAQe1BKzbEllmM
wa0y0/La/zBsk77wMhxXng4ggSxMqTe43pF2zPXxB91TtpOlIlUDAJI9JzyBs28yb7C5HFksjCH+
H4JXCqnePru6yryNgjJ1ElQY4NaM/E+2bWOqeUFNFC8NdxQ0SDd2VgUHW75LcAhn/aWfC6NSSUT0
ye4g1R+RtUsZbweYpnRxYZ6bbAQB8QBL+9gd6E8yanBTeppW2UAWRJCCaX068ENTe7NQ1MlhsWJw
AkKXflSW2Z5eO9buuExFBGDAryLTKBoRio9vrvAGs7AJuZcXM4D8EReY3QqWF2pFOidHHhUUmyCw
ZTHRkGnE8JAHQLyta6HtmJRThGCA7FDY9U2V1qulRq9m3fVfRDTGy8CU0B7+jp9qmyNJOY8lK1wV
j30U8b0KpTeGXLpW91Biuv+AJjBNbqWLBDwt8OY9tXUI60Ojio7UA+4TXZM4Z2qGsZel28+Ig+Fx
yy9q+I1ufwgV2fpSen6GeT4bx2FO/ztNExJpCVMQXT94tW34LOhFNpi3vZJBLDnxbr5wslkWaKyU
CMWflXthBemBqZCEj5oQ+f5/SaEw5QU/fLLIqcbVvfBZcU0J8kMjWrkkBbtBFEc0fgT4QvPMDO7K
R/hb5Tue30Y+bKeRaff61NM7Hfixo3QlL6nauyV9rqqRwvant4XN+JpjTIdJ+C6O6Ni5hQlAdOc8
Tmd2TwCQ01qeRFjxxgBOuuMV8G14tLMWWccGZ5/bnkIzlpXfvH7JLfRxAUM4GyfhJChhBtRWG+LE
rkS6qW+AneNC417AUvoI9WADAdXBCmD6ncybYf/Hsoe1myhOamOazHqYB3/CP2D5AOEz2RBqLXBO
h4JqseEd4b1jpslTZlfnaNob038CMBD3qmVggFnuW57Qyfw/ciMLOeo/0AfCHUYG1GGmpYuZXMtd
gYuYd13bHE/uI4nqC7IzZTKPXHgUNyqk8VBfNFbnNgbp1kGAxRYHK/pyYIQBkay+x9lVt0Dzsq7z
M3sbaTNIhJzfD2tdLKDa7TpEXlJfPnT3LONy2n/dYTr5n84i/96/hYXAFeYX+F2cyM3Or1uHVDqN
/ktIETvreobY+FegsWFN5yl8xtqKCsYNUCT44/4JvTA5jeSwDAIouukMXN4bSJuQI/fUQ9UfrRRw
qSruSszbalJsldoO+YYuOoCih/AYaoLc9Ib0jTmCkLjgaEB4kmjC7OyKbCV3AmvlSATZPoOrIBwn
zWxQMUb7yfC3zOxq7wNFl8p8Ev5c9ZK4iszzll7AZqtgg0pMFaZKx4DBD+1OpRfNk022WjVuHUy8
O7PXAIYKzwrdtJHgSqCN9RLW5kPNFgORiuBDrK7YfyqrrAXr/Qjm3GyuOA3YqIiP7a28ZSUnR0BI
NPeJQ9fDm/L0GwOkqG1rYMCncPEPrpfFVyUg46vz4IQwmyVKv1XljBJm5pbYfyCvUeUQpOsoiVfV
IhXMjHunuxhwH3er9BFBSSYyZ89Bk5ktrzbwpYd6nNJ011uGJtVFHnHcVA+eia+y8wQ72xaJAigv
/V7Vn5u38YPI3bz+ddXGBaAB+VRfWoow+oWP82qW4pljlBO/OE8DHDL6AZhgCkoNB2BKMT0k+OFx
PDuMLacVUUqefFwpyLoAaRxPqLxI7F0HvSjznrcCE1f6uO8fEoFVBb4Ow/xtEVDm+jT6lBjiJ4KE
XW3wG/V7hpGtVoqbex5Q59MEShdsh5ngNAR2zmz1pNjTiqSjp/QQmbeGKdNVRrXgfVm6GrAe2B7o
N+3dmtfz+p1xnD9qEByeyTCLWPYzRazKVmgJRg1DzkeK8jeKj861z7FXP0yqbYGWTPa4qLoRiIcN
63kLmC+AOzswxSRJ0yC1ELMRXcGVF2BvBzRXwa70lktvEe54gXhpv7pzxIUa87kkTOv7jaN2HLis
lAyaPlNOXJrwUEa69KXafF3DDs4VSRpPVDBknmD5b2bfDgHo5fUJ7FumdssRSkFHTZ73Lhtvf/bd
+YF72GtGbxypssXMWsP+W2YR1p8cUHMzlXkZc5wVg8sE371YlKQWsn0kkN68j54GunWXiguoRwKc
Qs27T3WqK83dEja5zi3JIfi55GpI3hKxOcxd16qgljKb5FKEtumD8/5wT58NCzONALiPpRug89dv
LS+X17dhgdqn1Xw75R0015MeKLwkkOnlDrsENbRXuvN1xkaAhAb8TSjWWiC7aqcSLh3Ol51j+Pom
gPX0OCbz91eKa+P7L58vCT6j8cD9uDyoJuISyusrNkW8DPBw2+UzXrMgUfA3uW76zNSffMXqxrFU
jTN5uVZTdDe9sd52EAhGSUsLM0zB1fWQmdwZkLPiNJdpoQay6SM9bxHP1NVdPQoslf1fZRsJNgE1
FJpsKw9UTKe+XVH3u1qaEmIRlIc4GhwNHlVnPOnBqvHkN2sMNBC65VrmWS7SH6GF0orH0hAoQhVv
Dcszje8fFvRz1uYxqdPH2t3JyLQzeo9/mYECxpnJWZf7xqxXXkcfwD4gC5yBQ22j8/bDXp5saKcW
/LXXvhAgyqKMSIOYKgIewg/TWXUcer01Frgy9o6AiIwT2QIt44yVhdHU0tpp3i7L311vs2139AAY
6fnB1V6kHLRWqAs7yG7u3zyqsl0+qEAg7QjhO6M5ONoSVQtqyljzodEIauL6yZgWlo/1SBKB13Eh
wN3Xlhh0TZuldnjKU1XJk7+PZuPJc5dR4D/RMAgPgHPpzxAWPd1l1dPrzCxoEjpEDPHtJBEiXt7p
GfQxGG8cJRFZYZedJL4Mw0HUaQ+SAknQEICWSHs6gQ8jx22srw/LOmUonCeXXElJFBoSj3CFAish
+9i94cN3pKOM8ECCRjoDp3xYbppNpVC3zIBDls+ukwsj86P3P7v/BO/QoC8ddv+SatNwO1ob4lmF
RqxJEFMat+uhrZQbjbIqdq0s2yWFMBIvRkIUhJTM9vgWx9g1nrha46Vj09qUVKY5e8OVukW9pltn
TSFtrVemFrwQ7OqItUZqxa6HBtKpdj0LoeSn2JPcxngOUCMf3f1tQQ1AkVdO1f8olZpyrTtP9T9K
Jh7Cb0jzT39guOjQ/scQWIAZQFG1tgxFX5JdpQ69frOUYpS/IfFwjeystb9OUc5j0R3Yr2WBLqWE
095e6y2e3Zll05qG5bJ58OnKZW+Sjdn44LiDDo8LNfYKcoAe3PYRXCDzZrUvvXAF0qHU1be++e2t
OrruxTSvspv5H8xIMWsFxnQooEaXx18gccJKALI/6wJLz0ML+93hX1hBPJN4u2IfTSLidFj4xRhq
1a1axEV2iZ2ghH600A8+Hu51hFX8U4hgWm6ezp4VQz/z0q5Ndbby60gY3ayaCKVClBISf7u6zaQ0
MG7gqa/+KvEDTr8m0rEI2Eu/OUA8t2ec5jwN4UghB2iL0cTVnvu6Xn9v+s+Ib7EoLHOoMoZ+droZ
hgLAyj3VzqJyr4ecw2xnFGqke+Ym0fUawcjnsb9d887Ud5vcZP8e/1lACrs0LtYVKoQ6SFIWxp0L
daXFx2INrtChm8ikHMFNcTAniiATSfuZGBmsbbCDVPkvi3lRvSJJXJzzsnuf3W0UlbT5tnggrk82
hmpsVo4nZH18dphMwZoEEto7JdmA5TsfQhwFmXJUCnjx50kgAzyC4ibE98UB4voQLntdYSj4/bBm
uRvSkvqJ5hZrGE+qUYdC6XxrhlDWIgyo/9mbUdoxDFjaHCUklWBzgRUOPKuSln01+OHrsa3WcLBQ
Pr3cbXN9y6I7RYHv7ak/T7nadRgIxdih/zojY1IIl2DAX9W1y0anyztQ1LU8cWTnfaGUXz56Zcnm
a8SQTe45SIQfvQqXr3S3JmBb/y4q9l12unmRbuB/YCJj0H8pscZB1fy6PoEnrTg5BqGLdqglCdTm
bg08z5HJ5RwBfasfgU/vewTzgLeoBdJfEzrX45D6/tmJ+Zdy9USJVyd9BaAmt6AR/oEhtp6RVE4Y
LbFPXTLyjvMOc9XHatYdYZRzPIouNeKN9dYKPPZleYiHnl0elAhG2pKVHNJJclVLMwM3gWc1UX3N
d7fObxUtFAiOJlB8Y47zib2Yv0jnjezM70XIHh9A3CaqVdcSwUu+KcAn7DXyJEUVMLDdMiC/wHqK
zclHspbi5dB756o36PqLfAtHM1cK1hnL+98feyDHiiypPo5CTFZ8zzl+ojM+Dg+EKqZidhCZx1xP
wQSoKuczRq4R2yFikQXzVAkedUi4rtI1VLKyKU8yut8zkV19OgKnLtg2zXRLibCOwA37fpU4xkeR
9vDXTELH5kidxLqgVpLyxe3Up/UBSNle+ctu4XsJOOn2KmnAo03Fg0LbYH3n+fL+PfsHC7+nq1BM
19PrS+pkk0XNvQm3EiSWmXNJzOlfiI7zJ2CPh6P67y2Hx2apHwu/KFSO91LeFjx4JJWMcfGSW33x
ozzkoN9QMwcZoC4a3N1Tmeb7Yi5UxYS9/ZIzo2e6sG2QcXRvia/u5vczt7ejPClJB7v5vdpodElA
odFqRvezEEhs0fdvgfrd5FHOCDW0BPUs1yY71nvEdfjknVcVmMsyFY4B7gO7gPnekmVUcejFmn79
cGflAfU9/hXhArzD8K/uLqhoG1c5ilJ+rAgHX2yTNUqrNGOPNN1Z83RKhfHQEzILkE7pIXkVCftO
olmeBce+2AQcx77SiSPfpVhkR2rG1cAq1wm6vpyCadei/yGmTVzQ5msy5xQ1iMV0O2mJheTjBnCN
YYDLQgmAX28osl7BJwuMyJWWOPiBmzf8MdttM11RMibtbJBpO8TTFluNQCTp5eEb1OS7D0AZOd+Y
OSwtgGt0KTY3s3T688Ac0FtoWiRmnqc4DRjGM67q3FAylpaqB4hwSylo8q0VaL04tgtX8QVB5y+2
gqaFbsRIsAOR3+IpQEZ7yjEQ0fWuMe7dW4K3q1UEsvPOISw3Y+Cjao823n14j2vPK7/+oYfuQI6Y
1wxAKcFsX43IWAhd5Ivqisgwxm1th8AUUIpBnpVGrOratOWi7PHyqDa5ttfRVTg7Yg6PdOT4WBlu
t5dBqp5W7sk2aDaO4KReA9IeeE7w5ehenrrNpOfKbdMSWQWmuG5ZWd2RPO97PFtIAwWcHvBvsksQ
RutFvCvhe0rNHsf9JJ4MNSK6byIfOtk2djL3Ayi8f/KrJI2WE+5PP8pSOsmL82dOIGzHQTAxY+Tv
MYHS/G+hvY8Y+vMmx1NKXV6MDgKQXgTQNO3tdT95cT3QxXNC0pJJQ/7nHyvcGbrrUoxjgUfr5ScL
LsR4Bqp2j5mxNz+NSX0JZedUW+Js/fVQYgYlUvnbDWsSWY3kFT22Z4TKNZg5Y/kriig613IQTSS6
xI5TfTKoghAy8f1dqAG+Pu83vYxXas3E6u7i9bOq7qgzFJncL3CLT1irjN2aPCfl8NvN7Qg6s1ej
+ekfXPeP8LlODdcFnqDF/r3wL+3U6QfPxcXpOefxZlWPLTx4NzN4O+XTd0vzZSMGUzjIuT6P+Cbq
ClhB3Yv+WKyu8ZzHChZcK5lL5hrqD/J8WFLYpd4+uErFVc40X5TxV61wBfw/5seIwtA8ciR04Tbk
qXnkKvaARMrHPm0v64i5nfEOOui0Ey3WGFUK65QUrwWLQvZdUNOX1jYmAL2JtFSEaoLV8QCcrrAa
GVB0kwiACn5b/ZfEJxMov3bC+aXuyV9CJCbPs9DPPb7WAODIKte99P06jh6fW920vP+8fBeLZv23
5wK0nAIq5U7x+Unu+4ydgsrZ4BV9Yz9sk32SSXDdS9zucqeNrg4++PH+z9yQjSwQNW+FTn+EUWJz
G353n4ApIfQ52+mKnSoLisgZQFNrwve7S2AtVMSpDZME0nsO3QZ3fP3BY8Srt5pyRa9K8GhLLSkU
eMJFafdBGdEvTUcuK51Tn6NlP6p1kKFPTS14xSzjU7uhFWVM2cWrx2dUaxULMqwwst+v3jDDf2yE
SQeGTR3Aowm08HvGrFtiReJHyoRXTYIO1BLw7ncVonIavTWYc2wWrsIaa0VemRqLUv+6Ce0wWb9v
dd8BvFNKiztMJY1yorIUeR+4g44f3zNr3oy2PIbXSnIF97/D/1xHGBYOCtO1uViiLqXLMQF//y6n
LE1MFsOwtGigZLl0F821gH4z26qNe+N47psWnyttwPtfm5mKxWlvzge7XUlyvwjPmxpqYSfdfZo1
wrfafRPwtDH36I61VVD3zzzzuG146moQ7vy5wJ6N4/+6SS67g9DimwRQ/Q/EUAONwTqoNtKxg1Nf
x4e2pFsrzCMsJvES8CYfoJl103BXx8Ql13dJxyJJFddcCQyYNBJIrf5s1Kv/WwAZFzud/mKKkyyR
JjMSbafSLimHMZtgiOVCbX0+L3U2Vyb3PdJgEwiKTOZDc5UpMQYeho+/CZ76GWaTZQ68+zgFDywl
lREJFjSQR0j4u//o0OXRegGDEIPh7VetEmGRkF/L2re3Ebmh+qfRXnLRqy1uqM8LSJ5/cFc0TE5T
qPmxlA64XuJJcrZar4/u2j2RaAI3LHpYZUofOX04NWD/XLb6UZJvxewNV3Gc4jZohddFqPPLxoQl
sjdFpoACk0Nd6rdPqwqEgno24W42mGTS9SmPY3sAhpiMElzni+HXs3XOM5Fu0KtDuqvCcZVmFLcr
+Yq1eRzXG/7bxDOgepWOLWrt4n7y0md/bpSYGuhA7n3ZvKjKNCK/RbJuaUYZfDeDe6zff3eeTA/8
YP2as92SECspolO8Qk9I4Ribzogb58qeiO4LvB6gXZMPNxcC9RChWTEzqA6QY2Fq/npPSLzL/Opn
U+ZFVhhvuQGNLd183lzEs56IhvT7x8x1Y5qbxw6E8ow4IDiUh7/Lr4bBrX0szSSpHvaoqZyENOSo
rupmHwYA86buTHiL39Ta4+5s0sfkpNp8A0wZdPVAoYfHdcciH+bkXq0eiZzwSHifKBP07JgZTLV4
4NZpuaASD8JCGFIxCIVaAYN13aldTCJMjJIQIpnEgenYwhcZZSBxFasPhyvGxGgDA+G0NpWGGn0v
W3DJaBuPQRr7byTZsWukf0rVCDK4EQGYqRhIo6lEhz4taW5qzr0OYsBRuOFrRkEH/6lu3mjjqZ2L
/q6+kcBqi0qFWi+f5PFwvnmlIAmWdXWDCTjsvGkvoa6+Vn6G8KqRBqgE7CVvc+n9nUFSkkMOB7s6
b7C+pBhi4XFgZy89H8WqMUrJQJjs+YpdDG4zA677GTE98B0KARWMCDEo4uKlSpIHpFPcQWAmF+Wi
jkMcCphdOQ4+i1NIY6dc9NGyv4a+qpWyD6BR75eb7dmHddmFc4N8dEMOScytC7R9w5p/m6JdoYkp
tUJmQRIjLJa29iDo+jk0VjNvbOSXL8Fe+WUVYyzx86Y8D/hCOyJzM7tX8ehTXQPTAnTXhySfUgNA
Vq12iTOk/+NVgS0g21JmwbAUerQiBATEfLqfkNh7FPVF8h9uy1wNeIketQ1KXI3m+lMxfZI63aV+
RbfrpfuCBkIv2VxAplMlo34YJEKqIYbHXEZP2oYfb/tLhWNsG/pNPawJoIUJj9DSi4etkswqS96s
IFRZRtU8urh+wVAWWqUd2h4l92V4DY3rx2XCynq+W9n9GORAXllbN3pgdq6HIx9feby2Kjh9xpC8
ygF0K4nDwbrMllTC03jKtHT31KbIkZM9w78sMqqNfP3hj+wPGKYSoFRvEqiudKW6Rmzxay2tb1Pl
jMOa+pnPEkgFIFUY31ZFzCyowTUAIR4OtaQe+ZMeeYPaGmYzd/TwFWR7dEZEafdz+RxKmx1s12Gq
IJauOF5Jf2cmJqFfQXvw+mf9dT5Gq+SvNvGa9CNuufiO/hHeAFkN/dt7AVyDXkKRAWGO6ZErxOrs
obLhSwVd8BmpZXZxC9I6xU8WSVR6QvpNvW19ODxo1zg8LBVKrt8N6DwfsrNXk8h5GAYZwYiT779p
bGr0U9Wwfflcrhy3hu9nj8TXzwadjUmjx0s6penkrgquJqTlclNlUkPeWVLxgceKs3n8L9msnehN
XeEacK+8rkRQ/ieTJ+G6/UWGGwGR2RF5AkdsIm3Ui8/S7Ej2Gl+UY7jofS63Q5NU23o16DDTFu3u
beGjlNBs50MfGApb/lARoIoDQnmXrQusPYS5qpB0j+h76C/bV4qhvYtUwxpcVNVsXfqDhI4F5Qzt
RJV2pVyT6Uvu0xoTQBSZYCcmNb+q7ah65SiJD4qfI9L0N9BgX2+sknXwF9YsMas4L4e+3UCXPHbf
zSg96j5Eppbk8nTq/A/Ra+GKw1v8muX18RVyeekV42LCfgm+DuCF06X39LukQmObkunT3pIXr4CV
ppdzOX+3zQqbvgmhpfRlqcP5gXu77vEPzkUwZomKOI0TCxEFFvcEjq9W6rjvfBi4ATbfT7krw8MD
kWYX34/zNUnooMSUt6WBv1ZJ+TMEejeShQxsLIWdK8fPLxAB7dGBkn880PZKL/SXrrhpPMw/wfmK
sl9vb9md79FVfL7RSvdNVwvC3KLwlKw/NzuOPFcD1nR9wnz47qspoqD+vBcs6E8oXPw+vbR+1BsF
JBYK7kJJhNTnFSnxnf8ClRUJ5RXiFkaieftBHZsH/4/mFvdGAEt1N2I2kf4PAzsvJrxvelM8Y29z
XWJrH5qnvaqTKIn3g2jCpZ7ww2T/1G5/CE+ZuTMarsqstqVpxG5lOQPjA+M2fZoLZxa3qEhlWoWQ
PNYc6BPN7BCPJ1FevV1EiBg91OA7au6Lp15B6sRTrHeSz5LX+tczNXEWoEAQSCRHCxQhv7yINSid
uvaAiP5YSBATMtghotFvX448ivYi+7OXYrUKGsBS6x8v1fcVAsYqGHPWrOZc0ouNVk/h9pDECetv
rnFIDfp1Xh+kAhs0hI2YnxozGddZlcng6PHJjNilRrfTQXRExtUM7fiFYxsg5vYWN5BXaMABJj3F
WaZseE8tepvs8mXmNqIFOG9fzYKpNZ2Yv8yw6XOq1UYzVS7NxYMAQH+vzAnkYEqMU37UMJibrds9
JKHZRFcq9XQ2p3Bo+r7m8rD0TCNyBhLHjETjpmgNgXGNnzI9n58AH3n8no2ekfWLy8OrUJKwXfDe
PdW3QxOBNG/GpXm3UJT38l2DJpDrCd/8n38nIf3WmNjYvFfRFMT2eGU32XtZPmqE5LKEKRXxXNL+
vpTOelZo+hlkWpAcNZDNsz6dxEtbutkt9mfC0Qqbwn+Bkz1hnumf3x8NWtkM2RavI0A+xAaqr6mf
FDxVpx2HwJ8egBpsYdjvHJNhZWcXAiw0GqParl4HAKzMA66JHJpSYkURcyaVX543AhMEsHXL1xpt
ctUx4It38x4ovztlUSe60LAGlM15UURCmA0cgdAUhV/wAMTOyM9IWe0h27FTkob/HX1FhpweR3I+
VH60jXSWtGLlxoy33XG/wINe2MOHXdjyNIdadEysGsrEYI01L/Y/yVbUGGLs+DgNVtsYuRnTQ9JG
RlkgJtUS83aAyamTRM65g2T9luw7s/jvvlJJGN/aw9VWBarh3mVWQnGeZrrychgQP+HjoaY5M1wl
JirkHoF+hTStjQn++KDlI0Ftj5fEfzVzeFaRYprXnJfgWoh7KVNTIPDHVdw9fx9MX1nP2tUln7JW
eW+CrfGchOHqt10S4oPpqfBv2127+QK800u/qiZyqwqfK3Q9w3JzIuiISNc484/Xg2SecteWZpxT
3n+UIs265Jx1K4KSd9N9YosNAM8PlfuWK5V27VlQvOUH7bgueIDPXKHy8oTcN7LoPcborKFgPCng
HW5n4ON+0ni1ZfB74Rd/DJNhtc5R7GGRTF5YZnbGLGWWPu1uBzWJLoBSWM91DAfhF4vcrfiEKRA8
QyTCkFXqn1HGNI8A0ivktHsHofwaNRSJorwvHkhzrQw5+wERGhm9X8lhgKj+NCdeuOr+xdc562zX
BK/+ylerj+se9Uer8eAXnDmZ/kIOTrVwV/1onlAxLsrgOAdwPrrQX/9rAd5q5JNhc30hrWkyl1wu
YXV2b3m9pbVCM8i5dd8Bj2krp5dES5k4yubmWbBOg4NHFGPoBJ+W93HohoRiTJ8SXDOJql3Pb2yB
UG88r4Q+USLXeyVrJiBd53DAI0dFUCRKV1XnMJxqmdswgNFyK3MLkmXaLGT2G6LiAbezZ+ppwnhy
Hfl2C9JaQtxKGGbrWBFznEL+iO8EZmQXe6KEhu/1s76GYWAQIBR8ZNUUiFHmWtKrjBoLXyFvP09G
noR6mGThAsXsYOgDm0v4aBgP2EqC4Q044j74AWbbIl03cTKr0uJShFNHRW5iQnKAw2EYKZ+JMP3F
DXvPjj33XeNsYJ4NHWgP2K2vpHrMqtmDCS/InuTw7dwu/NCkUlOsNGdOfpmZ64Xb6A9Kvu6WyAMC
bs3/9Yxo11tVY0VpXAFPsoebaYtvKvxsaidv0+lRMuxaosYUIbKBETNR7uK/5BCNUnBiGrdFzpmi
anQqVhFea1udWmu1AHlXSiC5ykQbe5hkhD5t92M3IZr7YFJYYfv1vIKkkSdFvL38h/qTqMj3uF7f
U2BrO3OZcx7ZlP5c4j4PCWTMur7XcidB2GXQv92R3l24aRTOhSbfPbpsssyO6wEyI+e4t4v7mde2
5KyXMmnlSpYGXTQk6nF6e2PLh8I3oxC7vT+u8fZrSBOhrLkiz0EUebSzsNrBMlDe92PntR9qwhVF
R7RsF7255owUChw3hrwkxq+c2mLcpfv71MW2mYT9CskMutCAjaKjowTt/qSc95U3gNoFqdNI+OJJ
NC2P7zHnmYrsskxqcArYWFh62bvqE3lKzBbk0GiMK2anCZh4Eaejh7ki4GZwBhIEeCz0NDUgrLig
ghLLnUyQtn1emI81XqMKGiFhbTiCILkuS5Wl73bcPoDYuwsTCLAYB6W28GRK4x1BvyZPWlzkrUQq
oUnpN/f46aQzR0cgulfx8r2i6gMnE+oWy8+rMsIc0jb1iPGmVq4+r15lzfXEwN8dOwvnnvBsKymJ
aW2d4XZ/kX+QbcyiEdWE1pbh4AlxYIi/tJwS8fq0t4C5C6pm/yXThN1HU6SPyN7qjStGXBibHkeu
Wchx8akCkJ7r3AXgN9UsxAvDd5AA6GTuVVM0ACf2jz/fm/WRLsGmeKD6ym+4f83bX1y/RPYMi4yD
HsZEjr6WSiCHWEGr3uiqukROF7xj0KXR3dIJ7Tqgausrn84p4NncUpX7z9qMz3mXM09qbVGwhfbg
8zY9fswX9hsmUJmTbxVuj3u09dgoKLtj1SUiQlVUmuBaCWTefYtQdHyGca6jAtTQS6p1XfBAlySo
E5zLG3c23a5xTw9XO+SEqwoJQ5/aNNVAlRMYEpmPqX4viUeggGHpVZP+SbIHxLeScowcRbnO2ESU
tO2Q80QBuFZNqc+PmIGwT29ZpMQnWYSbHuf5h7OM/QNeBg52UWgg348A10kxnRO+lbDhDFJ+vPwh
IbhZzKYP0XlwdIBGjDCs69A6SjlwdyyJxVMoQUw1M7kLOO2F8hCGHoKvfDE84bpBZ2mgjRVftOyP
ta0RiEGtE7GKA9e+1Gs6q1gVNS/GCOcCtRziHnXTkK8wgfCu38VuMCvHBXUhQQ9k9Y+RXFKP4P17
J2x9WBYXPWKiAB9xrJ1HApyxEXkgBfnY1MotSVVz+2/CqA6kgHTvwAhL9rolyVn09mHfQyj5lnSX
hTJU8WJCIjKCQenE1e6/UgZhE2xrVlJhEMqlZwoujOh3PefH7lzRrpUM7bWR9vZqVN4yzkFljsnG
tTkPsGVowU4XqG2bG9zdsdLThlrcIJ4iiqQa91Plldih79mON7K6qKBzOuEkt9CYuXBACbsN6I1O
NSB5O0mokbn84mXUYzIvql+RLQtySYu4SRb7pygSGuQ7JlufAFla8xwJLWPpN8DxgMMyyfMUY+2h
NZbO9/L+6H2FrN/geFBPAesWR05H1kIG58FI1vjcRP1MPMQaUfh32xso+xclxRpYMdzdtmvvwDPt
vG7ttQcft5p2qtQ6NYsY5XJDLEUdso2PRa3Hw9MlL/FI1gWC5xfNScVI/4zIdvqjCG4q++z+Qn3u
hIDyCo1PesTZCwd7Ixjh+YJ88EemdpNf9TdeKX0mb8aCmYgPKS90B+SPmNd3b4GJpjCojagty/mn
SsSrmYCeSZxxS9bWsvswB8nkai5pUOS6UJ3BtAjqauPPc2b7jFLXTIUTycQ91XBGw/P2q15l4NHM
y+a73EpID2+hUjQpm32MXVyemQQtNGuOERCN6/ATznx1qvq+jpMz9wASd1Nhr7hUFJ+KJW4fuN4k
OYoZJq808iAvVNPAtDfu37Pcy5BpkVfAC4Er2/e8XNBOXkfxqPEXQzi5e2GC10WvTxtwvqgC3SqT
RFiIbIhZShmVE5bpeg1RUhDeTbVIf97QpJR07fDAqgnejZ2iXr2jZkyEUcJw4c+o7SEU2/Fh+rIr
vW4U50EKD2Fg/EM8yKBUyXVrwGYDaxzuO2RbV/3kmCWL9vkQyyTtBghPU3aRhP6UpYPk3xxrk9UX
1CtmuxVp8a5Yd9o4a9HaLSHYN+M1GgOicK+FKb46jCUZRqhxq7KZ3/nlM/KM0kf3wmd/rS/EMOFn
g1HpfEHW/1PrgFO7v5vvuHP2jCk27v4EvrYFxchWyf7fgWH+HAZLdnYw4vWVerXfdJFEcJM3MTBc
qPxn9CRPFX6PLk162OY7zl/G6tqqYH80y1T/o2CBVdRvcuza4ApkIJ6PSforoWtMUYyklikduKOM
roCjlmHAPxOlCjqZXhNOkinwwdBy+B0Xc5FbFt22M+BZngB7FErq/zehBKPddDSxMKvv+7tr9/I9
cGn4ZmTvZjA+akwTzggQI2j5z+bIVyB+GEHJkD0IQlo3QW8I8TtbaORsxJ+I0dYgIGIuBgaM52ex
NJRYdq5UjD2az18bC5S/F9yORDan/JZhOPmPIDhodW0mxtOmS4qZU/PyUV+BWYgwgBlOHuhvho1g
xOh6H+Uzic5NBuenBAVht6hythU05lLAgeoXNvxXcn2z/ZtLXWt2LTeyTSi3gVGkEdDZWo5j7Y1d
eJ8cnptV7zRsMUnTpMV9VpPwICupXeycM25Fh33dinsbrLQTJK7SvmyRr0OkYMohUXNEBiKEmYrv
exFAHCAQ7QNYqdEDj1szv3JXkoRwO6n79uwTe6VR7Pr12kiTPSbCBTaos5EsE+IjE7viVbbHGWuk
0OK41g4PWONOa4edCqglMCCx39ERc/yRIAuGKiZECgn33pNsc/AAlDpRmyXVaqNFB9PGCa++Xwaf
mKkaEydpB7XJJ3CA5gIaXBtrexTiSdDQM7GsM+TYryE2+s68HG99G/WcH3ro+5gH1BS9R/7QeIsG
oJQjCpd0vCu+LcaAxOf36JgUus4J35uF8hhG2BpD/IpRqylN/i9bFEHKihO09xjq37e0GxZBhcrm
L/DCYMfFsddaOPozmDMHI8COcHzsAy2uwNpfNifFhqCKBd8cUtLzWKcuyfZt4nv99H2325tUIwXS
jXDibKcrF26Fa0uCn9priLQqcVNzMtJI8llqg2fTYJCP8kLSz6brbnmKk7UUZsyT2PWj0uhQjejK
F7+uTTs84/7YDTxsZHFFDAhJ6J4k92zOZqV8wxnOyL3utog17aMDd7I3JYvr4wr8e4rC+l+f0hK2
Bm/WxyVygxbYXC8z6T/MG4Ym11ma4Tysj97SOatx+l6ja7etTIvVNlieV+S6RoBNXTlDIIgMkLV2
ifTXgK0z/KBKIFWoCj0hBj4jrTIAWWfO6P66ZKDpS0E0K/5RJfjVtiutVI6DTIt9cFA/W1Yeyp/c
aN3bQ1Rcu7+zQtiywANJOik1ew6HS/G/3jZhwmDl4tEEh2Xg7E4waernOSCmUa8twv0/RkboSrP2
5fIFH/2ozeZ4MKhx1WY6RBKG5UQIa9ciN/U8oYtUCksICZQD7EzyGeIlGCeb5w5LnLiaaacvD953
n2yZxe3kp3Hp/G0reX8xDyCNrHgtUkQryUiVGueeyMP8Q7ECFv87YSdH3+iccol0sAu4t2mGOG9P
8W9gwcyPcdufhMp4tB54HJfwbkLTqTgPeTUqHrpCWZT3cvHOz1CxUlxzwFH6QMgzTbnTmL4xSppt
+YMqpHINX/CsCiTUEMB2ntyIGVN/PAgwK5dUMPJFn5Zr9E79NGgn8/FoAZMwnz7xPI3gW5jecOJc
W4lziF4ncroja6xm8TXpcD/RDW7c9MmhPtsoGHA4Fnu6b3u9YzbA0Z2p1mjhDbIL2JAorlWFtZNh
LNQDAszI8rOMn54F2T6xTbOv1xhIblNs0hKme31Mq3jcxK9F1NdAk4UxFzdjEQhgpbLtMBL+jITP
5WuWxdwiJ7NPb+JIrNtgG2UGHA84S4KcHPO8Nvt6jR4qKQoetszwI8LoXykEYRZx6CmFxjBH4TyB
FbgjkF9LnGZ2pSRyMEXuzT5904mk+IFTL4O4hDQ3F9iA72kyWJm+iN7PYMwxT8l24mtu21xZX9Xx
+h+OF+kC+ImfHOJxJ2JTy5TvUfnjzTiTNKpmWvIBYUIQUpJq903U9FYU/0/AOkvNhFH6UoBt2rPV
TWtRmagkg8J+c7KMRRsShA0uKNBKndW7SmXURa8UGa/ISaAqmFF0u/wQGac88FWuxyuzmSYgVqqh
S31KN7PZKRAn9pzb4XU0oMs4L5ySDOOnHL3/grFbMZ/U2bihpX4AzI1jUt1lozHx8YMTDF2XDNyb
IJo0r+Kc91qU5sYxmqD4db74kf5+B+nCAx/KwmzIU2NopSCMKyIiR2IJZsJBj88Ovz/1w1zHeHXx
FwC7R1/BEeYk9TeUccLeAVkk8RTBlJFs/vvA2dwEH2UBbaP3AHSyyDLw70oI/Zp7P0ECqmtfJwln
lm+vJZ0oisOgdN5Uikp1ko7YBXnqmfBT5+UWrlT0gqx/DC+KY1HTvAjaNiqCERonfHxUARUEIdww
zNu4fiWjhVAK6WdyF6e0KlE9Iet8iAzxiEKyF5jkheXpjcWJs0CK4cIS2aHV2sNMqkSkMaiSKup/
cGSbUg2LGOvtzag68Ak/EqxNcbkmVIW42f6KAHm6sIAL2YI+tvzGKL4VRfd6++Qg7ZegV5a0r0yX
fO+nquvR4walieOMrK358ga9uj87GqHtuBUJxNyGuf6Q6s5oCqM3UIB/y3fc3/TnwhyfWTI9a2EB
oO8hqpu9n3tUq+CuIcsLbkqpQx0ycIqEG+8h1j+2mhl1Fei6qLBRkjoKDqaUhLOxf0o7gw5jw9Ye
6HRKlpaWV7VjX03wEiJ48mjiOr1qsB7V8rjzp6Pw3qM1KUpOO1d9RPVyytw9r4uAJs2z8aZZN91i
wMpAT41ueRIC1tAhQ2cMxn+eK8R6ubdRcE+L7BDRPAf+453gvZQQK6P9bu/DFvBqIgdJ+rE5lqur
coHc04GX9ECqeRGemFZ0vb1ViIKUmIGLM2e2VYtbLj8Mxftbf858duiWKvNhJJNgiwA9mxUO1euD
u8JUXfltQxWvn8O2NwoRECW151CBNb8M9fBil22gA9IpBXeHZth/o16/m15zSGLCYDoU6aS/dzSA
UTuU7D5Op5UByxXNCepXSZJD9GLvYyvcYcAZ5LRdwPCM7wKl3b8Y5zeVoRCK8EKFPzBiVyBz9nsb
mZ4sUDHxc/hew0eoy/FV8u2l6MMtq/+Mb3AvWEA9B3PvqJKyeGlc1e2Pmp31jI5CoU04UOR3DvyZ
t1924Prvaes8E7PJwnC4H2h1nehzg3O6AytyT6f4y7qyLYLVL0bcED1O/dRiVeQPHB8yS40sVwf8
REWyZGguucm14V2tqlToKIOcpPyxqyvDcF5lBP3NCabiqSeQZixNN/Rc0vCEw5BZqwmzZ9UZLFfj
a2zYSl9JyL6Bd9heSvmsQCz008QrCS/mpWRleAD677i4wDH9UPVCagntS/99GHe31I6in7KGhCYQ
xr+xM+JtT1YfLhVJTMH08FvPKYT+Oq/339MpKXUfoCdPPuG2SKzXls198fMo7RMLsVXFl5HKkbhJ
h+t4XQcJD1IqL5IFzDDd4KzWEr/rUV7mkp1lorqk6DKTmLlIWJy4LV7CoCaDc2ol/7UOnw8QmfIj
6rU1nPDxp167y+5KlDUIJGFgxmj9lXaafVXL6FyF/5jrJZGDI2N0GS6Vf0iu4Mw3qcs+4+GGrHin
uQYF7J8rHdsj1EncQiv1wgqRrC6XENWTC+TixFBw2K5m0juFuEkv67dT4dFdRnF0rBLWXGdMxE+S
4cwygoZ2ql166a1UIq9AmxYE3jpHCBaAAnyuLvsGW3XiHj8vAJxnKVUgTPiApEK0zWEYg0h9kyym
cGk1GAdY297dSieyj/B7Qmp0R+XFo1D0ary6mZR86f+GzL4ID/68eHPTXBEnNszOUZ7yzPSJ25VD
AAvjGOXotgNNxx7GoJNyFEKjQ/U6TGoUtjczPLaAFqkS0zoD0s7O/eC9CesrGPtsEbKDLYJitE55
gYN1Kdh26pJ6E0aZYoOiHniFBwK6Ufc+L2EvaLK+KdFQKSYUdNIfIz3w0QEmr4x/NVk9a7EKG158
RcpHp4a7anV7QVuMw2j1qel5udBy5V8hw4qYahXx70EB0S1EAt+NVQ6oM65YIsd4rfRVgiPPkW1J
gJuJxZ7lHHAcS4U3Ha0k8dRwpUrqnJE+G1XfPbeCrJEMMlgP3kO+gX4S/P+ozPvpA6+pxJivPwOQ
J8Em7oPY2cgbgC5zjRS7hnaiBCv+d0sxXfQul4VHWIFWxGhkMMAe/2Ubvyuk/+Mg+V2zveIdvJ9j
3ER0dZMSlNt/Qdy4q724+5oVHObaBMXKOrhAK3lOjPhrt9Tm/8cnnMPcoSfZw4yMWPB1i37BVsDv
x+1Zzo0fAU9HPTuUx37laGuq8bfxYbiPB5bR+r43N6NHq9Cib+CN5fCqiVZMro9qQirrVgNxwH89
LmtT0aDvNVQEx1REyPxrC7eZcyNiHkR7V+0sG2MMIhV2NZ1xV+d7o3yShvMlCnkC0d2vV1ZdTrp+
ti5MFvnUL5eSmhn0X9PnRiEGaly/m/L5U0s0zNaeai9cA8UWw18WJPg3OYIWRlaMYfN/ALUV88Ey
KjOKTEjhNiSFjaFW8xBwreRDW84fnw+HgJLW9bFqQwHKDmd/iEphSqy0Nt1zdZl41MirldVwze90
y0FdI//SrPdcRBLSURXevuQTrYrz10uM+7E7equtZSSseyheqxJOdSEQQFfCnt0IykL2WyyWNCGi
mJ08PvYPQWJu/G/7d2Ran3wtj+Qjme2LLxwKMp13aNwm2weI7SOd0W5R281//WhvaL7XtW/jBsbG
N/C8g3iSnUcdAstC8LWpwQzMa1+lqAu8FBwg05nYYNyodu+vvPwR1ytoTsxztrVyFm4tT6t6hv5B
QLOPNVBaPtRWZi5tIaWMtMToVfRlI9pJkwV+A/l2So0kpESgEMP/G9ukto/ijl0KbbN5Yw+4WLB5
NAfZ4SvgHX8UfNkPDIuz+vYcufwH1PIiM7Akpu/hZjhDBAs4S8N1q+lOsg9F5KEO853GmEPI+4Cx
1Uso/pe7LJ0n/2iHnauQXVu4I3rWHmNaRyDzpVubIKkWW5QABjIXMA5fkHi+cvIt0eSz6UMexAEK
MQpzJV0hMICqXR4a8CeAxICSArsr/ziOcMUBlTcSXLYYtBxjB4Z9uEMaV2xGDHSgJzxUgz+dPyIw
R5BVz9bj8w+eMx+ZSbElEgYl2ipC1X/O366+ElyZTTpP1ZMqjr/PxSK1rFqVymKV+gmh+PGoPlxR
OaoFSc1V7T/Ye9G4RLZg+14pp6l6h+WD6fJx8+fnr5jUuv3sNMKRwjbZmNJLz13YEgjSqMo6aC8+
5A3AUqH9oVNuZArRFVoD/ne+H7dgt/xDq+ztFJVMv2UH9fVU3zTJYHpTH06l1xUqljI9pTeQBscJ
HHRa0DaTcpnh1Z8QjeU7Tpu47XFgeoEeQFie5DczaXngVsHDdo+E5DoNoMiwcdlEguWuqSGB/OqT
Wlgw0seLmJ5IWTfm5IMXK5+qQyNRWlX1M7ehHZh2AaVCpc73qh8yeUbLdeZ2tdVEZHEqeYVIJQJz
cUa5k8npr0OsmdhSsEpGEqsls4mfv5zLg0qh8G4Q27UFG2wCnDzo4yhnwl2w9uQxUX1mTKNOXH2A
dWmJ9ZuFF/Po4RqGDxEXeblWtL5X8xCnVpuv6YB685SjJ53n09Nbsj38e9An7MUGQQpY2RnxnDU3
nGorZHvfTBOYHVJIeEwdhNPbsoTvixTH1cTJ1AhHd+sL2mdRJl4mg1b+F0chy9S1HB8+L1V4U0T0
1yXN1ieu5pfV318w76a/40CNQTTntfNlrBGqeCinyS7FQWlrrU4bl4V/gdlMqbkuEidW7tJ6jmOT
fA8uZ9AR0wNwIL62aNApR30+09iD2PuKSFsY/k/Z7gA28zMUbOZL95PUU5szGRTD8r0fyxzNe1ye
qC6mkzgl+c+/PJ7UO0kOOIO8hYwcgwi+3E79Nvg8RHwwj21ORseQgZ5LkTxOqGIcpY7HYQDAmHku
4lpuz/ysypmwyamLR2dnfv36CYHDR93A355JUn/79fDuBHaoDgCdl6BX3oBu3kV5KkcIvPbx6MKW
8kRkdQOECoPkXRZGln8koH9j7u3TLQDMVktmEhyhlpdRP37YD8YAcNlGTRYZ/LX1XJFRjfABLqn8
sivkYIvA0SjwPj2yIpPzLivu2+UPoEKgGuUQcrK7/gIxYkw13swpipBS4MD8DpGG3W2S+CrKtLPa
D9B07S//d9N5fUN9VqBtk1ewDW9QB1TSFym9NSM3py8oY8IBq/0TttKtK/DxRcqgzwZGMkgXRCuB
4AYKYrBzKh8LF09rzlLRJgPhRBIhyNcDrd4usSQFE73eK4qLbKN1XbU9hLZ8tNJGXJYkdgsXSEUJ
La8X9qEUWdN7pCJQZ0+o/eFsraRBA2bOv9asOdojuOnjLr2RnIAa6LckK7YF5l7M7wrq7KhUMKMo
699N0TmeNeLnB8ho2Y02VW1b7E8K4EdDgiqi6iT3/KZr6DJcjHkH4sVN4AAtnJfVGO9AZ8XIK4kU
LXZ8M2V2kqc9U6zv9S504q19KlHkwWq1CYQSFL+swAWd2H/Pqm6KHdKxj6hEO+WDYBacU6Z3MG0X
NxtOXAdp4UZXQpBbUmaqDajHJAhPBbBKc1BvERy2s6NWHTeWs2MRF0A47H7XeP9nV9HjyJdhZfwj
VeWrjyvtMTI0a7QoC6ZavuJfoSEPkcM+Ifc3z+ABAAeHVkxCJHXwMdRA/2VUftsNKYP3Xg0y8DqY
Q7XWZZKSm/LHntZvdEdI+4Zw9x9lo04J3Des/c18kY705RIdvQ/6qL88effpq6pBz8PoeVzvLFg9
KHa0E+cZqfj181igx17h6/8uTViMZn1lL7ZQNknFRItQmmYDLg3MpuHuuUmCYthlALWE1HIKs/xc
87hhGFT2axC5uvYGuIjtMRkLx32Pqw11pKcSd10BxQ9U8oYMZYVLHYj8FruSv4XXNwoszYYZSkc0
Qbu2loLOBFS3hrTnEiIMtiKbf3qaV2Ibb9Aqt2JeoY9pMtQIP3oQc8x2KVa9epyyfEL2gGkzFhLd
VCnZz9ZPqyzj4eCOyJIsDEvsu2C7B4ctTz3XnP310P0d88ssfuXTz8DN9uGrxQN/rHquRwr8QX/u
Q3Znq+rpuAB4jnY+elxlhfeuNQJPmrOlSSzTgDTDw+f3nbIQAalgWrmZ3gqP0QXynnQf2KmwjQPe
Gy0qLI3WR6K6Uy1obfjdjGMgPLRHBmDQo709nI5KAFKD1ry2ucSvi1FOMwEDBbEU5dZQE0bNA+GY
YKvdl4fqFszDCzF1z/s904vumHz3R1yQ4pi4RHXm2N1/JYhyIGgWhxSyGvFb5bancilyyfqmmix4
cIO3P+06hJ4/uGEbx7g2XTSjmIwNb9tyYmwkX1KWoiOCNCZRdeOWYo4x+bLnkg4yLg0gZ9FvZPpc
P7q0JpGllMZdUpTKntWRbi8sN4oNVks4PZALoKhxBcmVdvqe4fU3topZEOeI5ZenPkzAoZSd563W
K3lQlPUJIvLRoLixPAVvq6HOcBgl3r7F6TXs4w8yn3p0RQwRa7QDJzANv/PukfbzlT7Q+sBJ2cCa
aoz7gh1+uCRrF1Rt6lq83bCqqvaPANiRNJYiy+lOTyQzgIfTWG3CdulWaEYfTaN/HgDhL9IE/mqH
3STGvpkxnyz7pLnU6kyHFqF79FBMQf+ZR9nxre4b33I744aq98apX+EOD0nV8vnlbMukaUWfksZj
nO0rbefc6vmGkxj5a2AVtWCFjokg4mpw1AL3Jje/vjDfYtCMVirPDWNHFy817AS/nwo42XYxJS/E
fp9goRMIHEydDDJImZ4SNl5xHW6oSaP2ivgl64/3HM+tgAGyz51KQ8bvIuiNPSvrisiHH6RjefZx
EEZrfRcAVTof8oJwwuYrNLi2y2IxZH4u77YleEOwGfqc4tJVNSpMYh49Ru8oZOTfLIPI9/pYnxkn
EI01QRigPnVXjw1NxssfJ+ZZypmWyQPpELD2f2jEQ1zuFGQXfuJiOCOnVD4joDkkq6J7QxIp/gDJ
7xiGYU620e0QZy7cXs6+SoMDv93xqmxPzI4C6XQcqOosla7/RE+jcgVHR8kc26m77F5sKUxvIoy9
LzmoK+RJc/eHN4av+W8oPOjexsPWgGiZ4APoKKNyzwiusG348jrj7rF2J6ZtCI4ll+DK/hiejr/E
pGsoX7uBFv47hNklmpJzD7tQ38qVB+pEw1Kb/7u+/C6xYCijeBPDpP5EznO9nSH7vI4QJ2yZH3iQ
fnqhKLdDBZsEBE0dK80ZNwhMs4Ezh19rHsfeuqe+eRCQYWdyW1ZvoHBKfxPeK90l/bjPNN1ApwYT
nH32z2XX1K34GPGExExWsP7rQNaf2ydTIHTfcDU8KeAYR/EQX+42NgcFiChwKIlVbvm4thp6wKBe
XRdQlRCcziY5KGyBOB0jr4YBSrHU4Z3ja1moB92F6uqKhVle5BeD7Nc097Vq+Pomgm8IhOWOhiit
BWoHrGIrJnIVHfu3gS+lvv6qyvxyZFB1+fPovCDoXkQ8uDwgvLirMeUzd/DDxFlWqsj58fkfdt6/
/UEFJaf8C+4Xt/PqXRPhp9LKD3zaiKJX9CFSVFWMuKY0fniFR5zOrbX2tUkrh3NDzDSkRctIgyjl
DvTjbCcR0t9UuSNTCevoW76w+yk2CFNo7wDwBI3ClQWRxkN1g1iDfOr/v3MhYe9RRzmL28S5h1Om
UjMaHj1jbD+7KJNka5SaNBVoMcnEqJH2cVoxnEWz/cBJt5gkNn4X3b3kq5VSqFBom5Vr7ZaA8lb5
AYx79jiW10sfgsGcLByOoIG0cxgWsP7QBdQkH4OWkMm6W2Q9o6oFlUy+nqNVlONR8WSZzXRR9nGL
cv31DCEB5lqWyDBzjgjqPhF7jb2oNU1yksWLtnFVrrt1C+OtkGMyo39+9iTYLbslSjPhHho+8zm3
kJEDY65Z+PFBlmgjqZuzhOiJ7kyXTTD2XN0OiXJgmkuK335p+8q94OHxTAguAli1WBST9c2s2HyN
wn4XogKYjDaXifQ3WPEz29rD2JIfWO8I4Tp6rwfu8I7BQ9WX1woqf9H/rZE8CG05R1ghbiPx7uLW
ndv5NNqL70xW5cwHLCczZJviWpDBb1xtR64JQw2JQKHbirZiXlZv8yqQQmShWTcoUeMyGpL9r4Nj
MsxgipaIk8KGyhbA45bKdWjRsADrp3FWW+WFQaC4/lr0EaSfO3vuuRsfzMxewEtC/shgapQRWK3U
9fhuMHjYwv0zb5TGen6lE4NkKWKzuKsYlDro/eerRAZeweiCGo2wST85a8CeAO1qkTm7GV1YorK0
XsaZYant3Q4PBD69kwd2Xo12mpJd2g4FCtffL3hm13rfClx6cyYWDLzqWHH2ZjpWLYCG0wrCvvOe
2+eXNZRkXPqmH8+dN/2LOSMFBbm5lenVRNysfY2ttmqLN8W/jwq90GjNoBOEVMyI8WiQpsxAIlKy
d0W0iaenV/23tyDLjmkdMpKVz66uj0kxaqsq+BEtbO82HG8H4hjRIMibYHX93TPvmYIzz6k11f3e
PccoZvrsZ1Kuz645Mi+f2m8MjNPa4vaBni8daaWZuS4dRnSB/Dy9tqGWNU9AUGc5V+cV3k5iN9ww
PIXwEYZrehPU7q7EplzlawXaP+sEVgAvEKlrPHV2IABPnwnUm1DmVxrSdlcCJqHrn1OHW2kgO3SH
w8IoXiUZFBSluz8qt/EO6je1Euz33jQBSgG62k0XEmIEZ3/jPGpEuPLzkIXqawEPcAfEX6AZDqEn
zkc383HCY8cLmsAfRljqcWzAtNBd5eGxdmkSjldm7s421fBEJoZWBi+0IKtucvoC1xLXbu1RsMD3
8viFrXQxpANeOUks3uaERPJ5u9ekzoTaiBuHCt4fkaHdMR7qMUdVN5gCfGI5PjCyL7JuJcyJnKdV
lufPryaX3rmlepWpN438nE1s7fmNmBfDElG1a32PZa5DjHmpqe6UMAZ8PQqaQ0Tc6eKnEDJAa+KB
zfAeSlOeCrrLjHm/NMit8xT+nxc8VoYfgm3LoDF1ks8141I9j6c+06UjV4v7u9k+1BowSqGZvgsy
QYsJOXPBsptzbUtSbzsBpQ6XFq1p3urRn+V/OpLDMJSQC7si3KgYVSaXo5uYwkrIz1rKYLMBUkzR
uPYTkXKVeIOjiFfHVZ785kYNA3D43jPG6JvAcMn18zrj+YIoY8svtz7hA2itQddLy5zyW7dUKhy2
/f+WfDZkDQpK4LYDOR8LO7S9xXYytHN2vER5SPVd6P0Dr1DdsX/l6UQUT5GkXKA78Y/3nsdLq1JL
a7yxUhmmJ6eT3/ya1qIvXjAQMkKfUTpQIgvvf8a4WgZNhG+3KY/8TF4Gd8ertJx03T0vPV0oFL/8
xqdQIqn1kQzsZ1CrR1y1iQUcCFaU29WsH7QvWNZtNW3/r7onaUYF2mWBgxCZWkdVNC7zSl31nIQp
laYXzR75LsgmrWZ5ZFvYJBoKFOFoCSOq4FRvr/mgLvBusIAtf4ZrxfG2D0j0ymDwGsnEiwjRkgP6
T18LQSg6/CdPsqCuVMhuDElkZ0dyTnRcfmIGEeo2rYdqNGG11lQYgZL6QoExfTsdeq2YPkZbOXPS
rsAx5nrSAKT1MbrWMO08fDKG1mRxMBkKx34WrrqUpIY028GXgb7hMRTTDPvzK5bNWnjkXoSylSJu
vlQYrgeSDXl6ktP0f6fyY3SSC1fn+dsr+x1AbgnnjEYJsXwBLcQVWmAtkpjvb6j49vFyFgyFagX1
p+bIv+n7ykngFExrBhk3tQLiyS71WMOY2ZJDnfjX/koo/N9RPTMn9lGfMhhLBGyaFQbdCb8ZyWMX
wu1Z8hVPVESzG3M2dzolQlfyuYIjN6gSlA7KrCcHJuP10xNiD/nMEDr7d0g0I9ccdsp9y6ZQHdzO
OkWihDDZCM2xQaqbr/teD2oEf6e6OjxBt9IS0lEcrmt2zi2tdbe/5mnf8Tj8vfoyPILt5dJq80/Z
IueYYrNX6AjJFGcnO0r5B0GH19RRucGTfKxKXb1myw9TfDWp0vfhUxm3W2t3+c/JEFY6hdKPbkCs
h+5XphrZwCbP0ozq8TH2jQ1jgp5xFS1lc7btyGEAltxuQ/z2T3A7FTr00DNGRvfPOk368wGoqIX0
YDWxy8j9G42RAbtHlyNRyOlQd3YdH4x9qOilTOoJCjAnD4DHgN94imTITFo+Fe66X+imLD5Rv0gx
y8wAhX7mLzJlC9Yhcxb0kmgiPGS4wUs8dTAMgy+THliqZDUkbS6tdNlQ5dn0L0VARfV86VCX5//3
4VdjDtiUgN1qhEdIGvBFLN7ipmkDpFMVMEOCoGfPdytiWrF+u2phwRCSejVvf//49jfX3+2JEemg
KOn5anYQdkv6W+19sqvVRbtH5Zc/6kdbpgQl4Ggw0A1OnuI1vjGYITA+7bAbMsnI05rwqfwOAH+u
MkSi2IxopbDwMS4SbWfWelmNBohl3bSoiEUVhUXJEu3V25VAugANCfSgXtUK7jBlqxgM8CyvqR9p
5CiqR+g9ncjaWKq9vw4wM37NFYAY+bVtgh0SH6ZNOKRUG4N5SHvfB139CavimKavNF3QXCvBDzXZ
h+jWl2VBzZrtZdeLyFYithmp4hAujKn7o6s313IsLf+FdU/kDgZ4IBpJTon6lEiY4MwHBOU+oxrc
mxFeGAUyB8jsnhw4Zfi1/g36wKv2wIusdJNUvxBc+POaKqrIkzes1Hsk5HjjpEBK1TxzzxDVsQGK
NUODt/VzNF95Li/2SXE1L6XF2JJ8VDi89fggsdaIG2hcUX3ohkslzCuI2FNyG/tioUk6Up0HDj5o
ZUMCNc81IgWq0cYjG32+2xokwfT87qg6///L6e0KemKMxHTTnocN9m0A/lHBcTAfeklySbYLo80M
6BFVA7K+xNmtkieB4N363XCBQjdJ4XBlLT+Nutcs6PSz7OHi0cC5l+dZ7+Hg2V515OgLNwQOG32V
j6kaMlMtVUkrCd7nkkS83uRBX2xHK1yyaTJHND83JN+42TeRhhMZG4+0Uqp4ptqsfRP3cm58sstg
7XjTLwuiVOJFrE5DbGroEOn/8lcHNk9tddHBvxOkDz9y4g6u0C+Whp9YmmEBcg0x4FE5iaiAH222
MX/qB5SPCS31W49VNOdGeBWB1v6V1t5JfaePrXWrrlrXR1Tz3VIN3e4Zl43AY8jEyhi6HFLBxxPX
RY5z7cZiUKuuqBLXFVVSqaKrOnWQRzow9NVlM2RA352pJR8QJtXdceQLilE640fQkPMwNnx6ATKZ
PJ2su7LWCOPhcFZgybA4yh1kYtGmTmotHgniiaQ63zCneKIueRl7anFRrvLOHlQF8BhTC3j903SL
T39V0mULL8QAc40DT6I6JdpIxiX2HqE7Mi67sYvSMMaSvt5DkVOxaf/iOTh8vusjC8Z83NIVkpH/
3jQ56tnh7Zqevs6uJs/A3TiS9RJxWT8A/9BAUroeCGrUAG/oY3uZYlFF8OS1rIADAWBgbwrivq9j
6SLb7suzVcZNmF1VRBA7qzSwfiZkAMLofO5zKa+RMa2fyvHc87pKMB43RuI15UoJcggxB2+kHVJF
BsWwYoKCjfQqWm2T4cyM3Lsh0niT4IorwlWj03LHcxahgfeWtjU2i0cL+x5p7Tz333l+UNJfb9Fo
Z/ybQ/SfCRmiyhHukJzCJ7IqXr23RN1QYBJsZW9zMsMl/sNjomVJED5eX86OMhC1qZFvrUVQ9oWM
th1WVvCmeqYMFfINGz8W8+kXmSRU0/mCKEFOhxYXbh8MiOhwdL7naWriELOExlUnwSeKqzQZKJFw
7+wH40YdTnh+lnL/J+00w+qT+//e+CSujuGkgtOpgE5epx9u8mMCotDCwLB3y9OTyO7SuU2ABiAb
tMPHS3FXkrkAU+pN/Fn9jqs3ckMnBbsmhSVIRJ4pS/PECTZSQ5CPSHxDIlAM8RzoJmxlnoj9sG7e
wLWbC6l06a92MT5NuSyULBHIbq9LK/VGitrACE7vWNG9BsPJh5e6NHn2ST2mSOFpJ9m6fkS87ixt
O4MX1MeQdlgs/b50ZhmnpYuiiIiQlF0bL4yoB583sMGqN1B2LjkFAlaiPDcawKSBblJPzseEA0hV
cjE+nFWbrLPcGrBxkAlyTizwR+AKCuVgempvH1clNjxaug5D5MuuP7wy5dhnWFdOGZfM0oGUhkuo
wMhmwEZ9IqnCtH9eM49Yoro73tC5mLyr1U/MCS8MQ+ae7899b+F5JYwTKJUNqJqlPcixq8NOVOVc
nvIHObt7feG6VnG5QVbOK/+5q2IfzQE/23mTbMQJ1VmYgQMkkUPee5c7+jzdEKOlHigOPaKOJGb/
7eZRNlbp5yraywJXPhqQcsx3FsmzdCbQlqPbpeyjmSsVEoXiYeJ/0tcj5aPW+NVfY2zsO0GhGeLp
EiaFRGyXQh78SUBpDOMcvDY8slIg0WHP4E/0Dwsu/J8ejNyucoBVmU6Zadmz0AJXPBJ3P/3YJM1p
WD5oCjTdUfZBX9IP9HMEMAXZJz9yV9CX5wQ+2blytNVPLAj5Mr/44M+g2a/ukC3B6tB4d0cfyY1X
hR1GAApdVpdj4NjGPL5IhFm+VzxcwciRUQWzMLv9ZJBkPPv15lSXJhofPdPTcHkyq/uGP0NvwMiT
wsk8erTeL+lv7EvBKzuSw7JxaRSV+23fOdoOgoBXY9NI4PRo0t354+BHYDSEAyPt3iEIgC8Yuo4q
eZQ12KtVxvTNEOReXkOUYl/ptDBMnNYnOV0UFAzu0Jl8VVLqkcyYoy6FmtmAxq7bnF0a33yX5uKx
csuIjtBhvXCIcRiF7R/gQWhD2ZQZ0RbUBMHAjTpPRd+4hCzWF2oZUPUBo8Rp9M6JolPB8vStDthU
GgACtxVMr4Gz4ZjKpxUWQ11XBuBrt1TFCWVdbN7vEy8dHGuaInZ/o2Purto9ByujNZYhFJDDWKuq
sSoJ4n6ceFyyW8dg+tvR+rZ6IHC0LkzghdkMv21+2OzY5vKQirqSeS6a2SRO0XBQ1Mzo9w9XAuLR
EAr38YvsjRfmiJ0K8SUG+l6r0ifuTW2cc2UhHM4xAQ0cQvcywndSgB8eaEh7AiarGfBom3DG96By
NqECZLPg/fWzZm9lcffvf+qJeJoeU+8aPBDueEuDrjclpWe090bXwC5b1wKzO7XdeKRQBKf6+FuC
n5NiZrBYq09o5aqYUTwEHUZCmCb3iQ+C7S91ecoJ1bHit9765t+XsxPc7ewRYtRXbNP5Sfa+dVcZ
LR5IhIxBpmexAntYK51S58TPYTtUkrJZUdf3PkP+ge8aUtxtwaAZdt+2xnxy9hCFN6ZASz97G8RQ
oLQ+OygVhQ3pn+gQOmQ1hv43SqMGeEkiMycniESuFoAf9WJB4dxf8tKKIU7vLpgQExpo8SAKmgRj
riQPhRZhLbyWJBtlwDf6igfY39HKo4srhzGGiA0J82lAUhVIcGe7axt9SmJzlOiXghXX2gCMxk+Q
MHxfELaal6rtMD2O31M9AAiro363yRpfub4dMRIJ1y+Cgae/xXe7mbMLdnl7aHXqfcDEliWaO5bU
0eKIgXBeQMx6sCq9BzLTz5swiiph5S+OaZXAmFDtdj1PRoTJypeQtDgpHKh9EpWqQrp/MOFoXvG0
9K4EeUEBkQYlypiAgbV6ZvH4xkb57srDLkTdd0SNY3nWMgAGx7lrkza2xGn8RJgw4YfBh64Ap4ya
XgvZFtnzXjw/Os5On2DfQ5GjuFfD3dfoufzCjRrG+s1/AEHv8rfn3fXsLzW44Gh5Fl94aUC1exUX
DaGcX9ifUHDfPP/9OhCHrT3fNE4/B/2NqSDCe1EkXc/gRqHaYa9SNTMH1PeZ2iucJRgEut7kzM2t
yFJ7Rk/yl+Wy1F5rflp6JCGqB6ckuRKQIpPzdhb49fU5V5a3ZkZDKVkpUqOcToMEm9Pc6rGgh86k
EYnfqYGYqAiTDVTHHP+KbltrIKQ0LFZJgdqV0P3f2GORA2luMXpuBIG7d1/+3iI/VwGzLx6y7zXh
vJioG/SiEUlC7yCnE+ZLspGWmpwbSOCYClT/M7xVYFV76hGz+hCmpXELTmT9Ac22/WuPve5C5vOi
8FpXYiXGI8qvetqoQf679Vt6XiqSDy7PZQe/ch+EIK5eag+TBfbklITbl6jrVzynN1K2ZhWgXS9y
vIUS6KW+Ko017nyBDVxzq6M66ncCi17+6otXnafO9XzDsQr3F85U0Vo17JzrbpnG6gvRSbhVbfwa
f+7dNZ4jUYdZBNuoFV7J/Mn+k7bzjPropIT3QO5o2XptnpA7av704daJGa/nNce6Eh/JEYBEqM9N
Fo8ggp371sehn3/9Z01/T3/qp6pIg+hGh0tVCelZIvIdPHp/bS9wpN3cOhYiMpWeCe1DE3vBKCCM
pjsAXRNpYwmMk4K8Qwkr2wbWWR7/BmHTqSRy4lgaKuqpvDP3G1oo+X4N+ffrYumETLvKMIWxJTNJ
Pes1GRmcmwfzwUCSkfJebWojRX1uFqXk3CznIwyjiMj/oI5xsIRRmCnOlFh3R/FnRxQstAXBVPwh
cIQPBMe6AwmIdA7SN9U/zXLilpMobpSQWJqGc4pmvN4upl2KDbnJ1fqRb/fZyuCrwyQ9yBoufDeE
zJJXhk6OXboQDVyjbmV1lh++H5RLb4MlsOaPxzIgNJNQkfZ+CUxaDIOD1XHQdUAkGu4BriLekr3t
yQHzw2ArnH5e75ke701NRyBx3kNAMlZ4JcOq7eB2RmEK9pJ+MkoKGunPLVOSOxstIYxMaxpT+lqI
3JAISHQuZ5w+P63cgo6DSUqtudhBDMt1VI1JXk4TSlTUpXZ+hD63NP7TAF4OjTC3ymi36dq9eOsz
29MBxEx+wCVLyhJlx8thHUu3j4X33jvTlVsWOTjqINlKqiH23I5h+fADbOQANSKzltPTa5t9alrf
MQ50I6m2dFqmt1qXzvEGfzf+isHX8z6Hfr8XdnzXEZZsVXjE7WdxvorS3DjysYXVLcow9cVn2sfC
6CmlZTW7gOnkQvCgBry7w+4pg17KJvIOYDb4Roxygo6x9MU5GZ4e4UaC/MB6iLOq6cXv3rbGbiNY
Qa/As5DSd6o6E5FaDth9YNhvl/Zmce2mjNcs0Bi62ULkuJlTpclbKy+TpyMuIK4x6fq+angLoa2R
7JynBAezm0T3PeHbvpf23bwUIIoCTe7L3W6f8IPHYwKpEJkJF92UDdBrqiMuWpZzLvUY9KSoCKtT
gRfoGR6cg+CtH3ouHAyMqCxTdcp1x4ft+fZThzl5phSwdzRv4J42wAkkEjXcaRGA67ggyxQk4Lq7
PdFwCXWVJ4ymf/84XYGvQUTqpSkuL7eI6YuQT56dksn3y2S/dql1HxqXg3BtHaHl4NcaKzlV5S/9
eh/E7P31ZsRAciDUX6HWVXwDKujDnt87rmOb+ifjQVfUXU6LPagK0b4kfQEZrSHUBtB0nFGH1KU2
xXiud1o/tXMzEUVSb/TrR8fkw8fGei5cfwAQpD+HkHk0+6jb0F2XTTy+g9dduWoSbGkfXAmjy0sL
/AjEltsUnAc1vkTnQGRCRDnnZtMXitZEolwHmTZ4BqIaGei3UXDX9aQ59G5ZJze/Qi6eAaWc9BSq
Ny2isMPz557RCW1G1Q0AnOR3o0Gs7cGC/u8Q3WEjylq5FO1EQ5xkkQJSMOvFsqWbOfwZf1ZrTH9v
xbJ0XV1NFtUFoyYHA+U8EAi1bFIt9AsiqCLQZf11iGb4Zi8tqysX4h7uPbHQEH+yhIBSuur4x1ta
OSo7mlRojTfNDebFF4JTQpwZ9TMDka6SwjrgemniWT63hVGcHvCe6W6gX0KxTPmBhYothNLd0wKA
kzyRNHe1gvVPMlcAxx6AZ3bzeTNA4so38JxGmVsUUrxRg/Bw1EXmZGRAffsRPh1vK5ZirxmZnXr/
iGxYcwK7dJUngNTX8O/BbmPTMZpgb4cG5jj9dSDcmGaxio1x15aV3aHwbb5PJpIkZ6JkQmd+iui0
TKZBDapRXUhe9Re0lRvaAKFTYKUUJ0raNq2fxsdSEqnc1n0Drkzr5jo/SYh/lvt3mMHsv8mv2LIB
jIgBuLptF5UTA8FzZdoa0f/m5cq+2rWx6LKh4mpHSqVR1Z8URypPFYrqvf6gxzKOMGPmwIbVRTx8
eUrcP+tPfuni1lJgLd0G5CoJGIDheDxtaj2PdQ5+HCMRj4gS8oajgpj7BuK+6EHjRGkq+14LX4KN
xeY982zEEQuBQAkv+nDF5Ju25kwR3wsZ9VKgirGgJ/BabNysBtVm/iby+CBzmyb+PxRiaAIKdtWb
qMjyQKgM+evH+68x1A1Nm0rkSfcpq7NwGB7/jQ6GBvM3e4kizBg6QiDzCSHGlzlHg8eHGCfKaCR1
6C71M2cWbvgw83OlOy5JbD+Q52clbhG4YR9clhXPVPEQFv8NC5wFNjlJWlAwSETdBFvq8tfubMtG
Ga+bD6/Wm41DatpFZSKrPj7N0saAAjsGT01Cy5C2rh5gD9JrE/g5KuJt9akoS/oJRNIR2hZw6rwq
GZMOOUH7bwMYoEThw/OE/K/yGnxa2z8ob3JDdBTCyKp+cHqIG3M8+N8KhyTSigqkgVFzFjmXD6jH
Y2X/bB9tmNuOWfxQwTILuCAWW4lcVpBU+YDeAmsZWgnSyGlR/8pj1R3vaI7eGbjHoVRBEp6d0vZY
TptvTfYbJ989I+kC93qbZbYILRStbt/ZuVtnsc3jk/5wArCLtlgxOiCCnA6axqBoEReQu7s4u6qN
o6/q5dUPYAm1nhAfqGDuT8vObUfWvR7afJP7cYjqXytYHjwBhzixgeXR3q17jsiBDSlClqiORWb/
S5umFRnmumeIUEUC1wisy/ud8zOYZiEJjELNSKUz+Xbx+D7+D5El458x3pLggQXcG1Bwd7ELVluJ
SrzJ14llOf4ui5AWP1inGWV/FhoEgQ68dsFhXqdOt0qnPYCn2w/q+x31t0fiIL7fL4eMHzSq8Bni
FsvZ6p98MISAx1cKEF+4lMC/Goe8b59XQq2LsJbr9Kopq4/7ynMmOHWP9m5BADU1mDpBZI/j251M
V/5MyhAh/RdW73XFA+w40TgIRFI5HQewMX3wkJWvV4fvP9iqoBE02OZ2+apUK89zWCTjJulbvrjM
lOaZDe8BBtRNCeq7Gb63UuU2HsjV5qGUCGrdiwY7EF0QtA/1sgHlhzKsHgfvRBwKX5VqGs9mlAI0
wDwflOaIcHqrOopZomLmQpZnxTnNi/zM32O3J/WP9k2bF1u0lG4z1LhgN1FB4IcsA91dBltKYU+I
67i4THLZnR8e+1ZW2e3qv9MXngN79AkAp0AA9eb3cNyYOahiG4alXrM+qYMmRjZqWWHSo8qvNv2u
lhDi7SGuUr8yMjM6Eh3amg6guaTetgNFI6hA9j89fVfg+TJlYjPe3+w4jZX1CefgpmLF1/saGjJi
HcKw3vqWDk/U6DgZ+wJZY8u6TQSwMalVRChLRD4Uvl1ILlgoQI1akENUlFWmMpd7u4tpBMH0N5HC
p9YTbidsAxtZSysB24oh4ix1gnWf0nDWAWgQYU4FbeVxo75Qa7q+iGP9kkGHELw3jszMSTtObND5
C2AUt4anaP5HTsFY8aUgGG0/nVXYOgDs4/X8XwgPwnVrYUITtJHeo9NJP5LH+g5W1u8m5zveTDrk
JE7x8Jjjyk8iEJ6OwyyduQYiDqIS7JMaFNVG/rmaL2RU3XAR18dXKc/851ZOzHnuCl4ZuOBZ5gSP
8utflnlzEzLdc8H/32kOq/k8BhxPaxU2EvRDi0lpAUrfJs44Rv1HqEgvN0+6X5DDkN6gbmiSAM1+
TCZBGCzdetEf1yYXjiG56H4u05mzzej90Jjkeuqt+YnlcZThkcwbhKIVWuZnc/xZvWYDdvEfjMP9
X6siqUs5HpCzM1mOBGYr2g7Vwklu7jqpZ3det9f67r6qMhU4jYc0ZpeSOkenw1n+d3nUoA7qasx8
B8A4xmecVNRArbfhEKCohri71lQXlazgS7fYqeuy8cmXEhKjxrsC5Crj/AXOOvGvHzTeI5RIAWM9
VgoYJkEEqHhyllMjUaxK5V7kgYLw0Efir3bfAqLOOLxisc/Ah1fGqn7eKX+XxB1Wj921yVtR3asS
+qTHPplStKFhRSpqi5kr7gmfQv5fba1xzRsYIleiqLFMTGknHpy7QM8VQUL1EDO2IPSXM7ThNAbo
G0fMBzstvWH1iAC/tlhL4TssPv0IsPFj8DVfinAjqa5A6FUQllNoCtqUW5iAROt873R0oTTNWz1B
LlOXyX1BKlIUfo1yTg+K3GeUta1Wh53Qob5dKBm0DnoumtHQS61/GslPTENE3iT9VYPsPLYvwveH
EG8DplUjnJKtMg2cit/gyUb7qeq3SGLvJ2aJLcKScGB0OiLP+5FJpZTR9wHwRU17BJMN+BSXCo+B
P8eckmJdW/G2MSPegRIb2Dqjhm7h0+Q+Fhl0T1Y1S4nyDYq16H535AER1XtAqNQp6FeMVNaaPJ7I
0VpF2H9B1x7+OedEAEQX1ud/zX3VxmSzmDQd5eluUmGUCecXDFo8xOj39ZbTZ03zwzQRj5x4caii
pxCIhtt9kSlnCsGaBhJW0dNaTkb8qZNC7ec/up8BN8ilr/BWMPV/YOGhkqwIeCyJ9U3IwGczg82n
CiXGftIt6wu+bRSVlxapgihDVWxIxU/w/Qm7COzUdS/MpX1WPSZjNCeCC3eoVh1MeaOyaAksmrc2
Nwa29/rDeiEXjQ5ygLwDfSkYdavHcP+sNRuNo86e+qez5IGlGNprfpyJRNGhNNuBuiKK5fN3p+hz
4iSTtu09tclCo5o8kjpBmDwTk7TE8TYnAMNo9RU7oEgXBCJSr6P2stdKJD69RLT2YYzT1tQwddjX
y7VDdePaIhrX+hfTw0TqYKN+pE6zxFku4bise6XmN0ToxS1VWxaJWWlnlWwumAEvfdCIkK3GlrbI
TMwtAfOu1xR1wwf+YApfbO6GjItAuoqz138ifzzhyop6d/Y5D2oBsnclf5J8NhzGktpE2ZlaPh+6
Xo8E6oagcdAqeYC9+BkYuk+52T5y4UyiaSF+6u1IJCNfJ5N0ezW9ieH6QaTSgXTmTzmcFS88sjvu
A/4ZSZRAVX4YiYxxpMWXbGrZ3gRgLtvhTDsDp68+zInrIshQt0aM7BY3A8Xbht+21rJSx3tW/4a5
qxgOHhvqe9EMkveWJjghJjvX/7NYsHoW4z5KFEH8M9RU8eAx9BSLG3t1hODLAscT1zlEAajws1hV
/3LVuseRTuD8o5QXjt6gfwFZlksqMz1nfEk3Ohhe8wozlPXd0MUrQTLsyiaHTkJmTYDYWbIiwFrr
0tKk73ERmKLjI7D2qWUcsTS/mnd21NtzAaT1oEm99YCazq8CuU1JgLeTo0fs9uJyX3tmw2m34CwK
6UtdcQmPpsmNNE386Yfiqxt0hMh26qilbaCnQWYP8x+c6kS4a6emzCLc5YqIHRZ8uGq6biyHvyAJ
KD7lWn+szJ2fVKrUbRWhhZTdk+Gu9gJHQVPqfBPScXSJWe2/Z3734rFeYrVWbyZI/eAaRDIpPTlM
KrK0CT18dnU7UOBcmLZRaRLBOeauxzeF7Id2I+U6Ca97wnN1A8edLH2hllKgVgW13PiHxMiVyZ5d
+cHw52gy3LEQ8P0z8aZK6Bsv29aTCn/eYaiCcX/6zsMbHBszGAjO731Rx3GmFfmhUgyvyoh/CsOk
9xxhdBv0hCrv2RcN5JpGhvobKTJno38vRXkP79xanFvbdTWALXkikvRJwIuyK/kD0Mwwr8bm9c4d
4+I8BMkqCSWNHAbzHMwv/23MMt5mYp3ig58c/yOtahulRfQyO1jXlbgNXLzclE2vihec84zkUBlT
X3QTD6q8jq6f7e+T9eHF0F8O6SJKSPMlD/Xjgxhwk7vftGb6ZJQsNdyhlxH+WSGK0C1WH5wmJ3PU
sC7Fg1BYTWm5tX7yY4rTBcedUnPxPk4kQC48PHsMOsZur46vD/BGbWaasArR8VnVJyB5Ld74xzvf
isYt0LfCRP4Ppsvsdb7tcn4hIfhMEXhhS1W1Ai4+GzG0aytX1xuRf6sWkE6JNLAb4JxBJyKEKAC5
DUFnT353zTC0qyupfeC+rCC+XYeYucJ+kSDfVVCYSr8K9jvo0Q0nAmO8NTzvpYgtRs7BnVRTd1Fp
kr73LQKGkkfCtcNdXtjTGSAGPNgqQxM7TvgV0TPx6Oe3LSiCAlFS/An/W6OQBVT/oQQEOcNHzIxf
qGNPu6gIGxRYLNAa3tiV2/vSkig2ko8mMf+w7mDGhaPHquVVO1xGdiCBonFTLSvWMgRLDiA9AOsk
irYfvssVn/KVrg0XuQ5RJHO5sC4o9kuRI6KRVftK8mSHS12Y5VJQtiiiQnZA9uljtIg/hVaNm11w
J0oqsofHnQLYOWTKaIbElaJ+Q/TSPAvScBl7K1+hAy7392G3hJVnZ1fLlpgbmIcUMgPQkWXJGGzv
88Ef2W+seb/bu3cgQjlAKpedQYwzQN5G4c02M8tWeqqbUDIVpM5ytfUU7tffsqJJqk9Cpchwt9xO
BNosiTuKFKQDbMbJLv3n3oBePMJE62ucFQrJuF2WiR4i+CePFtq7I0O0/IxDfMLW+sF8HPjuKesc
8BDWPDNNCvp4LQ7V4z7/Mogtu5vsocueanKqs8x0Fd6WtGWAwTU+hP2Wz+CYHH7lfp6ttGwAzi/l
0vBFGfBMHoHkUeJJ2h7iULjQZ2FdV5A/5oAxb+zzjaip2yUATMhaMx+/MSVzQg5ZOD9Cfnul+grS
egHhjabclfPXiSa9cVw2cFg2vLmAtd1F2vymlrBVuuiQ9R4gB410VA3z4ErcATnThoC+J0syFEf0
iGsNsMYInIRKHIhoJ2/2Llvnaji32FWfOMncYfaWUpj8TCO/oeK3bsAoK/P0KsKihy5xhBdGlL6C
5FfJ0N3VgdcpBwsrv4nUVbERZGb7+xwbceff1Qd7fF0Qr+5oWqobfp4yNzNbdx5e+PlfgZLqO2bT
CsS+jGni/q54HmNqgCqKieiw8DjxhiPayZP5zZLGPZ0tLr2NZrPZj7aeOtPcFcfZZF/uEgFfIRy+
oINvzIGMzp8VbCDP6lCg7O8SrESxmZVe52ZHjWplIz1iMwlDyfBqJhPy699sYi6GPTdqlea1ZaWf
UCB17EnBqloobo12m4ArqJoh5E2/UR6dpFV+wHKWws+g7P2wQNNC3u2ynAzh+3jnixIxKO1//m6X
OGMroKxSq1zx/ALjOwYG84aYoLkT0J+b96oXr3/1FOBe4ZTbbCthxTqpj8MGfBle0dC3FVUdgJWf
ddDetFk60Jx/+7Qzw7WXfxvHc2P9JKO5SpGK2gGhiPh+WXZtM5koMXZLXGH4OTWmEqFupXn9fqjE
ZKyiQ3mkeTPWausyTMul4DrODgUXM8235T5NW+wB9EckpTenaRTKPChZL9qrYYMcuuYA9FoXLyg5
ybBQf+TcVYXhYlM6wlyMt51sbwIIxZDwUinkGRxyM+4Tm9xIMfh8exwHQaEafBDFHWgFyd2p2DWo
IF786svDDMy8K+z2I9dFfeOZxi6Qg108ySu9vKIQPuf4/PxFfIgXqLUqFIaCLwY/jMiO0l4bGTAj
I3xCWTb16l2+LFQu9Ie+MLv/CsEX0fH+D++D0+OuXJCKHJfCsivMDPpeM/vG8BQ4NGqHgfQNrxnL
ajQPqoDLna7h4iVlU9fPtBlN+/+PXt8nR1Oro3SvnpzCwuXLvLNTjBm3kD/xKa17Y4AFMjOyWlTU
RVMnE56TCBMaWYCB+ejf/18kcZLx7FFa/BeA9rXY5f+wQnf1mZKSg/uKY37MEHunvzCcF0/zfE8A
lZE9ciDZi7tjtqSXiD6RVqfwqnOTGZfCXdwr0uMfXmuhhhWzwvNGGIh4X73gviRTRL8qLBfqoWy5
5t0wDP7ozTVkc9RRrxuW3KmKVfeygFqn7lTg2nglzsFfD8PqBBxeJiOJfDUb+EashgQyUHclvJEt
NfcqLcATNhTkTv6D3S/tHAnZff/MmZXa9/x8gpfAhuXnwYLpNAAXVoBeAs+0SkFCuB6jOmE2mGEC
NyFSjfwFjummHpCyTtlxEH5nIDq/fA3pQds7YYHARIsCAs6oKAxRIHD358kn+o/4cVMyO6DoITaF
VmPCNlhnupS8SCzuv98cAovHOpTY5ln4/GBeV4gofm4JMeW8q9ppPA0j06fOzdgHh9TSnycewNly
lwgzXQ87q6sGVziI6PEbWogwGlZwWFdA4z7Ka29JN5wgyhY+EI0q0ifVHQnpBRPHjpCtrqxkB/pi
Fe4G+jwWKUKNKYx+Ekl7WX5ecwh1hWWtY2W2tWKgVFee+NvSRbyfFFtxt2VQ7kJm2hixtAIz+JI/
cTkGeb2n7DigneL0KN5S9dRlcv1PuijZtNq3AkDgGHYQzgYMk4A+4vcAX5QHzlZU/T7EeatpimEG
uYFajDoeC8D/y63zWK4kDD4Gb3vD5laUi6VTXjznJjrUzb3zVvJf5WlU8Z2Tgl58eAZtlmWl/ddA
EMxORmSK95C8b3y0kUKlJcyqypQZyZrjDfGP715Rr9Rj1if+hAIaDXCBXNIOTtn1IxwBbd39e3Z1
fepGDJEYSg2U2XcL/nPZ+j4J51Xb1lXJLXJpurv7TigreagQAG9R1uworZO3kvu/cyLlJQNLIFOp
P9IllR/ejfoufoxlQ1i4ekaHDep1uRq9JIlS4hw6axjG2q1uLQXIjJI1whF02IaKBSiRzonLnDyQ
ZBDRK0JBXlkNjvZEwVmbooYkeXR+3AAFGN2WEcI0BC44o3m0/8D2YKhrhMXWVCEKpiXNBg7Gxzw0
Z5pL2RS9FzNIEQgrGDbX5cH3Q0UGEztIYiBnEixrmy5Ab9WybjaATsXKvNs+JGjFCV74rt1A7ZmD
L0yFZLjnYBmaeQ2WyNfn14GOmgNoEjPkbfXI78hFFi0+aAeyX/tCYyS8pM3d1jPoZHo80EmPU/Ul
90opy++uPk+kBN+0JqH/FB6JOtpeHg+oF9tBu2LXt5Hn31VFgA3dUA82VxHfF+vCcqgzTcK3kdmH
G26N2RymDNz16RNGh13gXMdtJ3QQ+A2DLbdLX2uyTeUIlRewGQ2RK0AM8GEtBzRh+eUByoWW//uD
JTixt6jU8i1sJN+xs0qopl6diC2tItc0vzfqV3RyPg2I8//88ZY0oi1epeTKE1lf6eFP/E7BiHZO
jDhv3a2vjDz+VYNHpYJM3fCp48i8wLjLEmKCfv2zvIS/PH9d5x/aFkM4Lf6zsW55Tg15FcM42nQJ
3cqHzmeEQU0BpjVOtISVph/CZWVuapc4YE5OqG1sBgs+crgh3mng+KT7X0vb3CMZRGH0w2scaSGt
HUsGBJlJzc9/wBi7vjA/PMrZKSdpesnet4VYPZLq56+4Lj47keWa3gBN6tkvCXDH4ksbkB4mrHWY
sB2i9fHt86iq/vs/KxhGRU0IPAWkI67y9GjA6ShEcggMVQikKzcasIfs4078xXwLB/EUXC/BvNwp
lTYXpTrkXheADImcF66aKOsdWbGwYUpUw4ZrE558HO5LdI8Zi43wlVm+S9FFMsaP0gcB+oCzdsAQ
t0Cg8Tv+lWT4wELpeJk5VvEfibvjaW0K9A8P0hPcI469g1RdwqoeRTA9ba6WX2OD2yEPt7mEvtId
pjK5C8A7HEIxP5YYUbG61vzl/gALGxdBNB7xRu9MiYRq/GJy9/DZyaB/qOONOTOxvkzT5g0EUz3o
2DVgAjXQFNz5eXlSem7w3qxoDJtrAic9crlZEvYlyKLEFcLGcedP7xijVk3qgc78jAWCIF4btZiq
j500H9+EzofqQDkmfhknoVOPF/QvZI0uRl30PgzfVHS13lr4h+BgrD4Wj/DQXPkj5EZI7Az45jQE
MhJFusgNgSBsGN4qTjbceXjS83YFaSOaAcOKSQbCDWSutbD+X8Zy2KfDhaNnn2GNwrFXZ5K1zGdt
hWIxugsNKs0UlOk5/OkwZ+QQ2MK4e4pnipxk0QAVXdCKJE5bWCd+HQ0G8bjPt8GY5ozDNnef7f6V
6ZP8OIZP+FCek0HjDm6lVmMFm5WPPzTNODB7IG+fE/foEHkc65g25v+1EXhfuYIEcePQeU92cvnq
l+AAR5WImlKATd6vQZ4ygVPdjEmNBgmrBe85jA0iiV7ULoCQHDx1CYyja16GqlgTrHCKI0szZlUm
Pu3CAJOpsZunJDw1UQBTWnKV3SOgXxSJE7roV4xiKMIYkkiSHmnKp1lwDwiRTTWbt78w3TKad1w7
nncxlDU5MNKXMFPUslnrr2FgPb4uSFC8vpHW0FgufzOdxCk37hmaANOpRgXqCyLRpgcS14rNenk2
SOOvDOfG5fKdSYRW8zGjtZL8/z7zUwh5TVSemBoIHQz6l+klCl4f7uwJv5F76mRKIYqTP8NJtE2I
itMxVDRXJyKZfbG2A7fND84Yzr55MTgVCoCAfpJHAOlwDIHvuNxx+QUGjqopxPGtkZeW02Cnxqya
VoTIDK9DL6273IDMeJ8WNWUJwdGMZAblHvAKoKet6VwFsxmjYuEZJ9LtQmz2GPME80TZ56t7UoOl
1YDsGXx7UylRk4rBXQ9VvWf+OjcrMYCIOPUP/XLiRKSENL8VRA5j9QhqFNzjcJeV1CBKzR86ibnd
2ZcFJXgOnvbcdJPl/+QEZiS4TTQZ94GuZKjBllaAMz5D81fe8ItA5Ps9sSpYgkODhrE6KiRamJFo
AIYNuIFvSnq/Yx6Dlf7Oel4Rf5nbB9kVaCEaNlY5k9vBcvsvSunmOSIZQosauzFp461eyFNedg5b
A0QnqHcZy4j4CbtcJmab9IqpbQKsjjqHtmCtDatfI6F8aVZKMUw6xZGb+q9uLrMXiXaTDyRZf3B3
5pgYdbCjk6yVsmENGh8WDjzQAOnZ7/iP4jmLxI9cBHwgo6a5VRH8M1U2tjD9/4WOeivbcjrk5JQh
Q0tavAfBl123kRsm+xUagK13AMopGStQNxRaiuvnllrBKuG6CCrpmf9jcRloBAA8cLQmZCbziIps
OIz9iiZGsIZsmRDix1ofdbdZpJhwQZibpoPAr6ocaZa+p9i0NUM4VqNAyRvD0sIR0rUyI2QgcyFC
59O+D2H9mdPEJtRZy00IgfSOLWyneXUD4O6EIKXe+PYgZcmWtI6gpKbndOUUCcFjMHOQApdOgLep
tzQuwnHXo9hnZJPQJnf+fu0Uc5TkmmnzJMAoBHXjsPIJMn4qkt8m9ZDLG69jWi2vZls5fGkHaPOb
hkdrsa4N3M2vT3Kib+oyIiTNiNw0BLSJ5xYX4nSvP90RElUcK2xBjvqImYQeRFOrKVLxfSljrAWt
/2o/p3UEpTNzbePMxtv13tfit5ZnleQof9OLHPXmhCYEeZnGuOGROT4CHA1OokzIoYW46zU7Tsb2
Fg7Jp7fmCGZrNBAi42jVbWoT4xmghaFES9cWpWQzxIaWjico4OooVNxRSXE9eWFLypr1SSlMPDc1
8SsJ+osNh9b9pFGi2YDr31LCwRkKJoopL0lMOcFfVC/gSu0wnsc0SEKza7xmUa7nidxAsALJVflI
65dq1oDS529sPZo9k69o4ParUcOV2pFbJfF42THUGHroe37jc2dO3mdcgTg2m4/Xge0Aq1RsFOyi
DHU5VqI0Bl+qiTYAq+qb0fzi+4qYj/p0Yjf/uVthz7IqoeyY5sYuCnxn3R6OqgysGGKng0i0MiJ3
KthEH3rMYSl8tfqSuDRNHQlVnpu9hlSOQQ2HwEIDXL+WeudZi3nZulkzP0CHYc0hF/Mbw5l8m59u
Una84EQlkN0h652OQ/ARUVl1sRs/16VxX+XngOdMifb562gHyElw6UMyET+MLW99xFabnvcd/xPO
fIJszrHn7FLZC6OYEb0cQGuFpUO2DqvGZEXfLF21CmEBbgHXk5ioebZIElBN+wr6z6iRvjuR1JbR
eZJmJLtiftQhJ/rIs4dH4VbEPguQbIXxDOjlQiLM1tiJFUJ7XgvLpu+R1G4sUkOqS/NXSRPrpxmi
q9Xj0QyP+0D88/ZTz1RQiI/siuTMAbdwUU3hv5sMjbmVvic4PJ+XC64qEBDmRbaHsViEnv/5zHDD
S6JPlGhYPdQh7Ossd00R2I5UXaB3Y1hlFXM8Vd0+WE4l3Ov/GGbUErdRFQsdHUTvY9/NfiNQ2C99
AWMCqlV2X4cC6UX6mAT1xX/D2m7RRuID4QNEtsQSBxwDeOzX9CxMgDgy57OSNzcVwdQYWx2ml8KL
f3TZo66mbvq0YQBlwrCjkm5gK0XQkMGczniMQuuatXZbuQEwTmJ62yyfdGgXKocDS5XgYK0wVnvn
t3bZZ8Lbq86qJAVza9kuqbUVUiBu8FJ1aldYpJ/ObBM5FNlcHVW48FETt7e5Rc2dAWhgPHS0jhrG
hd27Y5SGeVo0Ey+JPujfsDHplu33QMkE8l/0ko1t1nz+woXzy0CQtS6N+WzdiHhzJfOiY5liWn+4
irz8BH7+jdsiN8NXBlgJKkNgIxKDRLHEKix5l/Xx5p7uhpxLYccrjdyDg0NdXWndJAKtwr6br9Lt
R7Q3G4c+oq93+Z0X7YHmgZ8Rv6YjRiv/E5/YnIC/mpKS3GlOf4bPG1+0olPv0HaxmtMumnQAu8nV
FSz8cIzVdSLKF1PQjgWgCceLxbq89/H+FnYq+UXdvWmR1f2e1VB/2Fhpt5Ekkf3gFDGU3iktb0Ba
Gq/FIM/kyHMebNXf8gyXPu4ChYpsYIElJ6Vdfpqb3z1JLM5nKK47YAy669dDnPOk7TFWlFf7ZJ5t
IJWIofCVHaMftCRv21nmTRahkcuwpvIp1l7cI8cgGQyNIzATZnDNdK4Zi3MY4Ri3qB6KyPmgfUvI
Z0jP+jbGHtJkC4Lg0MfKaQYNrz2MCIoe9/Ymwu0Sqp6GMX+5MvmjX0wA2fmYeLYzfLNAkcNgHrZL
gQ9tl46PZQbAU5yR/W/Q18nq1hVoLzzbhOw37MwMLk8Umo/rp+Cn/wOKsvOKpvyCy56lh7Yw8k/W
wWe+CBQSFNSuZjDY+2tckoW2z6MrKwmBfOJb7uFrVMOlFLoIian1wmCFzxCKYm4J+PlVPd6qN1oY
5NG+n4kYulGP9X6heWo7dDpEDyt4r/w0J4sCT59P/0/rTeOCTSgi/tTOGG6J6T8H+/P4wAOdILSc
CSe6uHiKyXrp0/hXvSi4PJ2df/J7jf288QSjPDPHTNR7XV8AV5pEnFaDrLFfxlxU1+K7TsjzgslG
MeYqv+POSqkMHKUlshAu1yezP/9t3ZuVSyYYhaDZVelDojoGXXKxbc5swSGQYNpJKdVQ0JzIWnH+
rUbf3Te1pS9sO1aHyVzqm0FnquVkL8D5j+kjB3Qt/J1XI17c7HUTZTfE/rjnT0Za2ufSadWg/TFI
s2xZWCcRVG1Tb6ssrNz71dMBA2SIDufc7G9a5PWXVRfySNvgrzLkFpWSawxd4rDeQ83irAU12O0w
Y5AnyaXnu460lSXN0C3sRUh2LPB5RTSfeMK3bQob1V2IvDfQpdNRvUg9tay7a8hmWz+K66TFflNL
wiIIhlo6Gpbn+Dbv7j3tr9GofQ9kxZPmylYmVZJr+3rZ3ZK9eqnnx7+wpCzAC3jx6MXNbkdeznfk
aM1hbLthSmRYuzoEEKb195nSC0vvcedZuMfMcj1Bb9+vf51lBQOqk9UmogeCFPXwtXiEVJ93xeoE
j0/cfT30lSvvHK/g5xLTnVRYgu5F5zrI6Zdg0IDYzwIDRjZoiyqiA5TT9dIdl8RIiLpT7jfa9ssm
tdl1yF4QswmT9QhtYQ+lIDO5shRwXHku/w6l+OqCjz7R/TkittzlwYSUTYah0ob3ZQgBeK9D8rxe
XgHXuHZQiKly3hWU6NVY3eaxM0/pIWL5lcpxxCY6ljTtNgEDHtQPPU5oaKpr8edq+YwRi8vHdSpJ
LHBhv+fOme+2e7gHDkmjlKvuhO3zUGNRy/DUTKU554VdUG8Vb0ifxEAcP+uoYkThMSg8+kfJkhw9
57GjJhsVFUWNU3Und5cAHRZra8oW88eXEFfj2q+p6tl0REYLyXXuTDLY5g0NA8pDvIhxR1gscfze
XBiGGEA5rWDKocaIj56yJiyc/UVjY3SeRX2GlUCSeGctTS2VKAEJWHjqyxKc25HYiASgc4JlnIpf
5syGQfl34YAXYiMkdIfkwU7xA30XwmdpcwHvCwTa+RMreOJsX1USO/IVypDcyuFWbZyUXnonZywU
sKlr7tZJZafYlIMAMAqnlr82PNvwNBBZxWi2IrzkAwg33cDEOV8q9Tv3jB0MIjV1TEeklNl1pEyj
X6YyhMlN4oHr3H0E+D5WlHGaH9CnJhcaOULItDIuEsPgwrGZPEsdPwZkUt1pAu5ooyJqY0ZByW3Q
Cw5p4hX+Pmx+OFj7Zj+HaSeB48p6X3hY44jaQaMLMsTrIKyhLQHqTMB41DAMVAk90fqJbFvdAMtw
qEIyWPf8ewXuj+XB8VpBEyks/0gTvrQFSqCC4OyrI/ACtyOWG6lNV9IlCldb1HAFgqsFtN5I31EX
YrcH3zm9gbbXr2/iru0YpTCkndxt2UDzEh/VuZDEBUeIUDHjUOGLzxoesDj9/ah2x3/4ti38UJAV
yjiIU8g8CcbZcceEP5DZyLllUnYofUvwwkbcrdJihhBdbMQvlf2frk/jcBmaGDg92gq5UU39f9uN
vqWDW0+j5zUGixoxAFLAWLt1lH63/KT3xUy5j3FhKxO3wQxPagL/fpmO1+jvQD/xidt6tGw5r+7R
qS7C6YGJWIkEtrk49S63hm+FetQjNzk2P5nXUkiMampbG/T09RAvcTM6bC62USRQw6ZcR2Lqr7cF
rvoHeS1XnxY/Xi6IXIisyPK+DaRQwm7x8niEKE9tjcFqzSXAIa+b/CHJkHaP6u0Nb0xX73/PT0mf
ndvotyNGADl+kFshb0huhuJ3CPw/J/GPdI6aOGK6IfyRmEn+siUbfZWbqCg5n81YFc2D3WYY2tS6
IE58E5HCHqsl8rCWcbShxOGXWuQU3eHIZzgN8h0J8xjlnZc4UqaMJ1BgPgafqwcbicTvtXn8VMgL
3C3llWPbxkbbeCtxjb4s6oVQUZpQvKdtvgbqF+jiIg2xK9Fdu22Vf72oIRMdDrKr8IYWOg6b6H6C
/m83hKegy1QHLPTz3chzyHnBZ/PVIUJpjQVI8ptpQvXTexZGBa5T14fLNdwPnhT9NedGWxqf+J35
EU39DKEkJtsbPWa86+yDbgPw70aC/65277IItzBIA0fWuPLq4zx2zIE/cbmyv7mbGmPfZesE+OHg
SL8ISwKSEdO+cmV+yDPX6/7bqM2lGan2bt4vHoYbxBp9YRVEvaDGqiMoVMfkKIn1NGoVuwBpRSMY
ZlpGgIhZmSZSnLEgbYVbKPviEhADGmLgv7opCHbV7qoy2gBnCLGJm+BJdELpakeSXccsQeZOC0qQ
6wnuV6yPW54g2GA44te8IhfJ49b+lmAYmDzxy92XNmuy3/EY0nqYxueId9eX5jP/fNU/CJHrhrLC
ikC4IdMqSVSMuKUj8f7u8ZvUtCHhfM1NqMSqgyuK10YtZeTG2ZcwOrQtEGr89nml3idWJvdO2+4a
ugliEYDeoT/a0dm+WazzNicAxpR+UqMxpkIKcPjIk8/P9TWwrAjig7PMO3oPCHJiyxwn3Ol+veu1
KJrfbxL6jc8yDIq1OBYR3Tf8SfwyXGX54o8tOnxSNpDDkHuCOZ2vnvk4WeVrGuSKmkEgOuPaZ8r8
zkr6t87yXGIUmLR8F9pmwBqAsizmk4d6mYRb7EsVfbw0fzq21asSlSkNFGD7nSWtu75tPNDMXhnX
XtROiPpxwEODiYGsRMts5rFnfvnrIsDVc7udlMFT+dA7bfv7UIvS1pAM8Fluqaz8XEssEjGmeHS1
Ut/hnUZvnatU3OYUcNosdISx7sINe/cTN/kSXoccPZMNaK2Av+f9d0kBF4wMujKICA2RMuWKIxYP
VQW8uGlfFIQsHc7SovEZndv2NZoSmKn4MpQ7TP9VCg6jb0hiZmPg33yb40xrGbD2+mHM7EPgnYoz
CfPX0Rd97VmYveMJDrvTGHYgzCLTiq8b456qgiiu2Y+TWuHPQx8+5v+aQSLxldjlnoMe7qr+0dXY
y6wMB4AjCh+TapDuoQrBFXrRTtu7NqPdzUIsEJ/vh0zH2c8a1SNdwQ4nr2ZLCNv4XxeGF8HjtOqb
T5jn2QVwTSfGUHq+I7A3w/dPwpGWbc+cLxPY5Vvv1/PhSKaicb8v7apxg37IwRnxyo93/xB/YW6F
RasgfYHMLBzNnZBHpJ7gH+DUdfQse51N9dKHJBp2aeABIfmF/YygE8nYMj+QEdAGVyXtnCg6tfmD
haXphjq9aRUn/8cZO8FNSRS0HjE5SUIAzrnoj5UePsNbH9OQKvNxRV9QCr2G6AgKQeiLkPsD5ACL
FJNr0J0xhVT9dbVI54triVngmV+nhEZCYw6k6vE94dRUVws4b0Ob9p+uHRLlh45Pn18yLm8e2oTY
KsUxKrE02RhqTxbGgbvcZayo6g221hNYbWdkm9unT2MuvEIVFOP3RxUKw1xiQx4SHA+yuooI1rHE
BRAlAoIh5TIdlzV0AUsJzHBxcEP+jFKFZpIIx2c9sbo1bV5SYC0XxCaWEdyOW6IigUAjL67H7Qkh
MGB8DnQWUrazvYKcTYJyfvte8GMyOhtkKY2oONhY0/PKr0Z6xEwGIkmQ5YuODe6EaqDRccVO1OUK
CSAEn4LwCUl46W4qdDdNrxSYWzAk/LHTlvWz7jRyXS6XehnrXdwmEXqu2zJVLFCAf8qbnbp++fDY
YMCQCLhlV8oZPc88ZzeQIvdj+jsEIAL7kACMdIXzDbD0n4NBBHYZMMhriIqhPnSN8e6dWJFyOeH4
sAMXEBKokDDzIDZfF94mCMrIADNt7eaQzo1wWJoiYw6rpFRT1s3VpcofSFRl5RkTrct3s6G35tZU
Fga/+HUSvByOqtb/Wm5/uHZRsai21A1HpXRBoqWOFv+QFNQ+Sl7ciGaje8d57pnzihCO42kmtW1Z
+qCs+abuDK6ilLTXFmSSfX9A2NfdbLk11FOK+kv43rIOQ5LJuOgUgb1at/BpeJzQNRF/Uuozd07Q
4zuTdo/wiSTE/calPbNuZa67bUScs2/Y6jycsUtmU7NgH/3mwD45u4G2ffCk8zLKX4P/MRSwwrR5
EKozxjkZPhzpg6K0RJHIQM37S1Qr/PGkUdgbmJOW+A3t7cx7tmS35kTtSkFV0Fbwv40fZI56A5gC
4Q1UeTlSO3jkHyVRKTWR/rbO8NSfZxLqVhLCOX/1M5gbonCAKvZ+s29MKcXS5Vm67iIazM0jvu9+
Z4s1gEHUUut2He+5H8YCOjh9Z2GnxB68antERYCCmPK6f4ldjospXIxvf6a+84tzEfGcXXMG1OGP
We5XHdB/W+kBM2tm+mj+8II1DcVnxVsAeodEDN0z29sFjYN8wRSClx1pWN20uvP/5bpTPlkdorMe
vg2OD6qmSQWTtgAXUX5MqVb0/HbJz/E7deTR2Ke0xNL4/6Cf8aVtqJiRzROpajhCzcSvOa7Iekd4
VEmSCXsEtLxu5aMQgv+QgBzElUXenkip2S2/rw+BxUEEWXDbM5MXlBseCCMnjay9E1W16HIp0lco
QdV7qRnBsx7aPdAcgtMb/kST1scai4YtUE8yt0ta7aZCmQuFik0OY1PrH1KE3VkKCPDCWVCxxfy5
9/YuVV7Zx+sS7wBYfdzFnAEwo4isgg3YW90hbKtHZYdmdyM+kVRxURiynUSCFDfugk3HOQlIFTyw
5WEX2Or/HDDBPSJEfro550sKns85dr08bJzC9ID5wxmPeQVMlK7Amn3HsXXlKdTNB4j4sauh54Gu
nJgfzU8u05CtbYLbRLwKbma8UViHy4otRXKcPlXOcs75y2B6A258AmVn6qHST2xDpz5s2j65SBEL
MqM/M/DumBysgnV6A7vsnP6fAaP4urCvcRPTwxnzM7gNFJ5p41CoxPDeLjCTEkqidNZmBViPctVL
IpPpfmCvz6robCsJQxRCcK1x3jS63dDlDpoKKZ8PcXV8yTpWz9oYl3IN6rIJnPF3ZBvhMc8ujbXS
pODZR4Djz4Watpbf4V1IbkeqyLnQgxNXZ0xdbEbsIppiElo/FL7oN5NJpsO0pG9pcFwNz8TbG+O8
Jnpi7nLhz4BnBaAZA/uuB6lUqfbdrlQatcwFYuzozCD5LdVCaj6BbZcPIQe8CwddhhWjCQIsXB6d
d/Z+FqPlOEgomJmUOg5GFAcHkfn4KWypcpmIKICpFve1Y4JUTngkJFliImP2XNCvcvoogic+PKlL
4qfVDjhkT1igqjyyhfxOypAm6/6QMA3XQMlh4BgrZG6ZwQwYjdt7K66v36LXNa5+cMfQVGS+i/3F
B2WpeiQUUG/dZDpavTL75zTPG94jNRZV4Pth6at2NzQYqcoRPvKmKdaXTFcUrpiNGUMB+FBATUpg
nCPalzTG1KbCP0/qwk168HYTSDNHDDWo2hQ5eMqB3C4xl1LGGUOFmicExwhxD6/hyQZUk/Sr3jEm
V5uVrhzXLMheM6CpkQEOHSTjIMCJEvouolLm1KivjrjLmHxybfhInDMEEMkGYe/0pip6FvJccA4m
UGX7y7T6BgHhYbwNmRWY8MNQKrIimSCvcXoTQEwMPH6aeSkmsIt9yNYDfxjp2PGdXRJB8YJ7sFHd
RhyPYoq7zSAFJgod8plP1l1au54oKWWUOOPlslOvII4lgqPBThUQjgwMmon1p8CDb8vUh7o+jORO
oFf00Gwm1lYqi3nSJe5jgYVJww4eJ93IKXNNKBvwkHu+pThTeatxzkF1IzHzgdAuw5XfYxclnTJm
5NE7wofaBPNKSeo6SDm0KtPOZgl8jQ6JDCNhrkUnIxkhDX9kMZq2I9Vxqh8vOBTl/RCWA08OP6l3
mhZqV8TZQpJ0EEeci8vAo+Ca/eKnUGX/o96sxyS0+QJPN00TjicQJoMfRbAQ9OI8CQWx+PkZM3zn
4Me6LKcLJg/m4V3MGB+qm0QoBoRs1g82e7c92VlgpDq1xyH/qge885VlP+avDe6y+c6JIsUVx1Em
dAec0VI8cqCFsEcJjX2mosAqoRYNgdfwnI/3OUvLOYPUz+mYwQKckyvK9x1Hn6SKgs99ud2DCpwh
JraXrDFltItpVIEU71kRNp9XpflILMKQybDbx+F1/wEaVnsZNp2pg9UA0nvI/CHo7+bk2DLWhf0P
qgL755lDwb0599X2ymSi/f+O3XLA3dUwkEz943UpoYt5RDV1237GKfujZ21kyGokGTifTqcNeRum
d3ZMB3lvaQSEnw5g6fg+CjaivKEuexje4xBFdFyNgXXuC2vml6Nmpjtg9bGKhooxuR2e215Zk1wR
9huu1eB6LQ7dHAqCXqgOJGNxbdqXdnkQ05ZJzn2QYDAdEhTiOJfSE/0eyWX+j68ogmwi3Fe4dFff
ILALeBoClylGuH5DdCfO7op/IvNS+y3HZbkPDu0o8x6GcoH45NyGhVoeOr6Iat8IeebrXP3fOmU0
2P1D+RJFV0yH1Y3EbYTC1iX6l3Xqk0Vhhv4ypyzFSAAPLzmf7VgfoCXq/zBHBaFQDa4LL5mrb9SK
vbcG5JDJMxkrr0/sn90CBg0Xejde5HrWNkymOXSubIWR0tIRIEVSaNNOXnBznquER1ahJS2whZcf
9rwBT8Rz654/O+Q5bqGNEAVjOrm85NJ7GuUFHJE2vfr/eUeL28jSGbo3Z00Agp/AqoiFpuzkOVNQ
5r4MiinZOKlwOb0PRytVXQx9gSUjDQSxnUesFMYMfx4LBre7Fhdls1s42x+tFkSgCItPBW8AZP1J
VMtj+hoA7gX9v0k8TLRoHlyWwtBmjUxhzIYxp7eRNSEKLI+MvKMZsNrG3ehtwvmPypGfOGzAxPtg
3QYg7bT9GiuIko4fH3AGopH2Xbb9r6SqZJuo1Qk7IlhvRofyrjFiPpJ8s24qfdpgwpCzcisK/s4K
Q6l933PwEKjSThVL3/eYczi51AdaOTyS4Go61hW/D7yYk/B5DuZEm1PM9DpuVd3tK6AbvJ8VQIRz
EY3Rg20tbB7QXRPLwdovtJWhowba3S1KUvyYGCWhWgqKV3lbaA0bwUbeyDfyTeNsvBdwhQF39t4F
X4+MgRNsQ2Sw7WX6s8yfioUj4irDg5er0wPdR8ULzIvoSHj2ptJVdNTIUmhEy3n4tvNh5kLq0Cvp
TPeEGiCXxB54BDHDi7Wq3ljwAcc89gTv5zZly9kf6V1mHTFBqcZBzq74jskZ6pHYtQ06mupaRZzP
nli2Z31UfAhDg0dJ/mPm33hRZaeNxboSYlGDcsW9TXGG+RhJUnHfqZOWGtbIgGV2pVd5Or2rUwKf
XmwTBcCx7PFrJuPt7JbIw9r4ReBsoGehhtwTQZm+vpvKrwKfPvxS8+umdBnyGm8Dn1YjUwRnUcon
yU7ZiplKT5WIbPWgCQOTNysjM8AGq5zLST6zLeig0/wfvB0dbDUqnHP6iXPec7zhntqQMkMQmRxo
ST1RiQDqOluZsoxiV4kZJ3Hq5vH7Uh7QYTsFchDfnOazDT8oLjIBF0xwENXZ5HRCi2aSO00RVNem
brxFESWS8Bz4EkaWzch5vE5biBc+e7DsYK1hsfNBrTucBVD1XCYHQJKgwa0AhO0sYHHbs6d521EA
Dtz3q04z05w2SimfyqmXmDJA6PR9BK4vt20mFCXFgcwFbg+7j/0iyiJrfSQv5oCVSxFEm3DPFesn
UjkDrSKaXGCqSJPBnOULleqn30Yj58UG8FDkK90fGDigxX2EZg3fTQN1LZaoTBTZt5Wgu5qaIXSq
ksPQ2p1YwJkNjG8lsjYCHqoSfpkdzhsJwlveqvRruR7RQHWk4j7jnML2T4b+mBCOfcO7/abPfE36
95V8qa8sxTByBeJqiOfXwHH7Cz7eWje7kz3sf9kvD10mWEsOM5to7KhcRaIOk2rYWt4cJdVc13d+
0U+fCmrMaU9i8eC9U3Zkjb2rUQCt+hSRAJjzieC5A4pWs63TAqkvL+ERoTPHOc9Nz7kx4sUkoyRU
TwLaw/mdy+hcTZJI3eBZyfFH1cAnK0t8xJ/tZKux95rkaAMK2Bv62aiZf5qcmryeZfHGhElz0n9C
aJwNpWhz8Okc+5ecf4wgv6/gMAZQ4XmMjW2y9Fyr8DufrfZW6ycK7fyPkKE7oB84/yagz+uyE03p
t7PJH8dPYs4vFxZ+MnwX3xYY9wd9bw0sdkn3ED3DxbYKHasvyKyQNGWEaDArwvK9hjOZWp1gkdKF
0CH7d9XDQP1vwIBN6oE1S4Q9FnekR9yOgEYjXZrggTeYYyIOMwffoNCWO40zFjAJycOvkH16SiH6
ZlumVEzI/TppRfojJ7bWs9AuFCc5zPnllugcRcocENwxJ6R6Z0UJ7y6NnLaGQE2DEZpER2zlWu2V
R7EqFX7E1LQjNEc5g6+yXubLL2hESGT0m1gP4dbNFK7xXeCGi20BJfOkalsHRL/H2sMw+jQftyEY
t1QZ8ujjuhRWI9jNk9G88BWo9VhLMx0BlZ94DHjXsfNLLScrMvGWiqAZFW7Ng4C58pvfy2fKyGmb
/QzwxY/uLQBYF13pN/Irb+7t/9QZVUqQwhv/pIELCypkqcW5Z/2pLWpolPqzVCu19FzfCUI6sh1c
DDS7Jdl2noPsX6FpmpmT7ZILg3VTZtTIsXAFtndo0doZ0DgVP0Y1i8fvf0TcTH96IiYMwYSgb+ew
YCjbr1LNJGTn0OK8ifYJJoB6w98t5bc1vOAff5MwGffskRewXYvwauNyaGPAddo7ifylzH11qCB9
9FF+MSdm+GLNx83B19hPYdvzEl4R4r+CDJ6gBGpeNETxzkFS9sO/VUxrv9FWlC1v/SeIoLj9PYW6
xygcfHXJz14uHPWaaoo4qwtJRhfsKRk74V3G838JTsPyHV9/wX1lIJ/KoiXeBpZ8+yB5+/X8LZi3
PGQ1WMkktPoHQc1fKUUDXb/moAz0AsVd6j2eSZaLzYUJKtory555nyWDqGgamVYt7Ho0v/C2U2dB
f+6+o+i9QXbdyJ5YuC0RHhr/XeQges9v6u7KJ9DLoPdkxC48llZXLJV8pNPIOWB/Qav8fqdo8ykz
ceOFbI0nXP/onL5Bfma132ao2VXnNdssECfBLj3yN4UZU9ibic3JYXLBzh/GvNcxZdq3BLrpcf0e
jm0t3M3nAwN4Na/QBEMH/0oNe0ZgsfiWYFjVUIjQICj79jK43zbdroM/9vUXcc63dW/7nu8nM1YA
YixrjMyqcaJtMwCjrpS1ZPeXJDImtd5G43vrYMw5w0zq8hzu9pC1lZh1a/gpsMYPQaGbVQIWG7Bi
0pHW1X1W6VIVGaQfW+CfAEO0tFOvvdtvyKeuVr3AQp7LRU77W/KIFnay3+ZrzcNEqmGUvdIPQz96
cxEJyRfpFltYw3rLv68ObOQQcFfa5hT586JKQxM1MDojfEf8ASdBcahcqHEIj4foKIEZ+zSEEZSd
EKG4ZisSU89bEHUrTBBkFgfOO2wSzfZkhpHaAtCB0PhAYmHVw4agtZYKVs8F7S8AcfDSALjC/HP+
9Wyz8MIZjEkWN6liRM/mKySMODlmEB5x/T0uAoGT9QXOWGM/hKx6OFMEUIxZFxuYvMQ4Ta5+EOT0
q495QzxrIBbkDfqCBFb/+8tyx+gdbOeCnPcJm4gUXwC4vaZDHPImVpUD1PO5ceRdlSkU/YtoJm6I
R2UjRcXYz4zrwavPkhDDASAf4XTgvSR0FJiAq4X1dyTIB1B1NqNRSueEsjN9d9wKDhHrsQ7l2Yav
nM29z2yH8DGBbhgD6dCZq8owvRYW2FvfsG+SxAzAFFWKxdu9NuCGtqXwQVzEnYK57aBi+MNDqCKV
FknrCj3oly0t7/QyNtpPcZI8oPMvu+NW80WcWkbwxPBzNInbS7yM2lxxoE+00TsCqcHKSWXMRadI
k7xEqmY3fZtr2Ny4IzJDQtzhxZuDJFGJxbRcMlQJUxg85+VVp1pjuj10zGmGsS0GLSE7mwY3oMOm
gbZTtpV1rxPZ71qtEZtqVi0nbeaB3NqmEq2Q7NH9nu9dxwVVS5D3FZytVM9j892iUNs8SKAdtoPl
hV9NPerC/enEEKWmUJFIkbJ9BYf9+T7au88nBlJA8a2c10juDepo8qsF0lN607JJcRTYA91OtwUw
Ig/O5IfK2bHqk3elIiTRT9dxG3ZNUBu6FS2c01B3y4Dfw2ofMVQe/luqyOmHMT3PoyQxVusFD5n1
PAC6GUotj1RG+O+GqazDF3JY6v9H8Wj9ztab2FkQDHCZxYYQ0FRStlFsljX9i+lU89wRT3PNi6iq
aF5lU2LVE3PoVPElnJvqIa+kIIoNr83PoBz+C7wwiTenqWcHUVzomNxmwt083jquTKECnw+lArdz
0O6aJzQH+kfUx3zaHIbLAuubdoSw9Aj3PnzzFxUMrS1Bm5/jqCVxl92htOLQ18jUo4nIrN0GYhn5
tI+h8WT7T2dDShV9X7f8voB7Z3DQIQqfS1WElaIWg6Zb66zBEwg775MIW6zdm8I5QzMDqH4aF5hm
ZBGn6MX/fwZ5FJuxh4psZRtHAywB4+txph6K6b2m2DsB1PVvyPbkMrKpio+kIvaDfiYp6Iagdjv6
9v//lH4T1wvLPbMPUV2wsIju1bbInLHjO7hlBuxED1yMzbXbI3GhDBVJL5rBtWP9ZRwDlC+5PvfA
2WQxlUHZLzzR0OaIByb63x9qOQFsJLNgnJYMhrQxHXlxaDi2qUb5ldvm9hLBmUK9k2dLigUNlPzw
3t2fGpaETGNd+poTUAuVjLv0ZxaZ06EGx+8GK9CWO20JWA0CvTNZO/7e85/i8zNvQOSi6+yQCHOA
I3HxCLoOQtbssv838qfQqSTAxmD03LNqWzuDRMqWjbbj15+OpGVw9KdMFswn4mgBh9sMNeFhjkxR
/zXPwJri2QYjJtlaYBtlzq+00dIU9RWXkutr7js4kWN5M3D5L4jlYkPjjti9lLUpYKItIeek7JMa
YI5DSTp0SKgzaTEftezE+r+UQMnnnHyXf2fkPOnagE7dpc8b8U38rWdM8eLHHpEx/SEf0hvX8+NR
pb1YYLcvnOWCq5QCD+v9KjmrtV9Xnq62XTBV1qNtEN43Nw7f1KAZYYg+da3grme5h3ORsbl6W7Vx
pY3Qw7cBaiUrVd1WHwM0juC8wHya/aQI4Ppq2gKt6Jrguo/fQVAccJ8h51LdU0oopAXO5N3Q4j07
xdLsL8n1vdCKI4sMEbL+AAFOOclhgJi2QLlXM8OE+X97cRKStUGIe5lMjAlCfiN4htsCYkv0TqAj
qvJYvFAZGrfcgYGCEMl2Z8+XEgn1B4QEWkgSn2uVItN8G93B560ZheZOEg2h+MYIcm1jGmnpDdua
AWEYITVb7ktyGZlsbSgCDsckaWI17XT8UCO5NvPGJiyFar9HvTiJHoZPsNNuVc8j5B0brzUsfryN
5iQZk5Z61E8R8Zfb24JsXyf0bszCsMAY6Gx+kDhf2gcAumQ47j08KqRqVPOxWDPUkzFGt+bKmIct
LTVv7yuh4sP8SaIzgRBLUFNvi05aV9xhWMWD+Pw/Pm/Cdd7UqKLmq8SKahnD+AOR1QVGBfdJLHRQ
Kav60iyTDA1HrMwrfVbk1e19Q4wvOKH3qDPVqcE9CJ1TWUwD7V8Xr/3b7vGXkf261YfUAMhvww9e
7tjs9b6cr/PDJYVzqlu7XClBsgNPbOKzcn/yRAypgwQ8HARUxxMD38jnNSJ/luvr1ihQ4MEdBwFY
b4rsOzeOI9Nur47pIef/0kLKMHGmKktb28x+3a1mvls9TdH5ZYkY3ugCbNqE53rwNU7eQJG+mmUK
jY4IIGCVvIoUy3hV+pf1JK5MTcX+UXR1M5uFNmKZGy107HEgCaM6Gt3YvnBuQxLsC/AsSKCef3QM
KDsThpFGgVVvvSsEWHCBrldEUhLtJaF0ecsGTzgSqjzJitFwkz/CLFLtzFkGw5RyrgejLK8mG+bA
F78Mg84ZBvyLy4BL2VtDuhuTKnqLfkbUoj6taZVKVEX3d+d3GnX7Hn5RHJulxI/npBQVm2dgRXRi
WhY/zYk37d50ctNdp9jP2GKgivU50F5QX1yEulOvDPxNpqROzvHaG9Zd0JA+5KGVInbhbWpBxNSo
+WiCFJRBjEE2lfX2jxdGgklXIHJYnuQUUjWjXF5ET4qNWO/BlGloXqkfObgClDoJ/+ciQvrYEqI/
PO9WkHWzlxzeUobIOmiKcTfo9/JAR1HDIN/QuUR3GAUxUcXjtpscoJp/MPSNS6/Ec2Ipw0iPPoLS
pQj+gelcl6yttGEueAV0O/+ypAuvxdox1DtquyF/0osp7fVlUjN6UhnxhQLk8YYcTtYHlj5pM1wx
C/4NT+AxE92AZCJeLuFT0GvtROcg/DYS6yp1Xyge0/5ol5mqUAlsSsf77xrESNt6i5wKCrxU9SFE
0/tJlCGAMrrHxX03MDDXVVuaJmXz40uizuZ0oYy810qKM57dGYXwHK3RTNWUg3jrh+xJw4chEl8S
vFFJ8HZb+1Ro7g9y3VpLln9aCaRYwP+Dthe7tUDOWA3MfmiHJ8Sd5VPGlXRM97Kfib5mtPAaW/gO
kOWV5zlD9yfhdkFYJes8OfDc4za+UGn7MrwnjsZ9tVSVohuylXgeOhEiNWFKTa9OZNr7kV8MLQFw
TR6ilfxej9wSZyBNeJMessBghYUGmUaR48FzYjmykx6exM75GNRcrN6+mfFSgyA9jDepRzKRNMAD
2tXpF9uEO3CA2AMqYD2RjUAC2ztGKRlS+RNPNGvkuO3L/IhVgtu3Ca0cTKxfKoHg2f39IovUoqgE
hYwdscGs+dVPoHKLMp61t84SO8P4et+H+iTN49FEsSC0d42mctTxx55BZyfxk6MTd4pDnTkE5+QW
O60vUNj06AEdTp6oBgEhDKBoY1VD76HYzx43mhXdUkVdvyQddSgxLFbjxRjDD9zoJjtZkZl/EQ6s
C7YnUS6G7F2cF26Dw/Bs3X0V2vO8oPuSvbI2Y9jpJOjC2jUfqXL2+PMFGYavGSrRqI2hz/Md9hDk
3oZvd0DfL7uz4gjjwGVy5M8EMaMPUuZeeySqewbxCl0Z5LE6zWOc1LPIiRYhFaoTtjEh3NQeAks2
w8rQq+cjZ+/VARnX7qPzDPK57j0z7vVU1zKYXLuzM4m7CQ4H9PoM4DU+SuBfnQfLkupRwRhQM5sy
z3ECvpF9vJ+ijqTwL4je2DySa+2bYTpb9djPAc+3KnK0PYM0GzKYce2UOXjSRjasEegLi2bBNoz4
O0CfunU2DKx9K3Q+ueManQn3ZROOBsXj4b6NFg68WPRvDeQLGF6bgzhfX8HSBy/ZgHekGadLJm/4
z9j/05WdcamAc+jsb96jqHei1hwNj0HmtlftyxcHCZK7/WXqD9Kb94n4pS4YOhE+aNf19BiXMU7n
7HO2wVDmNELhaPqGGLEfpiz85+a77eQseuF2ZtC2WzurAe3Yet0+xPnJSebYttlRO8S+8d2tlmQ1
hbuBGads4CbWeC6hJmR8yIJeutysqvT0ND61a5W5Eo/YmVtwdQCInJWmFLQs2+JQSdsN4XpWnlt2
GT5lURhSvXaG0ypeOYVVjLJ+MnoofAP9ELiNGJ7NmN2VtP8fIhTFJw9I61uWiWYsUTeyVP1C9/3D
01JNZhjsrwqZFaAUpIt97ID4jtwiWCIf3l4SOWjwO3zbl0QZRLAsHLwX4C9vUOqTdxxXnnrAQtcJ
G9mhnEuzL8bW7JQQ8i8jNwRsyjOhsfdBCMkUhmLvNn0azb99yLzlOJCBg6AHt7PguHG65VeGwqIy
c4ZXvaXgvA6qhTL52SMsC07Auq0/6Ynw2FYN9kltqcjQUkulKnkv+OiG8wXR9wkMRM5pnYW00fc+
bLC4dQKJ+qFeqldKxl6qqpnImfR9yWBSJg4iLE5ezJBibjh96NQPwq7ujRETCO45K4G+EgqQG+OV
Uzz4ZOStGaElg+z35wJDpEGj7d4OhMf/xOjSBieuPFJ0BIv4Fbu72ek3rSHHr8cIuEXZil6sR1bY
xy/z/8S+c/+sL8/UlBQiO5QzsrpdcWrSVgLxsx0pLZ9zYhrde8GGKPo7+roiIPTnRyzeC9EFrywE
vrGGqAOayGDFGnRJDtxJozgXwZE0US+ThQDGAGgt/DDNFDQVvGeaXCGTTg6BxbxH4jptuAbSV0/Q
duAZQxnHDSOXmVIDwVJhkEkhO/64AjWLpa/MY1QsclL49J/eIUWvn3YFbo3pMu2gIaQdo+qbOkj/
64P8/Y94QsosQqr56lpzNLEE1CqSN2YkTt9d86t8fFKgQK2ZXK5QSPomJwx59iBQFxBtAAf06Aw5
fER6f3jYfa1DQ9347QInmy8oG+Z36WZYeMN2rT6OU256d0rJJT95Xd1mm+lVjvyB8Xuhfc3cd+6W
5x4pJWuL8JUEWcxVip9LilBb5Q7ZNGotxA/Z1laK+as7SCvM87+rbYsYmr8lgpwPX+wlVm6sQVTm
9B3K3r1m7DIedyjOI7qU0AE78qTpjZC5ndR+GhCNShrBLDjUSTW60qGlrQslV/fpYSWVPyP+rngz
d5zIIIhDrjeqvyejJ1+uDQynMH7FBXCNO5BnbQgRaXvKXw4/wZU5ot8tX5E3YlQPsIF7u/ZSRlsR
OK0Rh70qVfg8UYheA9EgNhPTEnI0Iq9k43qshTo614GTBHOQfPrfrmkaX0kx9PHwCh/GwoxRuxz0
TvzqoD/Ua3DDaS3ukiutyO7eu1DDdtuNgwPb5KAx6Og+YkdGABQ/IKYdg3YodJ4//0VOb+rc4QrG
JaggNS/FdQziXwIOgZTog0ety8dskdbYooxiuLS5HV+Ie+fXWBf4Fz6hggPsNeyKcJHCiCfVXSef
EiGR4lhhhZZ9emWWHgn8JYc/hek/yaCW/eTOTwveS2VtPNEgzLU1+JmEZ4KoGdGerB2MlUZi5jsW
H6q9Dw3UqH+pD4sB9RKihQveL/wHGPQSOQnV7p/mutGS6pYqKjjhqBH6UW5h87OFvAWS1qk5frQb
naJG7j1IU6+Sw6k1l86QSO1QMBua87/GApTxzmRDye2XR48eV/h/CV2kSwLNMPWHk3XvQoiFj8HJ
Aweqazwf1ONo8AtSTq8ckUCaJx3kwjWqgV60Rtmakxeb1WqsWZ1Zcu7VA/CENiPAWS6dzrymJHzr
dobcEmS+R9JxlDo/ffQ04fzR7UvA+a+tMA+imwwVGC65iVii+mjBBpOnPctXMYUWrFmIjPhv2WwU
QES9xm2nGoLAuTzc9PVsFXIsU1R23h/xoAhi7t8JbvSOIy1T8Z3C7XLdoNC9Va+45A2XXeLsikDT
bQBgXne4BxKnPZBdnZ/7AbiYsWf3AqFsBZr9bHVxv1aQXso1b/sDgf4ohG0zf53Wa87APsrCdGNq
1SLSdooNp2CggFudGILPh9CDRIgf+W0wBt63H3xR81zlEUL9ivfgWicKsEtKPKVnTy3/QdpwAiq/
/1VNAaZinfSUxck3PFwUUmAPsPmcRtTKS2h8GI0Dt/Ono7DczgrssU11LY8nuPHfXo8D+xoSrXea
qlvFlE49IuD2P/Em1+RyXiKGRhbos87wBam55jIXYUZRHvVhHrYDdDh2AopbcWwp9PNaVC2cFHns
HFRRTZOTDaPF1hYXViGLulPgUSl+FjyAS4U4WspzDJoBEIKDAaDy95DkdPjYwpfHF5wEi5bJm+M1
sPMCo84H8i9LtaE5TqoE2bH1Zq5nkwbWJWugkc7XfHJKsDT+sh/+fId/dWPa9jI9vt7ofSMQJyiP
qB8y7vOBYJOk/YujHBn8yzL5tzYNplXOo9pNX21GoM6iAxbbkhO9nEhXmRScT1ueQquqZSjASZTV
dxXaLYWDNS04u3uBdjQNccRCJJ+TdPbpaX6RISeBEU56KjO/sHptr16H5tPKpA63oETrYp9QMhxZ
D3ZHKLwm/a/vN58iZGXCdm1CS8QjZOcdjKa0m6c1Pfb4DJcU6jn3aIrHibUfwqeIdMrD8fLZm/0u
ReRrQtP0KA8VOcX3q5FA0hCRIAdeWkylo2C+N6zR+BgLEXNqlSMMM2Ft0qCccxcxv1UgbB/g3+oR
ZiluF9p4xbQsZTdcshB90A4Eun4O2SaIGE1od8wq0PogJigO9YmEZT3rxH5BZdMQwt5MJ6/DE9dV
o/i2X+2IPXVU5gWIGj7NwHp7ItASXxqQXuwd147KmSMBPITfFiHR4viLhJM37Z6DY2jL/WqqEJKV
1d3vv2D2oL7mA6dbbk2L2f5kzMobwu7ZSyiZLNpFxXMLpWZNRuTpgYbz2Dy0pnKveGzHJ3o/fFQX
eFhaLcx9tWEpTGdDiPcaTVKRloqT+iGCOoPSUmM4LXwBZ2zJIXA9Yp36nW2HsNzHrfW9m7vh+fu/
M+4iJUazRmTOJt+IF9ZzHK1zbGLSja4g8VyxKno/OGCAYtyl8uIaYRrQmpUTWV48Yw21u4dDrA1x
Arlxq+b2dCewcblvPlZ+XMU+sCH3ZSPtPU8MeEdF777NcCgmwwXYzJ0fAYytOdALmwZEbcmCfSad
DiYzzIEasFFDmUT2GtBya8FicJwwKqMRp1xSVgpi0bxddvRLdxxiBluognk9JJi9TWveW5E9LS9N
OaPzZWe6/nv5KMuQPb3GdoQOxi5K1waYrpR4dwbrehgHWO6J/j5U5doSW6xLVeZZWZOScdiGcOX6
Xze/v3u7s47xwDOCHE6LquuBjEVGUGhbMqpi3vSpRk+xqqRH2qYBfvlaY8Hmhiz5k/Gq/bluqi8y
tVaMVxVLJp96TAy2ujPD15OMZJdlpFKoeTfkBPDKfVyPC2Bc/IxJg6mjRssWW76h7ef5LU4byWxs
RqgDS1heE1MHs+Q3PGw0cmccuojw+nQ1ztkDQO5Av/3oy/HV+vmrnTKd9z2Whz/VGW19alfKNbHj
uWpvFowUCM5znuNMaGB9h3GrP+s/DKSLg94KJ+WNylJse8fUeVk1jNMC+zzngBNTw8qKSMDzlXLu
H4dnSE48QAdktFPFK/ag1D4MRoH4K06KIg0zL+2S14zIAlFJbTCNhWXsLQQlmR88O8fQ1/N3QvFf
oJbvjlGOmTekjo2vE84Ayv7vgd+Gl4b1wvhM8nVvrpkFA0qLu6M0DsiA/XrKzkhl9bR8yQlC5Xov
iCoOPdEQzC4IyMTjLAzGPPjdvri7oR44gFMMTMB3VnfqUebiP5o6OR8w5M5b2Mbpka5ZQiGyaBuq
wY9sPsYRCY74Vi886fSTpCAguHKhBwZcHjqvFOp+GRXvLwdPaYna8VT4Lv8qs2Ef0QhY5yOcN4nM
/TfN+xApQkeL9djR9pVl2tw3R1EbxNZrcA8T3kah6oJdxboy7TtxT20gd7v3UNzzl4Bp5O9iWtEm
xt0i5V6PuUQDP2kuYzOmyKf81APK8+SxXU/ChzsQ9S8IJ0wqtxIrv+LmO8XbzGci4FJVRoqEy2Wj
LLa3n8ekgJZJvEv6PNo4klwGH3uyDHc+a3RvUzpA/gZPvYnV8eKt342D7xw/BsrOHlW6+ryDZRIf
F4NG+Ty6bjCkFkKCvu6QdeaYY0oc36VxRqe/F3T8uV864GBxk9uxgd1svNHr5YcL6I6Ki70PQOY3
d6V9ZFon8/ClUcK9pxilCp50sT/QNswd8yfYorRWPMXnKS9vjCkxmjosdDdwJgoV6x639wFIsb1k
BPT4eq6iDcMQeNT14T11Iwm+BXZMSxrVZgcDoIbq7jmArCBaRGgHOJYSdrTMif2MIJwUNY6BZm7b
XWUMLa/Dos/R93muS2TMkg3pZ2m85C/4GsHltV1xiYVGsZHqPQdCDUQ00Q39VUusOf4gt88eiKwN
lsTGXhz08sk+DSwQduULXAOzsbF5+/BiLwdmhxjOxTofX/M/YAzZf1istzXyCpGb1tRSFiIfnIZS
m06TYRznbiGd62hjQN7PtJohG8P1F2KrKR5CqoOCmFI22sOyGuSx9iMd5y1HIWl4GkUFISzs/rxA
0uOrQ/AHLkZP8tLZoz5IpZKI70benBl+jA5XWy2eVFzYt3ERR3TWwcHu0qP3XeS0l08uUkAWNyPg
z+tSBWUDMxQhFprfZN1BzVGwKqdOH2KGnIDAReAu8jkbAw6D7zqFCIy9d9LN1bn3ZJatpCJOXjPE
WgrWaATDcTMgdVK3dtBNkvEjyTgK8noyY1e4r3mUkiCZp4vvO259rPA4J1sb4+o6PxDcuUbvFCdP
M5ubRasT4AhONFh2lgl2y5cNzJegh9rxS+gu6NTSX83/pVKFpmNs0GpLCDlG+hiPJDSTfONXUG9e
vPTbiX4u4gtIiGjn/LFVjfd770MozBxB6MCa6tFA5WM5Ype+lnOSSqEsp+fMEoerjnZ/7poB5koJ
tctHJnWR8ju2W326TNuEi+QHK2ImTDgWK+U/o6G1arBQjHy7XA1bFyczx6tlnfXF0JRjh1v6hC2s
6xta9f5gdmHs5eEhG0QV7sbOOva8LTFr/Vlnlts6F0WuF7/Fo2ZUUx80SgJMIwFzbfSBHznNJsDM
pB1fRiBTCiKeKosEGKrwz9Z1ewuiXtuw0GzUsNP5VV26+JzpMAYsj1OdHWTKY/vxO+RRj4FAZg/f
+NE5SzboWVMVTHV6UIPrHL91yM6LP93Wou7QZez5wS8HEQowiXRiFTTG/5MUC/vtZ4qzywXeinwf
HKgA32OEIssqTMXa67f+aDj4jsVyWZJKtCByiiuL2aBwGD/2NO/RnKO14azLr2zTXcW8sb0GMQEY
tacireLZzs0E/cbpT9o3O/cyQwVRbpJoLtai+NUCuGgbv95dSRUiseAPdIelXoxy626o1VM4v0K/
8AncOkhgWW/6KJ/j6OE3PPplky0j5uQnyS1qUTkuYFZQRPibWgk6ERDLHXjbereZDSnIe7dR8Chl
c3Vkmr4UXvRHmDVybvS4B3BbrJcy9fIr9FbTH1tlqJNNJc4p501VzT0yPvpK6mT4TU8XjYYOj5R/
6U8KhrtxXE5nxrjZZTh79/EXEkXdcyXHKUwwFFO1h4Yo3GqAInhSvOSTRFuXXp3ycaCXVTFyRWXZ
I4u2xoO7ReDPS3Da97c93Uq7sPQp5DSrnpw31KJfJ+qCGcxo42Z0xiybFJUtrujiHGNh89zk/ZOH
vNwQ266YHBXIW4V+3+148r0HGl/LC/lhkzsZ9s2UF6EvN1Ujcngx7mRFjjvfUFd8V5H6VDeDKNfZ
Fe1ykW3qWyz0MmFqMDAMdLnTvIaun6ZZzkYVljO0Z1mVfWkkdMS2ylOxbk8d7eIzS8IFrzaB2ExU
SXh8ngun1HRf3lA14GagctBdsV+Y5YM0WBAosU4N8QYqzymaIVC0qfKsBW+IMrrkbFDq/kbDZS0N
5T7NHIiQdtKshtmCJWMEBJVhZ1XrSSNYREWxkGvQwNtIaUgn32e8/CO/F0tvjmKQvJ1j+f7hert0
bkl9ZnUnyUky8flCpUe8FAAhe54D8WCiKPUam+u/1C2XCL8dZHSYrIWiesyH5P4eaoi0n/99g7/a
U0IzXnZNqZ+uJePkyee7hqpszQeSY6OlN/zx2lK3X2nqUapeEOW/ZxZNTMDhCDMVnBqa8/r6XX46
TPqujxoYYOudXjJHA7/aU6mDmVVHNz0KqglkWKLI7W8oS7SpCaGHlQ7AyvFSRoFxTfHdiC7QdX4P
n6RGmAC8j3YboA+twAdFToFrbjBtUMd+pgGp/wudFnRdci3Dt0LYv8/2JWgj5ujVqRyp98kdWsRy
9LB27o0M+cuHQEo6FvMutHN4PL0l+GHAZq4TAOV4L6MGaAydGvDouBQYBoEe5PKElhtq8CDAuvrw
Ahbvbl3Vbm6b6XM8QRrbsM1/9Tb/+IvKaKCvMqxKwl/eFT50I/jccfQX7fbrN87aGBJbAbuAtQtU
gys9MXKB/p5ty+ge94uMbnvF77twBYTKIDI70uMWFqdeN7IFJGRWbdFLtRkfw4a6QcraJCXdyWvb
rEPP6PJuAcsBT6wKph6XrHhWhW1r42kj+LpQNuI6TOaTLarj9RURBbD7eXYKI+cFC45rYX/acfdp
c02A66BO/LP+jPuAhsDKWqay2b5ZvnlCwx3Xu71oM5vDTp5ZzbyhthnmKl7M63/GoyoTnDFaiL2C
DMXUh/XZ7WLqWvQGkKUXVpfrfq2KAgaqSKhcMMe5l4fbnX3ox3xBcHodAea7pNBIXWYjcaCgMryD
2Q6TWKYoLc9E6UkPmeFh/euUsMou0DO5sO7tHVvn3VnHKEzo/sKDi46p6Q4IBVmGLpLChCa29NEo
iI2E2v8JQTbWOzQk3NM8siQ3QpgTtGFxFsh1J45tuJR9qOb9DcHF6No7XF8GeCZnhlvF3r1X6kqE
wppq67szXXt2vduK3k/kjcM4h9KGqK3aVMSz7whFDm3QDU8+eypH3EDuVCAx5i56xARUVvUgJEw8
nBcBge5HdUcepQaEO43Pw6tmmQQu2EktupngVo8LHoQsT3VV7XO/Jx6d8/tBI5VRnWWmeAqbNBl0
hFNHp81YOKsJxdnWnPZtqN2K1AdHG7s7IWtkbqXT0zqtg7aewdPeku6iz19m4F+p3RYTwIwCWupu
KkkQMNEGBLgJ6ONYXSHUVv1qLrkP7SeRDjhD9JOdWpRMbvp+2RbFmr/3jndXu9kHUoOtDnm+JlpL
h4eUdH5LOr8yb8yYLT2E5oe7gpmeaTZRgHMDfCiKAoyUnvZsdWfFbXB7eNbIY/y+G9ND9qwxwAHY
suHBvLbaYPXLsvPDUhd94tjyKyUWYtbHWTtcyntt35bQZynFUI2Ukr1XtoWxF+/hCn/PQ0g8npNJ
nInhBq32ZSmqnKnS2CtFQazdvGX6Xxo1aV4ogBZ0JrbupeQmdgLOMibgzFVl1s0MJ93TyavF2QuH
Y+RNwCLgx0m+Up74NYDP4ExW4wOGQr3bAJqCYWuS6blMeckF0gSlJnOiLmzsPUQlQC++oNqzsE8O
vbzRgarSfP1bK8vMTMv5jgW7ROv0J2GNvWBxalV79zmaBrAJpu7aBv6JAFqCXm1G6ChK9HZZFRKt
/ciMWCMBtwZLEY24OWCkA8+hRED6GXM4wAldqf7I3C/QANDc01uO2PbsoW0mE69nb44pFyST2YHr
qplTl7FLPkS1Fchyd0AopAQcHRucuexW6FvXX30zko3fvRnsLxwgK+dj82MMep+e7OHvFl7GWh2z
YqqK7v7+DNdITj8vyivGOlIPN6OoU2tfoJhDmaNePiJfBsAaQorCvSOvm11vT7dBQJIrD/cg5dRu
M4ZBHQqBMs4qtTPqW2PDR9ewJBhY5Ru/ftbb155YLDaCNEindDaJlyQebT4fvNHHpkcRSyA0Zqc/
9Ia8wWI+HqNm+hGcfXub4xq64T4Lgwlhv089/62PN7W0LI8xKaDd/0pJ6YENgi4qCpBQlvfYg/ym
/3A3JqFA2iPX5RC+2oqPcx84eFibUw5JZ8lyNW5B7jK87iJ1t3QsIgbEVYl7AONQh5IKkiVFmK1c
u/joSxEbeg9UuSxu+CJ9XzDfnvwngcEXDiwgN52e6Cuc+Wpx9X4/MszqodQiU8T2ffwee+vkeHp1
UMGr0SrNDvF8Fr5Q8rDBH0/wqlaozRLay1rsiOMBke+bwSrDgo9M1T87j1UkmyzN3W1hY0SF4RAE
fcrW+sXD8bvJGM16WnC/3DZibFIDzvgz/dyhlW519LgRkkGUS++7gcm7/91OkzxIzGL2tIi3DHUB
mg5XFucqqeIlx2k0FTFnHu3wQrHYjoAMjFQOhcMrKoM2qHWLWfGOQG5WM4O0CZy2tY9sj/KhIuCa
VCWG6U2rPdXQqsBiWzRTErqfQVee/wJDmWoprOoIGwE6hvWhmjSIuCOiCHzkc8tXvFvwZkjXnKHV
nAC31SrK1m1KNfbSAan7VC5LjaeZsJEiTCwoASf+gOYTZQ/Pz2y6IA8unlTiKXcgPhvFTom49/qf
dJUsGPS86zL5Bcx1lqHrGIL+m3DTMj8HxSFm70DozVXxePps9HEEyOozSj01r95b94d0k3g/gIws
BgsP5066i911hn5EjZi03c35N2vDCL+D+lmqenBtMK3ky7e5oAvgrhv5j5x2QfeOXE91FWXWCAVD
oJH/KSi9KhhHG2Viy7rUX2aBhEbJUK+MNSAZzsvCE/2TzrJ6zokioYbvlpgWevvoKlup4qIMZt3h
fbNSQb1MpTmvftQwknuZEgXZXlUAuSpD66H96ru+j6xmehGF60kJxD72fOVm3DiDJzCmdsKsjXRg
KPfDMVZ1YtPUivCs3F4Hv5XnpRypKFtqqVE5/GvEKkdc+sRcKgNy8trK43HpK1TGENY/W7vXaigB
dw032aXfTT9RSx/pyUFOAZ7hrd1H3HBpqQO0bwh2HZbnkzm9w7pSLQPXMToE9k4/XIrmKzte+Z63
lQpSYoovz/mW3ApJ8dTe6scZE3h7MQdclfF9eKaG2wOKkN5tdR7jc3alHAdsuLTcgEXQOuVTdZE/
L6vuti0vs0WOcVOmNGkXMBQnJ+5HAFvBbBog07UgF+NaJT6AVLu3l5YRgVpY/S11JwZVRpYHuESO
i4MWGPwUxqym9Sn1q7r1ZG3oTGNnKkvxUsf8R7vLnBhheCeaS3HQEkjYI6yv/cDJX8IGrz0UDD7k
/5UFlT+sAe397mh9Vt4RGZYeEesbWqQQaip5H7KAiiU7Upc0EVAYUPcikuWLCQhOWfatAY1uA3UO
pdzwmQEUnLw8dAdAHs0CqiUIUuJqmtvEd0nKfRav5tdLANX8PeQdZvNB1KdIxBa/K0lSb828kJ9P
pHPEL2sEaDgu638ac7adBUWJEjkWpuN3utPuooZYbgaP6vPMlsg5fuX0VxyNN9TvOcH9uJgRRGy+
yrGE6CPL+HqZAnySS+2qC6/Sz9WDQhCnDBdKr5lPD0b853EutRurFfzayUAmVeRzQHGa9UGEnWko
Dprco/jllkh0Bh143YRONpDeLgVm5SXZOOIJQXHBzUmPbA5PV7G2dpm/WwXRBa/ZGoSin/SuAGKM
oeO7W5twbDvbD9MhHUl4ssckFt4DvivHpCqc2cz66ZOvVhYzp5e9fjT1j7pl1/HTikyHZyMODQcG
BK8hRDVlpsKb6rMc7M0yDR5kjB3/ubJ30r6ZHii4wpp+NslxOjx2yBoCR4v4tDCZUmWf9TLFQyjq
hg21zqyZOAbHf2UGjp+OtKpA75pnla7wEZv22EMeOgbGP7ORI/u+5XG8csU6Kf7yd3jgaPwmbzwm
QktH6omzbXEW04CtQxYWoWcI6050esaKY04/fMIVdy00vH55q20udRKcfwLAsu0kb0jNsK/cc6gj
3zKbfJzjjYEo80uEzNMG7phIS1D3qltqsq4twmP0h8XxDEMBPKmsnqO4pye3IxQ/j+pPcpI/YwXY
NzIh11Gaf07aK6L2AjpQ91MrXzaZUArDqgfWYJwV9zHE9WstFh94Fnq7GFXR3CGfGNKpYQwQrgaY
sx050oEtRdsJzpUADPDK9/D/pVrls6ZBXwX5tsTujot9VQSrMCS8PmDsK1BDXXMQpMCR+qWdXEWP
cXgtWf/mWkqEmwDDCvthihVD51quMzIgoWQovmx1QN9CzP2nw2gUwREY/WlxYlq4MR8tltnz1czq
l6xVbB6/M02OqXrJ4k4eFCDMIwJ8AQPHNdq1wMKRh/wWA7Emz3J9EdrfHlcVEng5LasUSPbpFDV6
ygdmW8loOBUlg+25+K43skyVlXCW/vEzqqnNIVFtj0/YV1LVDp2axMCHSNsOBM1A0v7UD0PWWHZf
Gxp8pEFMSxg7lQi47/yF8OTQw6mLrse4FJI5jaNgmvBK7kR3nR86vQk8VWSrO+VFtheCKRLkgGyZ
tfbKtXfhxDDVCL3shqli+ulRqb02NdAIuq4z7SpPXASPGUqebITD5U8VwHX7getreMpAOOpG3E1z
qiifmOYaMSY0ZxG9GiqGJT9pSy5cZgzKQVDGiH1p9zjrfZnNjX38DwRy33BhIWK+DSf+K29vuXBS
mARM/k5SmQZhPgl05p4evYPDuk3B3vRyhbvotflAHtK50lMXjEUwMwIr6vStu6WiAQE5L9bReE8Z
HmYuTLpPsho6yxAymvufR9YaXaMRsZAWA312SDnTCtghmDhN3U7yiD1m8BCQtyjON+oYGDbJOdlq
/Bto6Hw5DjAioCS24VcoYaEsI/3kffCPCXzBjJAB31oTxc97oFA8p6NaKZXvsCNCbfp21DAWonry
NhRp6ybxVzJcgpMMa2q+XP+waM840eqg5i8+IpjdFs1fyww6zukGyPpViV+214DVsySt5fYtoQJK
Jugtv30mW9r4RFkIqJhDb5Kf795CaY8hx5pBK0SJasMytu3WHYH/UlG3msZ6n6Nk8a7huJVVYTQP
oTbliOTzkLuacVUpMYZgSoVmU1cuuZfia3rJNarqgcF5YaP8NZkDWL0eKaONMXpKAnssxtytrCqV
6SwMCsEMuxH1wDiDoB4SiUjxJ6Teq0HvUIe43Nb5gb5CyfSsCb8jH329jCo8lY0mGWJkG5rqdZrt
C0wSNrf2uNjK5XfjOPLFOdhP2qZjVXT3K64jS4MYrGneR1R2tnsgIrfPmwze8m/9AMdG8Y1LBeKO
qMR8C8jxtO14kcM3hWANrMkDJ/r7J9CBDiFyk+FIKam0yyjpweSoFXmvWsgKySacwoY71sqnUpYb
Q2tS+0Wnfoq1z7XPCZEwuO7fD5PPoI+DkRZ32WQWJxE5ty6P30Nj+p2QA7sT/AQ/bdfrrtG4OjSw
qX9X3qmAsLpAmp55J/p2tsWLZL+deogCtXpF491gxoj241n0Ze3SNKEayA7LtC9CPI5xpKfbNPHH
QD/tL0v6rWfD6BMAJy5DgIAQwugRMS8TkWeGRjur6DVIdYmaumyLZ7Kef1thkIxW0dJTEP7xIqcU
9k+hg58pT5ORRn/B0/FCah9H08c1LgsGs0u0i0AMoZsJ2s0RjtBYPhkyx7hkfbvhfKxzXypookh2
BPGxcSIhzSay5Rq1QUo7V1nWCELg5MOwTKK4grqzHvIJPbJ85KMNW6qIs60l9OUitTYwoQzmD5oI
qXcKyJ7rR+ZjaaPluzWhdcFwlQ2xEG9zUBE7+sEkBSSjXj/bCGiJZZtbrdbEvZO+TyK7SexSbdDl
fZUW78XhxMvHLKKAt2dilao8gW9XFBkJIG/KhH9PMeaKJDncwiuQcuJES5fRxpuI4yjWGmTHLPeN
zB8nySj2Qe7l7XhL5P2rqFFFnU/ol2axG9XVtY0aXxss/uveaUNXMxM/LKSLHWWe9SSfRQQwuOwG
yxnWVi85jup56HkyaElcnXIQ4gfPyWqsFm/XfnkhKMxTrX20Jhb4XjaHtVx2GBoBjkeA4Ckrkt36
M8/zpoAeq4NNHmfBs4cAyUzKJFjgAhgTO4fCXMg5ZiyCZZ+SEE2sa7e/6lzog3mvoIS/drxpxFPP
IScvI2btfm9X8Utsx4u1WR3a7NKc8xThW8VbQxlRAk92W9NDPqeMwdAbXfIPEgZD/becKnlDAFnE
phERXfcjo+6wovGkg9Ro7u/x4dG0KRnOifG+Se8w8l3gEVWxM/ECjmsZLD6uK89L0YfHL/K7OumN
rjeIvuk1mnkRdm1g9Z0e4EtsTzSbtR1am3EHJGPCyHs6TRKzLokBCDhuBxvQczwu7SeJthFmsc8H
uoYzH5ZwPzn0i/0nkNSRJd3eNv+3TxDTnKNJW5YWPRUzWbk7bvCbqG/bXO7LE63OoQT+Nzdn0iPH
WlNHQ6Z6AZqcCmGESqW3xnVlxL33oJ85TVP5g1ly2fS1Kl5LTylUMBRjjf32XVwM9+YlRMfM5xJU
l/hmiteHDpghxLwYzLrYc/tBTjtHcA7s8ygAA0NVQMYDSl9Pl/0V5TB4dX/ReN3ITiMhG/BiooCO
xlk2B3i7uNXw8vMw1ZvvfegzzLO0sRtg9qGQ7e7E5FyqYdRiHYpgD0wm8tb7yMhyWkO75MeAjR7o
437BItgG/GCb5A7JUxsCftF4vY76VwIEZgKz1rtNm8ZHhPjU/0pa27sSxn6M2fMzQZN4TZqIKL3K
611WqSZUuuyrKNhXaSopaLHokPd92ISTIPoZkf42qDXh0fqetD+Wk/XBl9IJKgkhxqwin7H5G9mh
XafCnYRLnwTTYvJtovR3IwKx15JCS/0gatQS+nNAyuYFnf0FM88FA35Pc/C046D9I0yhxV+x8oIh
GHZdllt6ZeWKi+29k+Obg8lJ43dEkDNzOOaBi7p0DyuGFNZf1lBdGeeM1aQrvvtXrhHQ02MVjrZ8
tNe1Rwt8V/hJ6IVuY5PLJ0lRE4NBwvlaB71/ltu5XUtyuLxUFZsP72WWFD29rGzOIBgY1p3iRRYi
VIA2Eg/JZ8lHe3lVkMwxSWunAg7uL1eg7/nsRWNcdn4L2VpfyP6AG4bE51pYNZwqVEmcFgtnhPH4
MZyHoI+O2RnbvnTQO8hR+vKuhStvm2dzf2LuFhIEXOIwtxq5ORR/iP+wKe9FVpqQ7Qgu0kVxZ79b
B9LrIgHQKFp5smOcq9t/HhrX9KjOJd8yT4RPv7/IMQBpl5+rjaN+Y/A+RnHnyGbG/veRPn7oMj3i
S2pX8qmHS6yOO2J4MatM0mljROb8xp4oB+gmpy+104v35drCxBBhOOwuZn0zRo0AYh5Jg7uaNrKM
UCOr69f1MSmlCln+jR0UZzTFNpBmlE8pE7kU8C8Zzokxt7bZ2swReZFOIKWIvELNQ0PmmW4QIxRv
uIf+DtDnw3VsbKeDx+WUk6mhv+UOaPBkSvqnwpAf1NX6iI5d7r9auXJSP8HBx1Ag0YFaV8pJPkSx
PVtpffVj+BauQAaXX36d4UuS2xPJsC7aaVX+VWadd8/LBM0Ta5gDhxlUOol/34KX7tBYLNU+GiIl
KGg/8j8OC7i5hFcooMqr2hdS83Iin6AyrlMlLSQs+C1EHdulZdakpuCD2eSMPbuAQECuYwLwbSdO
+jZcGeE48tEXacTbzfLaXuD7ZkzC7rB2iTZhnuihp27Qlmw+7U0cpzAjqHeEmMCNTbx24MsfW8Ep
hujWyC03JcYRUU3MkS1V3Zwv7MVr7UwTLoSeriGMsYU6EaQbcG+b8R2qi1+/5j2mSUUnpFBDi06o
9O04WyvfC11Z1v1mmuRvBPiOAbmI/mtaWrnBu5Dut2sY9YLcFTJ2RXcjgemkF676eW+2XC25Hka7
kpwUrBIJFIiNGupRwsEKcekhwGgSuTxp6DEa2fRlNaN0l4V3cUEk8NbicfJNv7w2UmD67M2mI61Q
98nZ5ymPes09GvAYCkxg9jIUZ4RG6EPyheUZcmepXREjkJz8QaaLg+oYzKOkr8qAsKdvApjl87Yg
Ofjc4l8Eu2qEJKXsn+KXp5PvbN/Fz/IeTnqcjc7aKcRxgoVPJQR2pPpv1hvpRDWGb7qkZ+p33kH6
bT22GD11jAsxqZtAMRZlpuLK6qHqgMmTJmc0Zd7UtVFptMDPHYEMIwWPUoIC1mI2vmq/gmzWWQz0
hbWd/kQfqDBS7JpAjf995nISzYMqeILiEdpounj7YoLiCqGfVOn6b8QtskvgTzok7vuOjYslzWOL
vyfZlrcy+CCq8FquiIs2bS0PobheSWjqqRH57DdkgGmjxFbvbIUrexe/hhKnWTQ8SBGMRDH22dsB
IZ7VI4J+BZBTjBERh9ye41M2g2nampQcTkxNfNalRvpBM7mCCBQMROFEpXDyh8hcH9ReIkfwaBBm
8udpppyzgp9JE6qbCbNqoexx7gM8Ls71dkOyT77jcMKmLwRXgbQRDSfd78K7x44jF6PEHAEDLcq5
19KbZF8nLliDObKV1H4GD/wnIzun3IQ6W0aAMeqzSjk0dNRMsG26UEFqHMr1mXAuZ9nBrufPx/Sv
rDqurnHe5M2g2eJyRXmyGAO43OHQ+hcd6H6odeIdjiR+8ZI75nnQOIYuQN0dyT5e+pH+QxVIdwLh
qA4+ZSZEjFaIoOID3oVjHs3ynIqBVpi6Q9pNApOtVnxZTDeQNl9XJKfKdJGc7VldljbXpKqVn1YE
xgskKVn3K945inJ3XEVjIIMqKnx01k9DyTbBiPJZYeArvWa0WLzB6XHn2LE6GgjZWzOSdwPTPYH5
+Q/bWwgnuIEP0Rtpdeq7ut1gFoi4b7WwxxChLIm44XsTWMK8iPwAiSoTgpRdKq7Qyq2WbQHt5QOd
4oGh6d7ncpdldDNeb5rvlcJ3R837CIFxvucUMvYr3ksEZLRcJivVtj6/IknLX2UkdU5DPq/KzH4a
A3yHPho3xF+HvW7KvBHWIY4cLPMlUfw5hUAWYMXDg7b1plpW44Y4fuWpNJNkSwO+WVr5aP69BKLG
6PE1EKC54GQaSfBAfVKoncvmD8bCuBXqmM0tUqxhyO09qhmKM8BIy7PIle74g7CRkI+ZB6aUMJQ2
8uU2BdyliuhycBTD5onedqSeCEsQ2xjViKxBd2H7gaWRkLW0VyHDlS+r1bjDCJJ6UvsDTACnErr8
/qI6hTGrqYrZYvpCksGRmTLkVuTBSqPeMQQm7aLnbiIeqIEqLVYPt6gE4deLU1XBzypHs5QQrDI2
0Y6BMVg5Wuk+0c5r4foKQsyrpxW+1bZOzYc69B9m6GTvsKUPnj/INM/UKKaUKzHYyLFIldZnXLWK
uPpVHd6WiPrd8K+n7Q9ECCW+LtepW+keIjHU8+HJvswoytT6m4e3q2Iy64ct3wEwP09jdk4t/Hba
AViqNgGbLl2et6lkySvYRZPN9Pri83ziJ3I/Xk24WxwmIuzJbhT6R4cILCYBhfiSB2bpLDvfJxRG
NnLFri/zlqmu8AU1lHozg55YQbyakxU7mjdTfA6wc0Ew6Ce5mR1edyZog59YAQsBGudrOPae2zJd
so/rE2MHNjG30+KkgLlZagmkmX5TMvwxd+9b+NsD3et/GArOe5p14omlHKRy6uc5THVdZJ6FaGWS
NYFyTO+FwwtbapCbR9J/IAPooirLLpA9iiSv9EKnagwbbpq893re8E/7N6BkNgcOEEdMSHqtALkU
FFcq1LFFlNNhBBn9bH+gOwhgxz9AVYtHNUPuuxR63JpNCWkSTg15BPJwZKnmf95yldZhLf+lKF//
E8Xp9RWtJvrEQR3/iQ+wbKckBJvqbTobICy1/c51u8Tix8SIB6VDCu9Vp/6hZeX7+7GeE5T8/phJ
P3l9cDwOv7JnD5Ks6QDoVPVeWZLehuNKIs962i5xDio1buROIZMjoQAF7fwmM+x3S2tHCztOTOZr
FmRUn7/Ru29RpwH3WEl1M+LY7abXAD6V6t9b5zaD+eIMG8BhYBFsgdH6wlhc7ONx6oEUf4sQGelF
JX1BcKcEL4hKj4d3m/5S/olNLZWqfqi9gKKpPh/ObJA3ou1RDZDCkeqv1W35p9b/WiFYDzBhlQW/
KmzAc9ryennLnQ1ehf6ZufXbDjnocA+lvz2zuqzN1pJhBiI4CrvnclSi9++0+5Fve7cwhPz0XlbL
6pVHlU8nsldjmkdsCkV/zqkaDQrmG1Jx5xIoaFY3UqDgGQmpMuxOks9re62m0i2WEhObkJIsJp1x
RiG0/e+8EB0V/NSo3VkrFWc6A5aWO4vlYvDp398FwfcPv6E8r4/IoFggUYbWYfHwoBGGIViKvGGs
j1lz5odfS0yVPygu6UEod1+q5JZ4B5FGQBMW7jsNxsNmXcEhFb/x5LyKW99GFlS3sYun8dYdgB88
tXUkxfVN/J3TK0NvmKGixVpXEokW7WKYeRL0TpHGlOVC/tj2IIEbmGlt8+haZjrjWhsLaUtDKkgs
O1FRHuJxIdwGFxjCoZ7SzVkgaDdsuuOJb5EBfDr6+k4/gVgldkE1+OBwAGKHDV6OLO42lyK7J2Xu
grVghzHGWoPgsXkWaIQeSheRip/njWsExMh0zn2RStsIHOwtIbluTjJnhGhDthPd4ikl7fLnzzTD
vCSNh1Yz6Y9Aq3aY8cBxSpAyj/3/K7M13OxEgO8/gyb2pXEkKRHwleAyNiOzrJBHsXUfQV7lkhBl
wrcWDAwleFO0tOLNXr0PEnA+zILbqtV6gnfgT3+D4oAmyHqddYD+DAaa8AkzKPPTXm3RZrJiCVHL
6V907GsYWwReZTrR8d7ufpDkMbSsuaCUVu9O4woPq6DZm+AA4AQgsMS0PI5wDtiNf71ncV/fDs60
c5MMVmxSIIiY4sPbuZL8Z4uB5N9IU8cniBQtspwJmO2sgvwCTTTSl/bC1/n/wjSOpxREXM9EDGXk
70myFwCtXBxjy58jE2lYD+HYzAsPDLsreJnfAV64YLktaBrBrdLMB42VF7kumvak0XtgWJr6AZ3/
D6GOogtxQ1Wu+Q3+EhfdkBTUq2fNE6Qwlqp2CIRzzwNkOm3adO4XdeVifXL91OqFQRX/IyGQhshi
HAgCwRrg/8zDHPs0wluGtdPtq3BZYE6CGdW3iQdy997QuuEethXzHq1S9XhuLlf7HLi7P6clVbSv
3RcFgpHn+R5BJMX5X3ywq1NGLWvdbnBWL8GBFyUKjkGxJ8IF2gGBcDgZN4W6k1l/Fh7avOIJai7x
tcl8DEdqztzKgwpekh9+CeL6Z5M+sp6vnKSdD7lHeJQ5gB6T8iojlPyOje9krzeFK/a96BZQDGMv
PUB/jXEQFFeNwE3gd/P27NZZGht4J/R+n6G0YNBSP/3Q1wA8zlMPlj97vur6iH9oylbnMg7/nBVn
DEhiyfOFwUry4ztRTMlTxTQfWA8+XxYeAs3zx5/7xPYCks+Y/azQ0qxiNAAnfzdUvdAqoarRuw64
3Ya4Hr+Cqy1AAmlobEFUppanDrKzWLlqIkM+Duk2I4mFxHhjl3+1nDlb/DHL46rbS2HtMla7jcya
V37zEmG62SYLBvYQl2RYWj+waNED8vNhYaK6MSB+HRS2+wimCNZhCPW4Fyv2aVN/M5yMqkFJwqG8
ClqIDcKjDBpS5agOO6zcJkfXWjHWrt3TKnGpd8iB1BEkzz4SuLvDOj/s/d7gr9b/9ZOIcDhDvLDF
HoykFVs0eiRx/Os438XhUCi1UYX3xmNESju89suKtvJb+bl/s1DUYbu+AHXa2MpkHMg6a09Yh08m
o5wVtaZ6Tn5r2y8XGkO19quVbmTMnDp/V/sCun2Eu4Sve/PIcaiKiW9Ch/Mm4Zs/TPHDUvmlT8As
4n6TjAiLWpB36WhUPVq+V4f6zOy7h+YhRrIdPNS8mWGLfpDJwB02oCghjqQRFlvq2grlchWVSYWd
fMLx4ru3Oas3NCEri2Lt5e6sYgwWWcD/KPxUjUGKYvxU+0oNeGmkHZK6Ovw6ROJBmllGVj+DLwLN
rtyEOVhsXfjSaAvzaQmZ0B19OGTfOQ3HqXgwBiVawpV2FzHjvnOP1kgYYtElDAmsMOJ+L6aDiWzf
jxBgAoPoIRCaBlwRmvtDRfobgtX7jesIh57QnOBrK40de93TeR12hUlFV3gXUvXbKCcaO0Am7WcI
LJEWvrcU2ibCtyWOYwcxsAoBHwa8eN2BpqikD0WNVAMBZbtVA/EfbF0Ol4JNDG2G6iPREpXgz7BZ
oTVD8Xi8WCirIdIkEDF063XlhaR4TZXZcQoIehZ4+atbKnL+qN3uOCBt1UteX+WhT87wGH6bbA6g
vA8CGSh4PDUSYgF/ncFOIbFZdhvZri1P6ud12f1vX4h5T/4bCPT0xaHEYg7NwIGlqkY7UgeP9GC1
AD9rA2p2v2L0OKriIdXWEU+beqTQQh9pAFfuvYXuH0KsxkOGWplOjqhNwjxK+UHdRc1/x2BKJ0kh
rbiFd6cxlNJCeX/bwYruIgdtactgjP4OQYSXszMiPnkxmbAGLWvJm9Lag/qESDttWXdZhW0Mxn0/
yVycvkOI9EvNU96XpsZ9EE9KAzgDjhJ6GHHbQz2MXERCbogJLNCSS7d3+Gm+2HE9/HUyg4s5puzV
rI0SWV2O6LjDsFn9k4pMJa2QT6dY0NtWBNn2b1UTP+ic3V8WegOPx8OtounTtdJBPH/d7igL7uGI
w4A1DsNd5EfURfJk/ulRxchqjd6SJcohY6WtnLuAEAiowVrJa1GsesUAWhX3XhApECbP52YEGJpZ
90YfnicKWd9qmbD3TXYiBKIe+mEL/JfvAfmy+PS+cUfGjmZ9kEo+YFet/wlQCAjhyAvZbDBD/0th
7r9OgoA5QjFukToirg0Tko1D3GjLUzgQMphHnHQscmopco3mafHzA0GlgNedFtKeVS3z/02JoRX1
aae8DFxDZ8K5luiUMXRNNB6m5MWOpVln2sFToQ+alfVslqGWE26JVnmp4naWnSkK3/q8UfSkH29i
VOBTePrH9kdJJ5OYY9gFQL1yQcRze65EiLGyp5vA5LQ9OshX4eGkcIehr/LO3u/GteDkqdFq3dtC
WnTn3cWuomf7qk8NJjd6K2eneSglHKn6dLcxD2zMSV7U+8Tcso+EOdJ1PLqHqcgMdNj6LJFDMV8Q
H/Ag26vavMWueRYsbpFu62wGmWB3sDqjt1BSfmbRppZW9ArpIIQSaGcYyXdjk/8eTB8NGI9Jtz4m
VlcamHvIJRMoIJToB3cjT58p9muZTHuHnG+f4bEVCRV5kfhi9T/651Ip0uqkq6LXa9HKj9/o5p5/
5u9ZnDNTFZLRDlAjE0wZSEIJoQKTgNcdN8OPO6orpT2QeXtTBJvQD0Gk7B6eLBIIHkMxz0qwm9zA
5rWTcJEjlNkW2Cvt6IuQPGWuKCEsay+hqA86wvHfXAEz+DEN40fxRXE48bWXLslC48mrVbGWFd1o
AQq5G/18oVMiGLbC3Q9BtwHK8wNf7kT9eBFc96XCkWuhJW5M/ohg4kW+wbMtHLSB6xCbQuFhkj3q
Yo8hnsq6cZCkzPmcE4sy2R0iKi+9oVNoZ0beKIGcUbpwtg5mQFeFHdUnisf4GWe/lE78rOlAvwhV
OcY6v6eALR4jF2vVgiQ6ZXabr3cNfH3eFq12DBBUi6xeMajZpsQ4MPRaKlxFZa2soJhAUamxh+hS
1wOBsQ0A76C14rEZytzavGCSIH3xjzD+LbVO+xrOYBahs2fpIemYw8+a11ZTEZ0UnsWhMLNFiKC3
OqpRFBxSfGzsc4ZTzumeIFrQlTfvht4VjXj2y8u4j4SGGqyp4S/0fkC1WDKOPNUa8k6aOTlHezmH
AIeIxF7GZIkX+x0YtjIVLc+7rp352zysSWQ9P4injw+HXutUBmfUMha/8dpJLmY6zY5IJWlFbqcd
Emcbfwo7UqtXmfvgp4tiIIJkGkJ4z0NvOTXNXfGCJv5WbfbkXUnhZE4UzE8/NR2pZ/TvZv6UJPQX
j1QbKadY7lNLNTgUOMuiaqNz2t8tcxwOKeLiiIuuvdvu9O04VfHe7gwlr1CGgri64tffUdA9zajl
CiKFWwYG0MJk/u4wL3M4Php2YFkvWwMxy/OYVo3GOh6rTGsfnNY8s+AnvUdt2fw9+uERFNJg60M8
+HiMKspIZzVIC7SCt7ipqxC8fOASUvwbnlJ3ql/DrmxXnqSoch9iOotrv6aQbgMF1Uu7B640JRqr
PDrCwQhEfrWzwoT3/tb/W8hdLaGraOCfjsRHfKCpTp+dHlPb1kaKC/Ttz6MADxUQ4jd0s/EJRjRM
r7HEbUXONWtZCqdF8HqYmlvU5f/R71JYQewIg86C5D7FP2EXGLe23BIhpjRl9SDBc6EjsSTiG1UV
BxmOWPVELhsCvID+GR1KWytIVSZmYXaJ1LW+LEL1fkbUDlZiJ+/54bGjIcKq0iDCIkT5c7qzN/g/
8nMv61ptfRuBDW/AiaA7/2kbD78qBa8xxTncW79G7CIlsvR3U32zudFOn0LBWN09FDYJZG9V5ouJ
R+mIapBZ1+MDFw4GDdpSaZBxwvlyVGWR8/RNtbQ0BQDYoW+5cYApt+lYfGCI2UHWTB6mkPxAdgeU
QeaRr760kMdLcA4iIqvlNPuJMbqSpOwN58PKpYhf7gX+gIIozCDIu021ANA5Qg0hJ7/agE66Wa/Z
8lcDYicPPcwcT9botq/v7SlcDrtWT4mWBm8UqKq0bg1Oi/y7RLHExsmyeBVUP6kLpjdSdvl74kNu
Me73RKf+/Ep5iJ8caL682wrL7G7Lc9G4glg4iHD9vOf3GBJpLd8eavMj9dzTT03luFuX8i0pZ11F
SLpoa/ahvFxuyvu4PxKpyO8oyI9iNfdFGLnRmHPk9jP2l/scvgUlOTl2j1wtBtiXVkISNTjFTc4E
oon6pANu7K71S9tjlzLectfTW9jf6UX1lSDj3Z2Ei1ONd8I12UIslvHTiXo0jn8DANPHvhZv3qMy
V9dlQeObxUMvlf6XhHI6JRiiFg/CUQFw5Av108T9jc/lKandwBlKCXaMzOWTu9ixEwv3T//+DlfQ
MllSh27YZw8HUhJCkRqZajr+eblk8Y5h0ZHgXk8xmsCeGXyRIUWPv/9dNQ7MsO46Umoxg8M5rjES
po7vzvtll3zsU5rxgKu4ivzIEV2k9k8IWrKcpgsvFyO4x68eyPGVdPuVimoy+wiqcBT/NQbId18x
VYkHBoO70SLy7wjcPQSassKngZONMqT0yqzwr5AZtnw/uTlTB34QpXUXLpFi4BORMaBVwz9qYrLM
Lc6RZVPQIzhahLHWR5rGaQGJTLn8VgsggeFwr4mZLZofW9M+KEwrdkCwggQccOW258c93k7F0vLG
gUxwvooHglC6ulL/vZYBCeYRA3BSOJpHcdCM3YAwLIe++TpqPz39nWn0R8RXvclM0TGoF8TtvGWP
KZHDcXFo14/npYb/9yLi3aSTrHArQl++vmKSi7AdAGq2nKJQDXCqyJAX4GohMsuO8JGxs3lw/N92
f1vP91V4VJYeyR4/L9marYw7hBAkDqLhSmpD0dlu5Vuc0yPJUPJaECuBToIPZ53r84fdZobcz0aF
pWxb3czw8qSw6lJGFRoENTiYS2qxZYdaG1erO9dNKYEVL3TmCxC2cNAcYAol2ziAqkfUTvh2O70L
ZAm2Bdx0/YbMuqa+S4mUK2/E8t2kBM0k/gD6H7JC1x8DoNuuXgVBRgiu/NBaUk+w7iIH+ySKiVx/
61gwZhJEfVwW30/bPgA8fUs4cnLRTVAGYVKdM3KLGzWmtSilpdN/emVVyuuKCpvjIV9t9JhCJ2PP
ql5pT+E5zL4Ws+rI3V17z/DjO2q0Y27QRa7uUvqWaHCRcjXAZW/suQaEWIokhTgIr8OMONsONfRi
Oi07v0cfkKjsWZ3QJcxNUqcMmWe5qgW/Kok18FrkCTz2le0xVya78JRryrOf0Izba1yKa4XELexf
SDPcojTHFqk3V0oRUnQDv9dnNVHR/6Y7x9JUDpVBGRp2+YrpAJEf/Snwrz9qDavI6WEex5xBs15o
NIU3SPlsEaPvrR7s4j7TQefBneSrfMszRWlnm2/SdNiImbSPYo6lFv9CkzGTSbmpOfaj3p7NBqPi
wgIetspd3uazttz2rUBWhFUW65fc9fnp/8g9bZ3D2GPBMTwNuQRorQkeyfQjNmVsE9dB+xOs859H
HUibbx0Kypl5pQuQv/4ERZIqIrgQJctxVV3f1ZWwXsJjryHHNj1J+FW4EXpSVxutnpCT80m6D+H2
owoNFjLot/5UY6m9aQD+KDfW+mmTaIovpxR+SOPrUyocpbMtps5Egxhh0+6xFGCVWzuZIe7s1jJA
kTkZsXtegKCilRERF4I9piF9JmcA1lkAJhP5ETuedByiNAb/XzmJ0gFicVhziZbY5p7ogk5L9q4K
OqJ+LgZmLDnJANJDW3tsHul2hri34p1l8mqKM5n3t1P9As6mvzbDGj41r19/E/zr5+PSCHmClorj
5fgQX/qV4oUccRPWzNrQzEAqCdjmcbg0rLa4SAJCwdET71hKTBiYz63mKZzCUidsRvBJQuiIBj3Y
QIizuXVZLn9iesnN9RHjFufaQ6VSg25b/f+F1/CsUrqPbgmg2g+n3TnXqSNnnligSy8QzkyRmC7S
reIy4lxFlXIyzrtpUiAB7C+Nk4VcGljFcyDT8f1O59mGqjn/HZ452WyA6hs1XFXOketJIsyECgh3
roPs/oKBVLobYeUP6I+a2oa7Me2E/1BxHlTadIPBRbKqibZ23imDzgs3RqiED2jEyLRIcu4hSVK7
Pxo14aMN2pPFr+bawZvGrjtY+oXY8yyFan43L+ZXUC1jWaAlsaOZxNguaFBlktxc1BTdiXeCD6pO
7nPggMjzJ5i8n0Ov8BHwNHva8AOCR+CilpdtL53+hfEIpmvV7j+5LDHPKnXi3b/lIAmWo/5pktot
u6S+5ZcjecEXr/8jOdprpUO5gHvCxXJkMn+DQ4jAG77+0tbm7FiW1+FsuJLtYkg8aaKxOAhfahX5
hdvXik/JvFEWvty/s57XrfPPC6Zc6EtnUJiloGzqupPQ6OWF720mt0kJS4CgBXtnVhmIxkGwIZNS
vNJ3Y+5KHOEPy0kBjRL0vfntTmEJFe2oeNRHwrM6GBC4ITOC4W3Ugtm6oQ3YW1ThWhUJhGdelPet
IdmfVqrAbz2dtWKvv8s4cLvb5W3kNhOxpzNUwdVIxAtIzAtG0Hf20zNd7b6YgUd0E5Xspc7/zTXb
sUf6H/9ltAgiQrlXjOM/bZJGCVUGI6bkxDO9SC14Ljh85LTqMFRxUKRxWRpyv3jUVjpigvZQzwL5
9Q03BepNTUu2ZXQJDm+GSOg5R6nb5dMY/K3i+20zlljLmqAXGhN65a7Ms+R6klcinqW1TIGN96Oc
gxrGTVUt2Ex4sxj9ROZgVaEAzU2wXPuBrcuAriFwhPGqV6jobhs1v8vFcohb6f+J51Ceq1pUQyy/
ojFEVCSDsZ8ec1KeqymnQPqqBYikb4VP3NjiuMJg3ABWXNtzLWayDUISFb55pri1Ci6NxQjVjutV
32mdTmUb/wyFiQJW4OyAjCJBl4dUhmhJodgfKVasS4u+/5yZ0AoeR+56NT9B8LHQB9p3QItGTzTk
YyJdgOfbPGfDvh7v501RoLn/sdxmpwhtWGhUM7tFzZLRF1zvs2corrCMDzxSXS4aYBXF0eU7eP05
h6XAZ4C1oZAt4aiQwo/4cPU++P+OHNrNB6iAz4ubfEf2c0+nJocOogvPEcOd0+/35Zn3njz2YYiu
5H+jePEjMlAVze7BshVapRPjph1OyaSZ90n6OnoR+SGywtNrVYcMftn5S7L2Hyb51nvV5/UJOfMo
GZ8nvjYcoSVFAMDOI4K23vXiimlM3olHF39XI6Dp5Rb2U0LbVUDvY9JKlDgPF+8y9nEYxAF0sMWB
YqSCCAUKagOX+vCtDqPfC3EX6STqT6Fap0ww2fQBJ9MCnlkPbTxzT4M5NSgzOS6BLlmfI5GnLUpS
R1FEbM+RcScl6HmL+eok99mklh1rVaB5b/dWeCzcdLJhvhoHQlvJH8M2fxIffxiipcA6cAEDG1QN
XJ3ea0m3ipoMPZGbBI5JfB1KeOzmTn7+WNXci2RQSwmui92HZ7zCHI5DQ9RK1o07DEAm/gZiZnwH
5AbDJ7Et15+7dDT4m0i40+kssEMv74VT0zR1gGWl5Dnl3ckDYoeWeY6fJ9LrAd/+KjrfE4UJxe3f
TYiIvoqpPB+kA3nYvguinAz/1bjl/78c+U8ZlKjHvM2xuTUdOjNLBPHfOC6rwneehBF/bno/a4oS
S4G9VyRq43EJMRqlA/65niNGgUx3O1pYjV9bMFylyaRXpoDAGqqWHwZnGXWwQqhUsbqotMsxLG/7
SpAS5wuJ9urX1EwxynYR9SvHGlLgB7AP+Lz+wI7d2rm7oafLw9JsBIdCoMY/tc0/wsIqcqnD4InU
HRorWKNA6l1MQ6DX0vggMlEQiMaFihoi4KMDNA6fTBLC70b1Onz+1mcDkHcECFsBULfrVZqs4Xd8
IF+eeqVXAYsQpQsZ0fQdhboh4tLgYoZ1l7cFxqZ3VVBMKsGJfZ6Ndphf/5p4cVBRn/99uAQqMOSs
ibbdn/2GVBbrSPoqmzhsRzBjHJPuvbQnOjLuDkR+a7K+J2kJx9KAoYZ+K63EzyNKV3MqQahWJ+d0
M5dtWE57/S+koIy4JsXieiCCvrsI94FkDpIPigAzFo3zDEb6ARk8CvbDmnnohyW3KNQnmF86tI+p
mAfljgRilf/GzJbgdVn85pu4GWyXEbDmwMv8u6rug4D7TCvDv+dkpNwDIqlBZk7HtPv1g3MMqC+G
icg6dUha04R0WIX6ofqLNva424YryP7GhN7w9uyyNedYA4cAXUyxTlIMp4SsK6fqP2LOXI6VSa/g
nYJGFVV0aL9kHsgixXfpb9p0tYfyId7Hdu77mRQDnqKbOlf5PazIFdkbrX/FZWMKJ2xVvzNMCYO9
T9LN6F58Ywzh5knLPHX7XVSVD9BjlZPkub1MLfMgnuL4qaH7iBi4evugDTlDxQJM+IbA95AEGqal
mR9lX4iQi0iqyIEb4J6HsyRPlg/fQMLgWXcpk8XxBkhtbw36n+ZYYufFi24f/440uc2yPmfFeXcs
ljW3GdLdBJVGYuoITP31a4kelHYgI8AaR0pd4fJdIBA8xPShmxWBVyJiCYQQ9WpzGoEPGcxaBEgh
KtfSJNvgWBRM+keDIx4Oj41K6ViU+7grmKkCKyXRcjRfa1ZwXzEscak0U8S3hc7p+/cXtE+VmZdN
dJ1qItkJGj7gpAew///HqjZ8ukbxNqzpIk/JToEBCKcrfPSV12o3V+X5XwavqiPIYyynouxUodjc
MOCYLJ/z46XSkPuUCrc0akJAJTsyqAbc8gogxina2PTOGCef3mAk3cRjWcyTDXPUiMXeF6MH8EQX
omsXibZUKvnp6p8KfABxw8QDt3/BWjYgulS5qEcM6BQOpvxZkBtWbV0XZR88Cj8ewuNuOExSSCvh
foMDgeD6xwUtVW/Yxi/I8uTEFgOAKYleN6a8M9LzqVX91Xgy82wLHJ8TnF17WyY2fUVkOo3is8po
xdswcI3PLXiCuZcMvLl9Jo6diEDm4PWRVVJUMgc/V0Dv95ZmLjPGDK15SnxH6Ia2Fls7kEyCp1Al
NXjgtEUTQCf0+PwXTBwqSo5pd7vHV9sEUTYwMUbhpeyGV8P5Us5/an+qJJ9BnDuv9i8Qm28zFdA5
69lV9wjcyYgvT9xtqfFEn5QCGpWgWL1tuRd0xY5d8uDrEMOXTuDzmgHE5DCvI/Qb6P7+BegONOlR
4Az5K8+zKbBsEwKnLfvTmZEfxjIOvV42Ne/H538HcXntVmLFkODCmnOyIkLLRGclDUStGtdM8rKv
x1CR+cyXByCmhe8t+mM1rsu0/I93QjW1PbH5NGYwiTaq6UrCmzc2mVeKq8TcOjxgYigr7eOMkJkU
DdiQt+AklBJOn8/SwYa+Cy+f9nv7UyhEMo6IhhvdJ8aNlWteCgMe00HY2W+PLI2QbU0Jmjv+ik1W
URQ4092U4eG2lFNiGt1OwqkXs4b2ttbV6KhyZd+GDlsNgtWDPjINHkUtoGxyUmCWcqpx0640moBs
KO8DpTlNe8k8qL3YTvl4+n7Zx0CExTET4gWx7/esBBzmsh5AnZJrbS24Zcy3e5NkBtzS34rwfMa4
Suy0tgDoJ7B0qSuGhtVL6c71NcBeMoi9mZd/m6ldfKzzwuTunpC5NhTDqFSUYsuZkmdlKG/O0LRG
YAk8cIf7qP+RX8Kzx3i1dZpLrfEW3MoeLO8Y16XgfqQPjaxfm3/9ypWDdsf8hASMHMuE8TknZGi6
kW/TjsZrAFGMd6tRmUC3Q7zJjky1WM/kYxii6aWXLoBn7UQHLz6VPtMeYsqax+izssOwmiA1gFMa
dUQtplKe3fx4yQlZjKjimu+slwrhnnwjWwpOruGm09BlthHxoQpU6CbRLJ4XGgf06CIquNM2wBUV
52ty92Uq5oDXXGxS69eOTh9inxNVGmRYXFUfbxsL7sKUUNcswX7bKsRaxOSiMCbHQFpn28d709Sd
oBDqzBZLUKIFS0MwJ/eugCA8rFhphznAa9IzT2Dh1fbkB3s+DuxHhnE/APNLvL09gQpKVTsNo6oC
qKWaUfgrgRTAwJcoSUK8Sh+reGhuo4dz/JBKtuP04JaJFcJf9RfFZdTsZ5PNCrL080Jp+vuK9GBN
wtqq4ViKl4bDo512IxDRZVTXtLwQYbIDA02MSPqETPMjIvxqOnqtL78C8DCCRk7CAkIf73GVfOV6
9gAlZsDNvj0d1CfvDMvZrhvwYaVCGXUFo0+lD4WafaD5m9MpJRbNljNdmgrGtIBVSwqIsDwkHc6z
7DRHcM+MJRrp9S0CQMBKMPFPkyV6U3g4Im1JQFyfo/vaGC8yTN6Z7wGQEKwu2sJSLgevBOJj0RK7
3e6Qni0TrLeRebkCxPmnNAnyBCKWl1PBhP1IDltGN3wbNGr+SuIcdzcax7Wzg7vR9n071hnXqKzb
J7ggAveqaPqJnf2s7TR/qQngIJ6nBFcgPmUCQIGdeTMoyRiWnIu4oExySEO4XL/u5Okgm5CNOEnm
uA7oNA6WjXjq8go9Gj4lnA0brFFq6X0oqCIwNb1wd3+/7iBHmsa7JCXkiNYt5fw3QFSBb+xisteL
ZHNkGCaZJvWRrKBBIGmB/XknKdo+I+3rwG15v3H57pZEIaN9ZzHv1PWSeI4I1WhmsBSzyBrNWBJK
UpSHTjyqewb69A1palJDOWXipVKCFVep/GVSehHEEyv/d27FrkzVnD/QXRTWO/BfyVDIqXSHnpAv
v6Htxv10cnm6Hj74HjunY8UwtIfPOzfOD+jZnCTIxnsAatzseNYm4TKiscyvvZ+PFwLnlY+wDvOj
/VBI9P5wHHbcdYOdnVymN+d2een2zoVgrlTwDqqmqseWuP+AvTcMV/UmaUaVGKHLB98dB9I1VKMr
usuaSahD1LTfkXMbrIEY7G3SvhanIrz4OftEnQ7y8pdxcpuVqGxaKB1FpqG0Rzw8rxgs2AQehvXX
HlYSyI+xwG4IrIJU0PzLS90hG+c3h2R9cNSXp3gMrBkCx33V/1c58rv9vSjmnO+X6YwfcvIMrRpn
xNIiliGT5nvhSY3ZJW+hcM4VyvvAYLHVAAFEkUe3glvTKzCrzjw1U411QRBEEMfL5APNyu4Rw1b1
0LievHlf60imTjuX1wqaMJi4R4qSLt/15JjKPJ2A6Kn3KuUDwnit9ewfbFOtXWcYAERPKCJdHOuD
gmscCQcb3cXpPMUwtwpP7srYjo9YGQcHLY47K9oFlc77B96rohBzEwQuVN0pU98nCYjmxZdi/vaF
40MA333AsBFXUjLThrhA2heR9LUCT1a8AfB/pFWuIv5BzzMJG9AfMxT816AFsJ1kNmOwDXn66UJ/
mFGZtQ9Kjdpm+0TgF8eRT4PKZJNh9uT6oTExXXbK5PbboYIM831jbPWjZqxosmx75cikLXQVtAJr
MGlUuD4f19WkPdpr0M9cJVu5MDEBIhKhD59NQMGhn9SVMHbnBnyZHxXSaDtIbbklp6DcBe/EDOmk
wNUE/5cOOhtiuFgxFSn8gtjJvZeoDqGApd5fqXQ8epTHVZCxm2Jp32uodvvlftV8x2MbFEZln6kb
lU+342lDw0lGbAlbwCEgh+VU1GykU+4XH/eAIgnCKJ46oC+gXi/DmnNq3rSZ7oxKA+Xm46Uds3cB
7NVpsHCcGJFBONGWwhvyD9IOUA6n09VsiWSvPvECMk0dFtLEf9TkJo0kwJVv6P9DQXvifaFOknSH
Mmko6w1m523EJOOhswWR179wd/gi3/d6P6nzNRNWoZIwW6UReg/QqpmP5EGRZ2tlENTMeyJq9zzo
YfwPse/02r9CjBVKzf28paYACa3hdekUMwa+zeS33Xq6bMWE2Xv9H2jVfMj+vPfHtLy3+TpGDgfE
7YJkVVYYxQyElv41uuTm1Z6+5mdDVLQK+j2Xebhj7QQdhAgoYiAbNPqfNUUW4e7CdjEh4tH/ZUrK
8SS3IhVuYY8ObUyk5zvZBcvZqaYrm8ZyWTbxAnG3KIuwcf/TyF6h2oR7CGycp0GOshW2bmJ2jCPA
WzH3h3knVKRIwIXDpRwhJUJjx8ElM5ayA7gwy1WtW0XPCqqA2odJhvFCBgJbRbScC5rVrVDzmJDH
KGyybHbdXdSD/hlEf1VEXFtW33Dx35Nv/5Il7tFxQ7euIYt+CKEg8QHMWSogWlZ2JTQonyfqVNLb
aAl2jXXSGcOToFaDzniOzQjT8kpWGs01b+n+yTdqAezUWUD/82kW5aehuhSpRKeOk4Gx5QybP5QP
QzAUBYS8+StUE+K50qk3x4FO3DQz2WOg0+OtUdFoGmCHDpyIoazAEmrH2mXdl6kyslDKOgsRL5XT
tbEYkCwfBOmnv5mF7Sb3wrczr2qOmcum/0mfzzPDoMkSkNxpf5AuSSMevgomL7BzRXJJA3EVo3Fw
xb/dF9HliS1MqeVKOYEsAyd8/DZuEb+gG5Ws6DbuTEnCfcobBSzuSu5kMJvAx4+DISSsSMXBoR+G
8nb0ciaeO5cpGP7g/MStXHmsvc3VJK2vKVxLIUYKLuz4L0cJpUH+J1N0w5RgCZpmyEcUS/QqupYv
jOpGhp6Q2xCL9Adv8wOJz/JvZjPmz0kU3K6WSNWebegtB9cHbNE/syPTwegtEozOg1lZBGo4yQCz
MYCYbB01vf+xWqq9f1cdaHxOfH5jxysCKcmolPB7qT5KKcPgYKpZzgG5iZtPyTszHMAHW4CgrGmM
srypeeuTFgEsPMTWTniKVC4ySwe4bjBQYLLpfqNWMpE+9AiRbrO/Cig3KbtOQD7f+p7GkJpq+p0q
rKuCcZevkbDlgH0Iexk19SfcjMu1+SbzCcE3rKUEOmLqklrIZ9jQLT/xLIp60GizXRSvBqZEZvRD
oe2r6NdHFS8StZNxDHX8+p79n6gOpoW7kIp35O9YOkkfPqLfQ+0jso85Gd+ZErKbi6ODEzdTt4bE
eC3vGmfmDMkU+49NaQNyN+mfQwLEny3kYAzLmbgOj/TZLx9TlLTM3CvZ6hByyXG/mmvbjZGAnYwl
0PKeJr+yn65M8VS0Injc7vg11hkztoKCzsX+O6lcFxl45oWxhG4DBRMGtf3ukU5iaNVkXNhSMz6X
sAt/1uFA3PhpNf0RUNq0k3WnKy21y35i4eF1aIgqZmFzr9vO89p8YNWk4waalKEMzdhznF31fAEx
rAxWoQ3PWW9v+stcWoeR34CFKPVKFHIKOPY80fdlCEbmAC4Uo52KcBY3Pa8Yxp7Ok6vYxqTHX4NT
vqoAbHzN6MMTemXxezlxfOldjhnuPgcKjKEtcdId37H0T02aghLNlwH9SNN01S81nWcRa3mPj+2Q
fmcI7dgby03BPZCf5eC51585U+2dJxuIsLn3e4qHCUzoEFQ9C55RLccIqbiPSlIguRJMl1Vpt4Hl
xV2Y+f2mAvpPo6AN1ZVvV/1h6srZTfv+P/kMQRUCOn52pvqmKhNGaQ7LTIyCVcoukWoZeVsS8yow
1WxNAKPsa81xJUIWRhoC3nh+PpCchfS3+d+Svt/7/BpkXP+1hd8HXpOgTXTAh7M6j0c9C4Vkf8Rz
GhhKn7gARcgF1ZHCrtnDAKwvfdJJpubIE+2C9UXQei4MpPx+neCPplxPfhGSwwrPR+fOzfh7LIfV
mGzMgFNgKM9pBDDUEzyU+f2y9lUj1K0KUw8n9mqSFCfEipVs6E9NFJcORWWWAERvKJDPB+uPLEwU
ToymquQ8OOPMpvrqaBycJg0s0GiHYIlvBVUezOpGwzW5ilJDMItXO498pgTQHGzHU3S9RYOhr2Gs
WJVp2i00Cvqxotz65IdSR7Dv9iHepVKGuMCUP4QIAd0Tte/JU/zC5lajoNWeIpT5hCtxUKfK+BtR
x5UqRlArcitQU7AsDPlNCEdp9wMTmrc9xxKVG++XYd5JA+KLDo41iw9hL7TBM2Wrec4kitqGZ4To
L1EKXe1pVSRqAvbwA5WP1IOwtjbn3P80dQce+jqMT+7bAr/eYMZovMPBKVFUmBRN7kPVoM3HsqMn
phma7C5BcQSnVA1Geag7IVrhHf6brCPPtt7FxM5ATgV75LMkGMQ9Y+rsTDlNkoL8UMOIGIOn5Kmo
H0yZn9irN53okfXGAjySvrnLFIfqgUAFnrXYaq/Hf/IoAeoszTTld/T9no16p2/gzlrw+YfabN89
ewlooa4G79bWxjVWRgvmsu1gMYyfFRKoXDXsUtEKFm8AmV7Wnomz+FqxOM8CIEvDGKejCUkdmY2P
euybRcQa3/uDqPx76SU6zM/4chlH+Gsb0sEaXpfFe5lP9w7JsbcvTj2WEm/hZ9GvPsRC3beT79RE
5l8c6SuosP0A9oqpMOFSXPqQMrUlKyYNArqY2r29M+wUNgBZ0a8SQPW8E5JYbE5QOWfHlVWtlzwc
v97QSIARtGuoVWBnCqTV95cLuAn4QDhOeAho2cRokdtMNQdi7kzZDakDLa3O2/SInCQimurLL4gy
gISwOaDDQUtGhuPYsAfweKPMMEESKf2pEjNrdfsfstb6BRNizOcH2fKoFzEVmRh4CkWVTSwREuSH
Tmp2HXwNQXzgf3TgzOKnrO1Tu2ewJRU0L6vub7NNLyp1n99SWbiFxtN9lcyxLyIIAkVK1efFzfb4
tjRRN5YFxKLKCxqJbq4yiInzJP9oxh5MGNQ/eMLoWHbyjvDcQOsXZkjQPPFFMOMmJwBPU/8aMG8w
yxz+UP6W/lQRMrctuAEXCQMOs9BclQfjuNLu9Qui3a7zybgfKWbOCgo4f/euzXKtfht2lGnn+fP5
E5hTmgSY7Ui7AMmZjIfNlk+l4sTTl/cE3Y2I8ptZ28wMshl+ENgoxF3i8NdlyId99HkJB8Xi/9Io
xs77D6ZNK+cBtzOlHD2S0l7JD7PgP6Kn/mUXKn6Q2Va2FvOnVyLX0RT9ibNOofbiSDnuEQZIeELI
NI6NezQl+iRphzGK6wH9zWN6C3+RsgmCQS3DE9YSn4Tp87J+WvSK4UJV7YMRbdOg9dGRcHLJcpIw
Y+kzpRuSr4DFKV2EltvtkULd8/LzH07kGJDtN3k9Q7lF7uk0KJ8pYubtqY5DWyvHlJ6IvpQ2mTSy
CPnxK/4ZQdtqzG35W9vWh4pq36iCQaVGPmcROqo+ZHRJNyoqHW/p8BVobAv8ZQDg5ylZLeLUkR1b
micsnex8/sQo2QUVKoZvTmVJlT6iZZHItND8fPbwMCglZ34N/ZtWOqr0YSNQimUtAmSqPqb/bgb/
iy9DaTElXsTEpZFTmFOtppyynsPZwmGRqUTkTuSdJX+RuCDO+NaB5xfPiiEJNBPwFFXKoeTW8KWR
C0KfTP2E7xPfhn29UFLynzuMpLuTpmSejY0eOoSCIDvYBPyZKJwVTpbqK8whxzal3l3A9lZwvPcH
Zm/Jpr3dX4sd9SO2OclkgTFrJ7lpSCAgHwbPiQC4WPHITjRp4aHeDw1uDQ15D96i2Zh3Shy/4TXd
rcLShfudQSbGtq/DV5CnsT9A1wmCWD6xpyGZWT1zHPurgx34yaqNiNGu5uLFbX0H0E1R1j6W/kjM
Qyr0wPY1VDd7YiFL91nkjPLaGE5j6fgCDhlAQwNC+s3hqpF7SA4SNZmzGMAgx9Xg64HndLq0+8UK
Q9fXu8+HPwyOEzcW6ffFZSftEy6qG+3qSloluk2A3GU74zgJ1FZR2ELP/Rj5cK65ow0ekNY/pIlC
6uKyYnv5lpeR9mlQoFeshv2qwzoQS0McOEaAUYUBMtLQc7+3dQSFR8LoZSKqTGi3X2bftjA7Dom0
5ap3bZ3EQYqSjiZxbKG4xWXo0daQCqNXUqQbR2ZMb1rxLoUNrt9r+2gfV0YnPcJ4/VcyRXZUpkFq
lz7A+5aHR9c9sc2HN6CyTRDqzBZ5MlcJ4PO4x2AGSDDi9s0df4BGZ4ddvoszTF38nqUShuTdrqEn
IWeqSnqynkQFByLhsYXwTqozIOIT2Z8Rmtqge2TQGwJZPut1IJWvdPU/VPaNv6SzSFSCL2Mq4Hyk
4SLDPNPw0zD7IErTA60klfbiyfAfpTfyXUKCnqMX8Ad50aPwbi0wUCkLmjtMsXnjqROGts1GsYv/
Jh/hPEfOCzDZHDqXKmZAGoX+m3f3ys6KZSELTuimEykXQEPrbrKA+2sCWx2s75X2+Y+gi2B05OeN
lqKiO7d/bksgvvAWTVjssI2FE0nQtBJYxocBVhjh0+nL5dQm6ue7tAwkxuUWcBdNTjVgKJYerPPe
uPDFCz0KvSocTD/eM5sXQJRFhjj/0aaR+YcXihgBKG/411eliRruWjpgIDcGzEJae8YEAcGtYV20
ENHtWpIeeAoYLVKhvSW4Hrz49/6T6teXIeBPtNwQ47mWItUp6mf3BFklMNtZJ2QpbMeVjzgCqKMO
VxK9kI9R8DEjVnbx6Tg3U+ZUWbGuoeH/yY35hAbVHRwJvzTqD+cPyY7QuGD0GAyK4v8mWoGR9VL/
FMYQXixccnATxL7zqhWvXppeSzMAWqmkt9he8sx3JfuyC/E9gUY3drPvy7ivPLVlk9Orz8uVYiOH
Jr5p1WI71Ic9wdY1NOuyOtuzgRcHWP/sw8L1mXPs4sle33S7T/b562FiCMuiY9bizSO8W26ZHUpo
ht61RXQgNraSYF/cbCIAWtXmsClsP7HkXp5MziKbJRDDur1EaH3RMhs4i+MTh5Oun0dA/iJYkfv+
l6NgAvXVI/D39bhTJw3x7sRw6LgYZGEuSWxj1mspsIwp4gxJy+bjrc2JgxObjfs2Drv/W8xzhvt0
1M44bZG042u21huwoQxzXNOPC/7cq9bwcXZBE+x8mINvv3sNpqwFY+i+nXf1TKN/pZqO2xEkyBnQ
aw1d+91WACJ+ZFKGFkUT8sEGgPAsXb12DW2pwuRhnKfkgxB3xih6TFkgRqKphIjE8DvMjPftp49n
AivwzI/gTy7TqE5yqC7wN3PW3WeS0v9A9CbPAQKv1bNeD0sH5KbxaYAaaEVp02vWOjVLNi8TIkT0
vIVz37GlE1pFHehLO++qdQkGJuAYd9MUiA5uY6QSS+U2Xs3Asq2ulehfRDbSpIUsig7v02tBCukc
E00s6yD3JGYE8JC+Aw9y2gEeAfg5mCfYdmkUE8rXY3oSECVRS+UIAE2c6DogfysC/PNJ5NIQUKqM
AMeoPYjxIPxP6sO4uFkOlRMjwWPqr1ZdZFtm2/KRoR8KkAIOwvgsK8CyYiUOMyEj3CRS4Hkq1a4P
yHP4lj8FlI7xFOSRkcDgLxtWbrqL4oply8Lt1D4FedRMLa+ygFWfogxaLEnNrnwjNJJ5/p6eHJf4
QuvOMVcUIsRdghWRcJio59bXDBlGAkIGgVXRXlfrX/oUuHduQs3QUcfHQ9cLnvTJVP73uLNJlJZ5
gZjlm42+kyfBIN2qtC7/H2npxQ1+RZv+MSNIvfX0RrZkQ/hj8dOFaueLPtEo/4ajxN6tpTP7uOua
iKIYJzNCF4gPFrCD1iHtjlLIVWjipzvOB0gqxnuzmdkMOzOtiyke9LK97aRgCD6xu29MoJPA5bx/
qJr6M648uRXqtEa8VXEcPUv3XzCcLNxpuIrR8JdmnyhRjhmTz1mfG3y+dQF4k2NB7m5F7ldTJLSk
+r4nROOBEvAmbTlMLHdjkbKoLsSQr2U2O13XOvTfWdg9mt4txmAGj2WIlsg8tS6SvB1jUCnBPbYc
LTtMvMrXa5enGNhSS7xfGn9XrHm5T8qvEz1nLmzq51vZk7L0w7ElFl6duOPP8VW7ZW2rTxbcMpam
Winqz5V1TcDlkoProWtqucYw9+34OT3o5dVaTZOze1+MgEQBLENTRH/njfQ10KlZ/k6XpOu6xQmU
VmLUTwiq6T4ABHNN/8RzOabsY3dcpHBh3Z0G+WdY2yxtEsGhzejP3JQu6MWVuwscMYhKM2TKmfs8
KrQ3RweUnetv67wauHUAX1FagWCLnJD3r2N1FhJ6jy+gWy6O9xDrH/CYBpvr/HXWm2Rl+4Jnso+2
4Y387okvWrH55ssXXW4n4maCEwM3lnz83gbzuqymln1Amq0mIuLkCySZLIE12gAZoOTjeDe3oC5/
l32e/pDb0ctiTeVgLp9fm8XBd3/7AsZCGeREBQRgmqoCGTGZAzdqfF5wjC4APkXT6pJsJ9QvMDSe
2gwAjE0sDjyfA5BuiKBcQDSAa8gzhMnanZdLSd01I4n39KyLmzU478KJYJrYhgLa4sB9Ao284yqY
6IFzbAWe1pBwc/vjBWNpXmNAlta688Nz4/q7FQRDDotnHjhPvckSThK7YI+bHXuz211vUwMmNB6u
cglxVUbtrQ+yR864A8eBdPy2ayfBkr7y+qmo5t8m8gVOIlfafXYulVJZ2EJNhA6pYcyrVQKHn62w
TVnDcVn7eC4p/3Upa/fSjS084dd0cSOJoUUfWGu6rkXPohCC7rMTuX/wDipnN7xjHmuNCLJ45itJ
olU8laR0ROVgCcuGuRMADjj/jC/XlaURubVt8u2RSxjwGGUFvWzySOIATfRd9ZnQ5QjAkao+H+lF
Xa91vo8dUBhPoYsU1oZGtf4obWNYHD2KiuwbFlROkseI8CL5OzeOQk0b4asZ0LwA6aVo228mHlpn
aeK/DdH9wdPrTOXMuAbL1b1NdPvIO3DlpDmPcSrLCjVsCAMuAxwA6K6w8pJaY0HS+BFWL9rFl92t
iG8BOi9LymUf1/PspA3onSlFkrAS/eKT9Qq2XLF1kI/HFJUPpDY8NYLd45a7XA+ZrgMXSP/60cYB
+Kp+5R2d4uyXjBtJRXRsMdb1LMXAznfGzC2dIRIkQ+15+3X/2r/zAjQaXP7b4xmWdWQQvQSJ5Myy
+oLE+PEBUXnfIUcRGv4mM0FgsNTkZC2PQpc9CzVIS9cMr2ocSxse6qLIbbBwxNoB1htLZrcmAmne
JXVcpdtzd+NPBFHPQOOvtD+Y11qG9Q/doouxKl6mubyheUEoFDMpKvUul14fWEbffgu5PxXBSi9w
lo65CxggQBjgb7GSpO7+wDLKQiT36veHLpsLAesJ1T6ICV0TYgz+273on87fQ34bcrHmcglykup7
rfEAF1xmcPRbXJbqKBxvBPa0yhvWaREwJq+grxMnmNEMFfA2kYwQH3QH3KvkSdagHyn2S9axlAxH
diaiRCvu0HRydpTfeYorhScTFMBCpHOBMcG8gKs/q9ywuwqdsyo8ycXzQUU8YxQg/qPpeaHMvycM
cvPnC6zs4MP2bo/xPjfSmQxCQrWFbfE41vy22zG5c5N9tU0JBY3Z6HLLDeHspXyXdk/mkvpvSFjj
e5X0OViGLlJWL+BNDEdCLMsx6m7jfM06nb+xkjXOxCE58D+tFpAZcqoqu/3dY3sDLe66W6lecVYc
Cxw0zO9ObCGMY3jk1LsPqCdN9sgxyJcolciwdaiB+WVQGxjQs41wV/A/vcCURBAiSdH8Fw/31jWe
xbG5wvq62CcFN3fffM60F8j6icH/gnHB77HrnnYkeN9QNzs+DAHl2jud2e93c7z6n12A6yel6+mn
SQARev+OYmCyCfogxcOT8fN0R3Fi+4rKtNxNsj2e1yyuug4Hk5qjZBijydNjjnIQwBBa5EsuEqka
MnqXfEc4NnB1Aok+OEfVflDrkqqmhL1XKXhWdrfFALuxUvqwvrppnHaoD88KTLLUtJECdNnRQ536
cOkN3ENrFpUXpcRPnct5Lm/YX8jFSUjLd+vZtYa3DJIp2CFOvBITe+qbhyHlEcTyKK0fIiV/YqdE
WtHi0CIrr5xx+MU5UpObSJ6kkrIPdVUqsakJMM1tjllMtBBnjtc9YoO80fJ1eOPv+jY5BER1zFnV
mhC8ArRmUKezNtMjWc1vXl87E9pBfbLJzCggDhh90Zkl84h29OnbtzQM+MQdKWt6LJEhQ5VQZyq6
u62tt8+IwtqygB+2aQMPZ4oK8LQdTanC/q691d+ySgOCzgLHnhOJ52zdyRFnMPRnd53IDwFeyRkr
nhG5BkiEQMgbKgwZwtQ8tBtlsYgjaIvNI4PIoSr0QL7lOT06/co8Jts+f4z++wr9YNXRnCfabWWa
OM0UA7ojUW7phoTURbfjWUYZFV2NdbEXeJIgZr0PhJIStLMOhVFRgKUzvptvIsEQXKIMDVyEoHW1
7XzlWs4WTJWs/atDUM00tZPAvJ5ocUnbO1mvvQW7waAml1+u2WEvCHbosIV8F7VA9/qbJRoPjl6S
L+JnbKwavWM8iuoNZcu9p0BYN5wkA20XIHbAMCA0EAASDD3oqTlSqXTkJs/tsSopYpZ3v/oCulL7
w++9YM3s8P62T2Map14yLIQr7YakpRIi0nX6cMCYOlKUXL7K+Rjh8EHw4kVyB2VdLTrhIKdsM+BP
zhuCj9Lcs61K/PfuD2x0qtmg4FOodRsedA3QVQ/IjommwkCIazAOGd1qsG40WRfNarV/AbNmKB+F
Z2Cz1Md2bRxOwhzX6Ak2MZKFMk5iDA/PfPdMP2wi1fzYyOs5BdNhxu+GmuD2wISTziuSFmGFu7u6
NrISfLC9brEqM/h+YoZgm5ALTgMz4h86SRSQhfYeBz2TqGFaBFK/1VK2hgJI6X6ZAov0x4zhJM/L
ecGK1mY6GwDOB7hehd8tzjJOFPAnKGLMe7En7u3mhdVhebXxOsBS0HmeZ+oCpHYYYHTckDI6OnXd
r5Dtbb9hKroFxplWmR8lFQgoS3rJ4ymPcPM+g5DwzB5fD/4IUv+GFkFHKbusPQZcS2PKpW8Rr7Ne
FLtzH4uOecpr3WBFdfnIckYoZxWHK/dPhsD66LftT9DFj/P/o1b22IamJxD0bysKEKO+sCczviyL
jxd1uvgb5KZsoQ7CZBX8qFyT1lRzoSP/Y2bFJFQi2gqIQxQOi3qeJbdoH5X+VuaKUgJcNcKp7T6s
DyLlz862PLviZ/tOzjb8fSVRMsA6JcUfGCPi4FxMEV3dvG3VHGzBm3icDImSe1CJkrZssRoMHinm
pvg5dEP7/0GEsks7nrZYh2j1H9vAV7ILEUmZPu2LDiJIrtfmai139z8JX1vvrpUuTCX3aag1gsAT
W4m/M2I2/f21uEiOq9Yl51cMRIz/w3VrNB/3GgX5JIfipDWPN5aW51diIf4tPreRZBL3aM20MJ3u
P0J6d7h7iEVlOBxusbGiV9njWHB0oEUH8Ss2wHqzlcvYu9aKFUinCW4eqeMS2++MkxFcgOXhdFMc
0rbU8BZrFD4S5e7RMCWMxz4w7AyAatZFx9iqS8i89dZXOEP1TWI+/0b+9PpMrsh2kp3KRyDCOwwd
Z/LH9ebwa00CBfEpun7sgluvEtULAKQxgByFxcsLspalOLkXn4XJb8TchVZFc9fUcjZkBC1knzze
4Xgt2/jcdAcuAX3h/C9H2Bq4O6o6XAPMdEcIQiO83aXpMjHQ/05YirWS1+kq8evCycH3KjSBH6J7
vCH3aSwIgA8ymxRO50X944+qNSUXsI0Sv43nDXc5NAcPQCh4jlyqv7WFzfdH/p+KefbMCGU16pJH
J1SAmBeAud7gz9uKc0KIEpWwIbzuG7aGJr7idrxZR53RxkmP50IILIH4S5paibu6Qcp87iAMtDS9
NWWKsumBmolLBRRcsTfkPRTQj4J3+AAjQqLjL1vRWyCg6hXHakavmkDLU52rFaL5TLd02XJcD4v9
kjFm6LFpulgmk4MxrFFRvDipsUHxcwS7uQzABfDqzowkmrNLN2C744RJ/Rz7JdboY6qk/ed19fYx
dqqhyYyIhgX3e9k+8+WUT/GFSMdSk+KLUKiSjKL9KSEsIbWtgBZgBnMQwZd10Ft1yiObQG8HJggw
NhXB1kQ+DJQSxwGYSTvqH/3zOxcFt8lSJOrMBc5q8UL9FdV1z7itKnW685UV6xea8xADWRF7lCfl
qWrnCgrKGWF+KSJkPRve7kiymVz1aKkR5/DG9FiBAl1m+7C+7uCJnK10REtwgg41L6dzbHPz9x0L
zcqK65IdtHEx1GanaPh8EFISnQXhzvIGb/zObxb+wyYsFmGoMRN6MctgtpE3uxDZ4daHTpNAmCbj
TUN+dW+lmD5M7C+98CxY/3nSKBnoTrQZkKkrDK8tgGQl5FBM8E6GeJXJu2yvci5k+9lvtYYa6j08
rd25znfZ9djgcQgUj5knSq/vF07rIP5PU9hoV9pvvkyPQXvEAxdiI9YWnGchBIscjNF9T/Ad/Cn1
7pLJm5owy1xvzlxqepbG9lBeRnKrwVhSPmM2bGE5PjtbRzJp4xUaF9fJQvb/cn68ajyqpiXydgZ8
OG76xqO5/higRQDBolmCW9M+cbJBx21qgAs/TVBoHTFk4KvLdiDqhEsdf6fb8zoPDcXOYkHM3dqy
rX5LSSnDNTDmkOJ+GMVdYZUe5LqQjBA7PbtW+d76GF2xr+7PeoyQ4jRTYpyv9M3FEoNJk0POy5zC
BAnzP1kjauhwE2oiD7MQDWUyHbJOZTr7TJLyDcLYO0ms4axqWJG1f4FbqfSMf4KD/4yf594IKtxs
P//1Pochz8z4W0xTYuR63x3jgXEveCmHQk2fCER4zJOQZLTnxgYxV6+ypeOv2CLup5lKVlreJNrP
A2R0Y8yCzf6day80GDt3tAqLaR2CU9fh1Bx3HMlUFShu0NvArAr2AjEdN4eiML56K07ZU0PWdum8
6QrIiPYToqJ5qu99/9ppWqi18fZ/2No57P6fQ/Dp180Kti0NoXKlU5UjOTkr+T73S0hEcWz8yuUF
UDJFhXp5OnZDrXUtcESNZdFdCGV5rVYkfuonvvJUM6/C8VvfUZ4nOgDE6e72pfdNnq7L++VbZV6q
R68lh/E8y2az86QURlxi48yiy6wOCcfzRwICbjekDTdjCTBJQqX5XM96cSEyCxX+VmHSRzTQiY2C
DFLjGbz0Fk9vexDNsJ9klYskjpLB9MUj0vKkJTRn00vl6wcEcV20qXMIr+z5GvlMkjjHyj3com8+
CZyCXPK35KTdDwDkm2dM2dsgwqWaHIpVNQbqgiOgO2VBltMdBjLdsJN2/5SxLDp3xxipOklsSQF8
R/UP2AGgxCNaXrVtYJD5RqXGTroGOg1C31dRobKpOoTRLEhYMxbk7uUuG4pweY0SsmNWhlOT3JMh
XiGQVmnVEYroNlaTHyagm6iTX2hdfbYFMWjWco2BEjMQo4cphr8nKUO0VFDo2nOJQNSGoJprxwvm
fWc9azPwF6cLXMsUkwOMmHqDL4cWS1m9122XAd0TPRATv4W+jNVfRAAUmTklb0v2R8f5sd+QxQzo
zlfRjZ4sU/eZs5vlCG43CPWsLgsHNvCPiUChF11iJq8bLQShJjQZcQKGpTfJtHypIwt9gAwVqt0L
0Hmf3j8VqNAY0NGJKddBYq1igNFdPnGWjwHGIuE7tVVkHlA6BxwmTVPA2BZRfjswWjT1uel3HdWv
SFe4n6uud9eub+Gk3hT+NWchKNGsFOpB2wNRKbqnbzen3kkMEWKocqID/8NohRUWmnynnsIab+oZ
9X+wY/s7g8rZ4cqy7TvhGYQmwlxajywMW2FUeQthZnQ/Pt+xoQ7fAZFhZc3X0Hu7C+IITcFlSYGi
DXsktZi48idK9dH84LZx4zCwhI6pl76bigJ7esi8yJt2QkUj9GG+92ZeLmhjyZQr+sLhfkt7kZII
dy04OnY73quKr13dKfZj5ZJ7HprBpSEnmKQl/zc1BJAXqcGiX7SwwHZCSnW38Q+Z1XvipVRl2Ro7
b33aXXXi0QZ7puAP+lH80iw68TgStDvnnvNn+dQy2Bwz4Vd7PIEChWvHzGPz+oJ8fnaPOuQKiuS9
+cf8G69uOp8ZNxzy58kanAeYq6Nh99Hnyv23HPwnb2QoQXEmR3SirqEQviZPOBElzQdI1LCmAsGo
RP+J2zP2wNbA/tX16WAvgZDbU9Fe4vizhzaBnhKssGT5LHrlilG9TzHlhzruss0JAFNEWv3/qckX
15XKBVs0bnmZaEwFtemo7SiTD+05WoPlipIQAkPGOBwY5QIIdh+63PWMdXK4liG8QSruamGL0cNp
9AZMiK68b2nk5UGNfGnjwg6mnOIwSHL32WWoUOGp7qAFoQO6PhpVbyqCvgb90cbK0rWab9B9oFmt
uf4DKtghZjMHCnithfjviskhFIr3UExtwKN5VpOG4+ljcaz3ydCIQaN/hlhtm27/waYeF4AoWbpP
+g/5afXYSPq8geBfNKVeOxsBVrULcql7I4kVNtklMU/KUQUhAiX7KT1m2cVCoIuPb8FPZAGQTIGf
qM/9TRZj394Igq7jzmQtlNwtKiN4lD2g8/lVRiEX36HD02ovdNy1vSPVpKWKx+6JX7226zef5ZnR
oT3sNOGy3E8yU9jmFlSFmCMnYU9rlOmLIcuJfYnIkQ05dr8Ry09QvTdJUknbtOpAXTBhOEhS1iWw
z0J33UtZabG85vtP0Rcms1Jwx7bVTsGt1Wl03Q9+DR6mH77vnSkYF5XWSsmiZzYVsMInELQREckz
EL6U/rcupcxQozgdgIfH8l1yaCSn9ZT+yA4txz1SDbTmGID4p+VyF+5G12/ARWr/tL824JgsUuHM
lCXow7O9/qsBO+r/cZSLYYaGyQEPcNGgROx/t2Y+zPZeABNBA2ESj7gfTyXJL54wPAX4JhmJB1fi
b+chi7MIkAzgX4kL7pveSUelddHOUotZBWMXCCvuynzLjItGSVD3qhACVg8Arm6CYweaXBJvoyHl
ACX3Lk1DmH2BE1lSOZWBVvTQmt8Ds4PrWAoBb6IW4DJmrXtmA4FqP8lVdKxsBQkyfimGeUEBR0mP
t3xNeCDU5TtiXIPNmezIAyv0i1lIMqralF86ArZ2bf62lh4AATE94Xkd0pbj4iYERitB8tGeUaoI
64nBfRvSepQdkZg/vXZWWVYcp4lPaHk3ttF2KskDzu9rP3LHUgksMJZmD7uFnztGRJwQwaR56m20
OmB75WosFE88AhvOvqAAa6aNtld1Q09ey7TCnKFxcev2mQsoFYZiIayqhFdZmo74krY/SO7fpXuS
HNcONZnM6hNnvNrtt7LMS/8n4g5Rkqbi31HAxCzZCnssCgVU6hvGzjfb3H8nRBSQTfAXuuInVliW
kDPsCd3d80E2QZGuQIBZNJQbmzlKWOtx9Fsqn1msWI27uR2+YkT+6YzH3LSoPW/vDru5B6MEXbq0
RSmn87yCBNwslccz765Fvk93goFEoT1qC/lNG0LZm1jQLu/DGWu1OnseUSi7IKDXiAcY+TlHE43t
uIo0BfKe+hujYAcImCGk1ksSPZ9z6ubAU6XNDtHtPJ/+SPXeVaZV1MHyTA7AkwFzXs6wc2Rdt0fm
/SskgzQ1/985Ju/kJGL3R+MKRKwpTBDcMgHPOLzvn1V/rZKror8WO9EADd67fPgJPTK6ZKoZKEsn
UYhT1Ejh5BTHhSY1LNBud636byeULgvBVqytmGaTbTjfH/e+orZgmtpXPohHUclWsmBnuWtV6ilU
/Y5655sm9biZQ2gJkgNOQwjzD3kbAul99IuULhfuV1XChtn7FsaSbSDug0imAqpN+iQ7emdRKu2q
c5TrCgjTaZuCAjmCFE5H6+jNWOPMUfhP9NJnaL2jEfZS4pC9x5gfjcBe0uhGRYMGbo3wAaCCz8t6
ygwY6fbUL0Zc5GTskA6+MJwu+H7BVieIL0GmtEK/SyfSH81DlUB20rYZFtHHynpiLdIhADwRwHZj
YuQ0k/n89r2M/P5DZLTyB18knJYbv6EcmMJR2DzHFIiLSclUv6CKVkKx99eXWzeV6x+SYhMr4+qM
mvv6len2MPzx8T0rlF7xQnXU2PKb62iBbRTYMbnbj/7YGu8d+AYAbbrqBDYJexB1kDyaITqehpE4
4pBlUSytrx0tOw8JnhrNlddXMdHnxgFEZS+gPIyVdBdRSSCC1oFAwyQ1/R62YhPzWtSzN01K8uvc
0wEaihDhAyUzOjip8QJXKzKER2A6GacovlKN5XgVbteHynyByAI1ZMRQn4KNjPltSLTlO8zHmAkk
aC6UZhFJIFUIFMOCRB+39mX2ysOeQn94XENwjPRGNqBdUh/AvW/O/NNX2Lf6z3w+XUVfTwf3E7mB
3hb3F04hkhN3aLuX0lXaGDnfonLRKRkO4FgODEkkz4J0/Z03T1DPQraFu0Qz+iPpgOg//U9JcbVc
F0Ktw6CMrMXFYDbxJZORnAMg2KGo2+7b5G7i+yTwoD4EOxZ7sX2O0PFab6Ga9tb97ENr5pKr5Tqq
3N/ksGCzKjMUIVjccvsMoSDhyatgpgXLWh4CVo6i3mE2qEkiO7MoPOOlDk5c5/M/0qgVK0uRDrg7
rUdpU3wV3rwGpl4Q2HlOACZQp+4uXKlUFYk5wSd0PUWCHhmQOXBxTy3kzJz6W6uDUIyunBl6/zqS
N1GvRep0oak3UjejA5XcsffaejYvkrR8cci47YsvUq7DSSDwzaYlJ8QiInL4ncfHqYX8AhvoW8BQ
zTYjEX6eIAYsVgpyMIAsPOA+52QcgZAKYsmzGgxNVlBIvvZ4LXKU7v3mXUhsUbW+mGFYGsywVgPx
Zoy2mhX1KQUkplzYKLK++6ojjcnqPHKQuWt22Jqqx3G99TDgXBUC5+AW2ANWf4uMHQhfJOFKnQcl
oYquDMxlNPtN2HZZCBQTCs68Qjrt5YmM6ffjH8AoTZLco2ujSL99AuWXMWASFhGybqCTivvGEyaC
fFsEXDLIhsmuu2f73daBqp4BSYpN1Zcq2rQlQGxPRxJfSt3+OK4eWNTb/MT/dnDDbQDGxDPH/Cic
Km24gAN5uvuIe1ZRM2Ng2+j60qL/ExCjjnneSNqj0Q4nQyD2dMRzhqKjTLS0G14V84hNG+spFAnw
lLu9iV7HmFPXlaauAseO0BAP3NiWwd6VGH/+LRO0vzci5uPDVh9j2ChOIbUJx1R0PA2Y/z3TC93c
lCw1o/yUKNiu+E+zD/09Y58HcK61cBApxy9auW8qqWWXUVhUm0VDI+6sy8JET5xH5Q80bzGpW66d
t4QkQTDP5ao9MZGqaGVhbWfD5mBvqDuTm5Hef6wmJ57fJM2jbEFe9rbOCp/QxiVX0H9IKhrOQ468
aLH1WXNnpWKFprKkhDz4b89NYc6rgz4g8PJgY4V1U5jnw8Ofxx2OMqBWP990ki70hV0ueHxaGnk/
KrIVmsECVfhLknC3PGDSFxAodRoSIa83HBRteBE3VWu5mqdtn1ax6U0vNhjsJ/mNZbZQVb+m3H4I
ScAtzj+WgJtaCoGG9iuEK8e4vLQIwkLtbq81FOA+f5wuIFu1qmD1ho6FpNt5AUi8cjCkQfSNZjOL
fUl7zIX4ZGqkwNaQ5qqGRTUxocr9xJthXzAJGnG2M/7zoqPFKOTesJqhOAvA7IiIjckAyTtMI+wf
qKdSUZqAjcqTiRTeLGEy3C3uhnHyO46r3qC1rngObdQhgQRCzF9+7s2DRf0SnnLkoex6FXROKRiE
fMQ5kSbsCwl6wetEclTCd7auZEjmWfAm9YRBPQy99niprwR5U1KUhksregAEptGaqmfTKoBpATny
FeyQvx1GVeWZtqumZSZspQud7fJRcLb5et1JV4YpVuAGo4sY4Q1B0h6yTJlRXqgeUhX+ovueoXuE
wsNQyJ11DOqAi5kD3xuYxhhs2EAhze+ZxFXnyt1+mcZioDL+rIL7tSQg+iYlcdMaVcDPADvk4wof
tHEQdtpeWNkClI/eHGGDdbJipVdz0r9ubg6RdYjhMlqjdzHqavsoQlbfo7T3PLWe8Pugm0MbsvVT
egtzxznxUr3Tx6Pq8cysMMIXz0tgunBV25IctZwrGeRtNk44mbBm/Aj3K+JTOoVoiqciPlp4efY1
giZPgppCy1tS82FDyQv+95gqxc+NBI1WvZTRShlXgg5jLpnfsRe38f4yt83V7R0vmF71sQ0IDrU/
FgliQ9l5o2iETbfoOHh6zJT70QW7cu6NbOLHZspxiTdWrxTXw28fN248c8OUXGlHL0g4iJUeD7Z9
FLLBqL8c5UMEliqt6mhVQm3+WiMV8bx7N+EHAhl/A3GA1+gJxkQwBqEZFtDrv2sZiecsFDu3YqBQ
Z+eVVYGLt7AamN1ggKOIezZhenQBO/C5H5MJcYGo6ybBLfisQLu8Uj2D02o6TjcqCb2O4HXgjFxi
SnBL7D3sV3v1YFBYjMjapAtNp2s34s6hEECFuKy1XoryYHvKaYWLlljS9UX9/FslsWD7Ulb0lLtX
tOJO1f1DL411Sq1sNNotgt3oTBz0kyGKKOen0opEux+jMk6FVb7GXLtKuYD3qN+gdu5T4xm9L2C0
Of+cgXaupsA2fj5+4C4++DxOTizQGOPHXi2CRx308EwJapvmrcLAZ4lz+9tULk8YwL+6F6V0W99P
lbNEOE3+zQPFpMVl6Tvnsg1ri3/xg++diER4saOHmfYk6HdRfv3Rn81aUn2xmd/CF3rfAf4pC09r
nmCXsLg5YCVp8mEVj8HAb/DmAzqzoGcIBFh18ZAakh0NsOVOeMRqBd46gWheqYz2q5r0TrGNeVGV
sBE6KXU1cCEKWcONv5tnncBpe2IY76XWTXU/e4MkerdA5FGS9Indfii1Iq2hODH0H0JA7huErjBv
Krzt561FIEoZ3JQb3yEVKjzAbOXf0R+UsmYWKxb5VNbN8Xe7PK1PsZbDM04/ndImGIVBcCauZVmd
0c1b+V9QhK0OuEPqQNUwhrsfZygLsa2BJNUU11GIveA5ZXw/D45BFlXSJl/AAO2PXXRBERNjipOR
aNCpGrbpiT5JwY/QAFfmKaa5j8Hcz+hgkSYrlx8ewuBE0xIQLCpz2cU6c5Rt1Jb0nmI92oik+bnh
SmVprycn12KMsoYJ96WwwC20r1WbBU6UZRB6pmSDt1LA3AupTtYJz+j5uZdRKwclUE4NcT8Jdl8/
Pw140U07enNtZziIvNprbhuPF2JB1cTloxX2E+qDpdzitDAYnViA3D/kYNLPvdQMYyTzHM1rD1z6
tb9jXO8k123koNw04nbykTcpMSJuEufVAu361NCwpiIxW1qdrZWGSgCcJmnYX8ACxxcB5xKSqeS3
lOfy6/OqiqQJKheNZC5aCM1zGI8LiiwLK+LPf1hF+f0iQtD4hYhh1jbPMss5yFPZWCGB+b3h42hz
sivqra3HdazNGpWtmco+CFauSua926TMteOQ7jsLMb5szOgqB2/kyFru13+h9FZP5hKfOUi2i6/w
EFGq3yULLaok3MxcEiY4chTTNnmEH32LQ1RFqT0nC/HpYwU2jaDpphzk5ZsCxxkaFFrcjOrsqc37
IVX4OHRds1sfPdpUGq90ZYk++gRO3T4WCc1iUfdcbY2xfxDqtjCg614ChcLs8f+EYn6ei+VXAzFA
cI5DGhl3embXfkEj69txsrKWXPN8wmYf7wUoklnXotJRpj7vtnKMgPR4wDhSHkAX8p+XBcqQtELq
LgM9fZJTYnMPnUurht6aWsMmamIDQHIRh2M/HQtWRU/W6dGVql6/KfU6cAFRjqdPpM368YG9w1Nv
51lfUu+cEhxoYvi2gBvyELTtrlRJY+PwNbbG/uXb4njiQ+FP6H0NaAvkZDizA3robWgGcotpwveH
oR4Gvq7WcM5elMj7bTWTKru4OcdQTw5u/Bq17ZjCiISI6JqLzXvCKruwx3SxbuhNINE2CO4W1sAh
Qc4UoZLTHo+2nJcwunMx9QTg65S8DzpnhdVW6aX320ZmXZFGNMroHkabInxDddiUpY5qDvvijIRe
Is7pjV9psVjzwvj8z7fCM8Ee7ddr5+wzcwNznBEqVXK3NR814Y5Ff7BnHt4aWQYMF3SCQklXqb0G
ZP8p2gx2jFf3SBlg/8xC6g6w1iKKn82olBoQDvq2lr2UxCY1SwCsCNWyqahAWrJ11y2fjSWt65Q7
qPavjKUCm/sQ26iTuwV9SEhjOawvaWQe3Tj9jFYIHXfLsWhs+qeUH/kw0pR6gwFp4d6GdBUrr+5l
hV9Qz5l38+TbhgWS5+ikoeRTF3e6b3iEsiE4tndY43vwFCjzWjaRDW9r2iaXZHqjNz62yC4Pzejl
bDC55ZawttpTB1gd5jSj9v5KwI49lig7TOECmobkxXxVgo563oZwukzzEbRCoX21zr1hz0YXtEyW
J8kJO4rq4aRBn0+a7cktbkf+jIRIskZdl0/a40Yoq36dkTAEL+oh/ddTHozFND4O1evpPZjpFEDr
VXsSxsfMOxCtiL9QLIK32UjTN7RsWPIuJkHy6yCDQaPGoxttaawx1d1IGmc6Y+NOJeC29ATK0GFl
jBa1poma9m+evEWme7HN/ECfUaCEetVTWC7crWdGN//AoFdLCGpghcmkgbVROQBbzcH/htsttCdP
vlo2JKaac8CEmxd4KUk1QZpj3lv1koAXTnfMIhCK7sDNAmXwxIMadrSiq7ju12vvP5Y/IqglsUj8
rEJoWBrocwWSGSyHmUoIUyaZJIJOxnwGd2yxpXpD63xwF+ehQfMHIQwUyDA05nhpwVMQAQWSFdlI
lbbGGSxWPYOBiOBD8VgUXE8k0ZBVMOw8KUv6hY8Zi2ShtBbZzT/ysTMtGnmoAxlYw0sE09vbF3lw
Da7k9irm7l1Me/4nyFDdx4O9eoamY0Ba6+K1OHkKk9tXA9Ikr9aKSgtYgXBSSXIlbiNOZ8zIOKof
NUD1FyFcg4qGglNFM/7RCMT7ze6tccYzDKFErc9x9jgC6zNpwjDQc9PxF0Xwy3pKmWDd3bVFJvHG
xFlByFpk/paENhQk9Sa7vsC5Wur97FWJkimG1seiOSJ4M5VVQ1BsMP2qGjP3m9l5zL/+WVQ8rYmq
CcIn/eu+QttKc3TsPICWuPzmDhT/DpY+NtSVY3yse3BIiliPF83exch/PB22ob6YeLmXl8pcfNKK
mFst6waR8cYfRL1aQnudIazaJcSor13He7UeK0x2abimy7XZvNZlqncyIiYo6I2so6wC1LQzkAH6
wJW9kZyoqMVqxMDTYb/xgr0M92wdhefm2fA+lXplHOv/31a/OWnO+v6orQj5Rlhsg8ZG5oAw8AlS
rxne+qfYUB8LHdICtZZSKpvOpSyxHiXtNYDjn83TYoeYlNr8ZbJ/rw1uCVSSTdw1Ln5X6bfkvcKG
ISLf+G+EjusKa99XbmtOWwzvffSzrtlui4oKhpOr4bIT6ykmi8GipAxtrLS9UV44H9X843diPOk1
aizq+KFOllhGpNNI85Dt3gHHTPeAoafVltcAkiTpeuo6NqxF6zsxDnl4QdNtWUjC4amkB4p91XAU
NYtAzOUl532GEpRRQPG3H02EOT5oGd7tWEbnBRPdt48NW2lKvxXhmLkE5QMwfAtxeVXSvnr5/RaJ
KLvaZVMQN/PLdO2TL/LWO49aRkDGmDRe5H6B6w+G5yaZO9wVt28TD013i+57x2EjJUROWiFvde8/
WCOOUegdcxlbFMni+OP9xdDeFXnquJkcrCULvW4JfMLl4drMYond8ODmFZVOJ5rW9fykGdno56Am
x6e7AMmlE8o76XtHx3X+OJ/XfsZ7hNV4LqNryDTkMf9uKsT7gcy9X+oRUg7iU+Tb33PSqzStnQYD
oLzrY4OKv+ezO7AekWfWpf2URMBuq7AWnTLnGE5/D6N463V62/VJa/esqyezm/TWkJWQPBnCWjCR
9QvhEHbiB01hnpMSIvqSaqRhhdKWUDWWkQShjv3HUUVyYiVnlxITg1Dz7d0IFoffRFCsO0II1IKJ
uUTicsOX4Q47NchBCqB7pESs8l4qZihL4DXSGQFcKQg2oAa36WiJtSvUE8BPO7AwA/ylHZNvOZgg
6mJEVrF2GpNxeG7MidKibTHJXZskEKuiNI5Bry0ngmxxrgu59WPYS1l5HToBKsgs0WGH5boIUqBS
FknLOtIGWWbsNbYgfOZg5tff/C5eE8oXBbVkzwg6WuZm4/EQkpOutazyxRGcIBJe5sjgxTxeY76I
UtRDIgkB/I39Xo8If4OZKfUZvzs6r8149oDQOOei89oWCVBev1sG30TKULr3m5BdYuxs9/d2BzGC
FZP7psUzEnrJyLRr+wRV+mVdOsYeTS83IKZTAg8ow347+7lTyEzi+teDsxzQ7jULRtNq+8hR+3Gz
LDE7igim+UTQn+DYW8ZNG1xR8TYSCjifPLNU5BY0RsrBOAPqurjd0/H4TY/l70DNtx66mng0TsLh
f6CBM8e7t0yCn1parg96Cb2chMqx7kleYQR8o35FRJ73fLk4F+pw/jqOrKff6FZs0i3A+jjjFKvc
qsaXpiGWmnShCxPsGFbKYbNjQrJ5BPBZcApryc53xlltj0YewajYplydRVYf/5ZopZP98nG4+odt
1QNmAzyadJCwL6Br8SwPUtVj+3/eq/bE1tvVGW2YpnZxKoIUKW8O17OrTHyMyJe1yAYX9N105+sH
4t6kndcBMOB8K15/GxPvIlWoPseKuwnYf59NGGHra5IJv9AvIuTCWaO5KRJne29l2YAIDxnKCXHf
MU7ryRvREnItfP/GDbiyxpun0fNuXRCwISNbQK079aEQ1ep+8vwgqSvTn/YKUVQDzozgtprjb1Kc
HO4LiKYSixuiMLvvSy5ScnK6awcvChLBgPrQY6rSRIm4V3vdJaWvKJe41NdpZY2YCZRC+IdlNNv+
cW0WbrU2DhZA1GY5Rp78WjN32STZNR9Ye2hajXD5/zm+Wr1JSH1sAA1wWt2TM/4KTZ6SRfkY16rZ
hKsoLydBP1P/dqu8Iu2ek6t5tZZHMdpYJPaCNewy0GC6q5+gTp8YJaDF5wkRb1dTMD+YREfHd7b/
aj6kBHRfvblGQl+mZIg6SYL01eAH9N2ER2d8V3EFygurZmJ/HHO9XiwSqf267j9elzeBRwaU/vii
CFu6Np4wRU146DxTJglUlpHMDMow+GxJo7x/OUTMlxqYTF80153fHFy5fDCG7Ta4rmLhgDL6ZVJt
C794bisBoeZP7mfs0Ok/6U0AC21x/hSLvguYtIUVlTTNCyq1k9CZ+hiBUURXYvBuBMbZdzO7puo9
M/SzEPgkTgM3R1l55qkqP3ktQg/03JP80piY3xZTx5C2bZvIaiYtHB75MZq24+m3BIcfQ8dccbym
OIkZBHTvPYY+4hHucOqp8XBy7WlRmRyG2M1NjPdKmmvae1vrwmzi+BVHUnalKB4JKzkvjPinYVuF
wag2cY9H2R2B7p2Mi0E0HFSVdAd7L7Zbz+MgtNvz+qBaD/bBfFjAJW6jSXm438IsNZV7YnMZj7Vo
O7Qly6Ou5mK2d6+JefIj15gAxwnEH/8j3XF63PrPld4uC09YAvY2U73A/Wbiftpc8MPZt4zoaoqx
M6XcAWeMnE5LxPn44znnoKPSXKTGh1mqQo1r3WfLl52nVVjVqQzM8Al5fjGZCGGN65lqSgwIaFgR
/jqCevqPHCl84aL/wR9ZQY68SPMNR8xxkiTskChqHW8GyNvEu/Zi0LlkYPiSOEbFToVNtUuVdAPS
WS1x5g0cfYNe+B6g9WWQquYBCb72uwN0IbxtjqA8CJX8KVcj3Rozu+uvroBuBbN+OPEMHFOPNWVp
ULhD3z54EPiZSU0mfOfcXww/Dig1T3nH8KKf0gdYMD+GY9KCHvY3vtpGlNRWBXY8TqSrq6FFa7vM
q8AVBTHK5NStqZhp2nUxNGrWU5lu8mghocXPXtp58g//id0IkNPc9V4Kq8EC54k12PWeLByBVnBW
yrjCFzLNMsmho6UMCSi+iGzzh4B1puy0Q2zsAF7V5xzBpKzKSoPib6TT1zlKtV8kxAmz9ygoOIYA
Q4eHIgGGGv3Cbmgw0REXMEiKS78jgEI50zF7mE+MD4Lq42K9VqU2gVKpvMsTrEuICOeLXRP2ukTA
v012IC44ROYrBcvFlKXwfJi+K9f2eG0SKE3K1EqLuhZUj9lnDh14SsATac3e+K6Hfce/Q7KS4XjD
wkx0wx1lGX/eYhQB4eyMqv5PYZHM2kpO01SyFUfUOmbo54+FS+jvppucYAd89xi2SqOMV5O71YGC
xVoKB9m4oFLpSAg0gmxlZxlEUderMThFoW11ljI4ZwyU8zSThxnVIboJRbiZJ03E5OUfAaWV6hBl
tglxOEgACUh6284TPj8EKpB5j7HE1JNcLpIj7ojcYRBqaySSE68v4SAQlw+9buDtXsIDAkytGKub
Ni88IIVI8OvweaRICNH6TNUsNbG4DyzgI64vLoV2f8QGR7T8l1fpKjoh5QGwfE83o9AdYUUPhD+5
TnrR91DLZtC0MWy1HtkpaumY5fdVQCV9ighDkubYOf2AQjhp75eu+9xEZ/hfnqcz1hn8TiyuuhWH
SFAZsgey4mL79BjpkvbUqunUWBdtSVIfflOYeVgEUe4xlNdKQo0yH5DRHZCoD2nxZTAtagWSP1EZ
gcm+2a+vbuU0fityExEWLIBxOKDbsW05Q89p8Koo+u8r5byl2OlAWi11jhr3Joa3iB+w8VQKkVLf
Cx1e4sW3+CUTd7uCCzNxLgL272BHonaNLF1N8/hNSNL3Kywc199XLthRy7gXVO6umpUKQd+E51Vt
9qf0KPofPXaUoA+ozSPYx/W4LtKJPC3iQ+G68FWFCWTOuPO+EtmT3DLIrHWeAmNbqlucQ8LVsFBI
in0r3ruyLmWGJN3io+hmAZ6YlEd+vAjEfg2IFG+4R1Q2NLBMLSmnnYmwH6lCpHV2waQM5pmvH34h
dJuvOUqZnuohOxnliXzi0v/9ykdHM/QyaklUR0IEtnYawFHXLhZjxvVstb1ck3GayD72fYNj2t66
612W/Eph06w0iWZCD2dTbvgWfLFI+YfSxa2kw5UHjTCQwgYJ7y4QrHqdcbrGPuDo+8FP/ShU8IWC
CgZCi+P1i16k5Au+pZcRjVsqVV3msIJ/hRs4IAwLCGOen/9Ytj4mFohfwdj5nipfEPNzf5IAZGBm
YjR+DmYNHT+cX9BRCmY7LD6uTYCp6dBFqMICdilWpHvFdkBhifLIiS8AdJ4ghai5woJGieAuapru
QuvkOVox92v0VV0D5/EP9Y6WWSJtnOBLc8AVZstZ1Li8k4HtgILOmrGL2XKI39h7hdrX9pI072JE
mlsEF/EDCFjyzes+a/AkmKYSCjkTARpT6czMFuIQJzeZKrRuY1nWEt/5x6NqZiRtNJ4V1xaDdmX6
RaxDL5kWwT3y4Jxy7QmQmgaqF5Z4n1WZiZMmQy4B85frhf35jsrbjlkHxaeAr81os0q+DY/phNqR
UDay9tg/q8fa7UhkOmDp+Px54FawbPVdJ9lvMzwxAghlKMEulu39lLL3UmwdBUyX8Mk9o1BbR1F4
X9CP5iksmrkfRjJ9P3n5DrPwiTzfBNGK6stSUOWKNwn6xJ6zes4WFJx7ysTmYLj84qrmhKz6JmDF
MGDyweTNdCEA/TFQeC+txOo4e+pFU8xNcWI9IXFMvRk5UyAUCE5xBLYpAhWBSPN8C+XOji9+laAL
qrjCvtZEXAySqNchzturUxLJS8a8jM51VKgTGpYf5O2KmnpumlO25VoFtvvg+j6WVFSY38X3PGSN
jFbm99tmSbpYZsSFgMpmf9rwwfxwz3katPPMzOqQhGQ0+00Mvvk/y/Wdp/8u6/LagZ2g0NOHiheG
vhhNLKY1nlDVTyK5ZtTodxu+/U14oGjuaq/ua3PQVckXn4zGAed66FEz3EDhBbhCmnHqlzq0NmnO
DtaawoiE2kYSOD/YneRtDBWdm/cuUhx+X/IIgRZQ4LYgeC1/2kUqru30vAElXwgI4XOI1bMBpIY6
IP9kn3zY/2oSp4GeGRLJrFIvm02udgh1Dgh3IFizxgnWFnvu0OvLVSqWtviTlARFBKBfhgaYX2nf
cwTQYxM1QPAjbjxF7Adfivh34La45sFBPLlN4ripi/AoFX7nBrgJU+nG/M7UVpEoF9OrJ6WkQPLC
+siuLUAw0W0gWpikOo7IuRBXVB3uVQ8pLRedxElKL6mOeGbwYs7NXQPzgHDrunpODgkaIA+SxsuK
29H/QkqGij7p61QpckFSnb1wqcBWVyVFF2f5gC+wWArPfR/AoYn02oNhgo0B9XbWaVHXaG0GumXB
yZaOOUoLWd4jyR7LUlnNs9iTpSR2Wx3YUIfKn9PlAYbpNb71sUfjhEunUMLL90TziBMQPe+dgoGW
figBRz51Pm45S3OnMwTqdKJdhR2dMEwdhCJ8Hze0zzguC5Bq0LsKYotHb7UORJorl+ZxD7uwErmi
1VX1g+RT5S2iiVFHE6mQEdo2Ty5wnJg2H7cP/cLx3VvdcBVepkm5+Sel3SR2G2vs9WytWXty3cxc
KtQW4FM7fyeKWRxEF4nj/QaHOEVtEXy9ezzwNhaGHdTCr0rcCK0vSlBodC6CJvuIYdYvVJchOpGc
EhvPIpi2vLE0p/B+QbR4IIcMiT5SEInYjtsyJsl67VulXySUKpeAjlosyRv3ZBqGBCvx6mlBDxmb
imf92YpQTjKhZ4IuRmLeFTHBvZCAQVSrjuMHwGXsQ+OsIl1ZM4lonB1VOu/YBWQfwiztnML/teHU
I7+9XJIlUhWSRKCFCECgyGOpJskbRIldlhHt4ty/3i3Bs5J99jAUNMBypAqxxFpDzmSjVt3pwQPP
evTPfph3GtRhjvymINVknXYpqoxneXSzSLdYB18PFRG3vuyTahWR04hrX9VgurmgrOGmvglYLaMN
qX+mHT5Wg4ZAxDgxzo9bUH53/dZkpsulMPNxIt7Cq+yVPYTHRmV1IRDf0o+s1G6G6fALyoDRq5dC
uNab3J7XirWVemIP22SDCuBEDMwAjfCnTzhqzUcJlaI/qMdJ2gGLkc3QtWkJVUHSaCNrLVEqdSFy
Ayou9QByAAMi4xaDsg5UUL5zMMRxg0OTPC+8rIvXg2Hb6nXEgMKKd3yLwimqBDcOZUO12QL82RKp
0QKHtITbkHrpAvkFLb7oe8uzRf3kp7+E9JvuqAuGP/B23zOYD9xC2jIqO8Niw4IgN99qFQrh5GP+
6j+OQZWaTctqJxQaJ8pIUojtTnQXw6fkiBwk4BX+5wL4BhKq3W8C7la6aPzU6Xd1FbebWSK6cQ+u
PSPQjVTs7hCVWz9o/aYgNi072Kemr6qMq0Zu0STQkIZC8vK2K8tYSLymkASxrChM3tkw/dw1F11k
3IZblxLaWMA77/sCktv15VgXGBEt4SF6AVEc9cat+PofB/VPGhpaPyTkYL5b5efygnsDhlLxUP2Y
q0N1vFhSP0XwxGZtdEDnnpccxepuPnfdcWEuQxfZrGryFGW14kntBj1mnQhafHvNUzzz9syVlBvL
TuNiSi89m0Ac3RC3+uDWB/l0rGVOZ91dfV4bzkSK75EPWnMl6PkAFQKEvfvBMsIbgxm2vLohJhDe
UlzsvlXPi9/qU7C2zdqphlMoElOjNYNdjaCKXdjKPjLCJ/KjuWR2bMw6dlydeL5CIXpqndDDpobL
SJJ1UGIUVIVDskgqXPGFfVOLwwz/6c1Nkb8zJyKOBGELiGqoUKmA8qqEBCiYFAjOa466tfO24vI2
Sb7E6tILkOtOUTN20lWQ6ULNvdM7LxDQRXQ8xZrnPefNR819EmhcXwFi4rBcnEU/AHNUXS32MXd2
gciPH0bUiDP6Lb+qX9gSVV5e63LWYNtisjLOslH16ALlaW9u7QXfi4XxIUzlvUnnPOqMzt+kt8m0
A6I17G9UxUFFqk5T9bWwAGdFeVrp24wKVzE11Eb6aURPbYLCa3CWVNYOiXVr019GNu/i63mlJ6vn
WTPQqPv8rsWpnmI94fRN49f1POepyfmblATs2iNC0OWH00xDKoObLOd9niTK4mpjp5aEAW+k8Qdp
HgYKRhNmUq7jivY4mQ/hC8K6Rh5uTcCQ8q4Drzzr3NhxbX5QNjKZY4rjFzFBbf8jCehlyTkv4+Za
618K0QhVQIGmtArWPtmtU/3uuZEXb/bqa0687ZURfA705DgjDOK8/T1y0oC8RNlkkYsb9/Qz6GA6
m4+qltM+9R7hAzd9KBF2V7sP0oeGxBddwyJKOa3F7SCccMQj43C/tWCZsuy8I6OSW2EHSKlMJ8XC
zkNiO5ogOY4JODo+VvscW79NRHpDpPzYKDiC/gJASDIaj5O+WbQr+QvrEcakw7oGEN01E4lX//3S
yI0x27Dt32p09+y4D80V+Jes9CHdpdWJpfBltchHsO8mYcMs7xpFl5RdLBABB4jqj24feb5XLP1L
cp5WVtDXdWv1a8GbK8YIx9ZEYtc4Qkis1XcC4b/LGMslFWrKC8BOLVeVNhijkDEhJ/ZPKg+qxsaK
BSFyKpXl6AXdS66SadsbxqfYpgMxMJN6CL0FONp+DE2uiazttrZfjOpX0EbZ1w0ICW2iMfs4HlFW
5RRrEP7ysD96m9Wzc+bwZVPgfqr+JETP2SYEmhcuSNZ7EFR0Y3Y9G9DljcqO/G8mIyZxqWCV6SOp
8CDjwWqkEaB6BqV9IzD6MVPFBjRmtJDLnC0NFsJf+Rn0Nk63580ml0yrqAaCWuv0YVQXa/k48vpW
HjR1z2ydeKBpt45Sk7XicwveW9Z8U6j91NmpFYSVBsuEsH/ivd9/6S+SuMyt5qOG2zbVeHowIE3Y
QfYafNRqyzyCm1qXOmA6UZl7Qcnyoo8tzGKe+tHC40jLGyyrlxzSpcnzw5XmVrc5gRZXmxiFrC1Q
qjabiTuHbv/H/69U8aeUsAl4D+OZCKHCbyb2rwo+wV5DjG7xyHYQ/rDl364ZDxNWhCudmuoZLOZU
wciEPIJQJll4CnqEXy4KjXIea3t7DjAbryawMZXMweszzfXyq1GZ/z9ckd5Ty1sTwf4NP4TkK1Qm
ZLu2XLKsUsp9CpgUXP8dWZngN/fVBC36Ur99S8P/LAsVXj//ypZWUK4yj//2kegneTTG4OMPI5pc
jmgoaC9WaeeGfu1FpjK6yD3NVeAoj/zNzlA5Z+t1fG0PMIq41dX2YaKMWCpffwpsJbrzvsT+IIt+
jYpr/iE21IcQjeUSSBg9J+Uxytp5i0F4jp9fgATQxlcCzdV204478CuUMZ/s+1mkpYcdpUMd5q/h
OL3wLAZPaztkgsgS9sp5iUsciWZTMor5SldbofCOWpRB0wZ2p6ZEhAQB5luJfzPuK47ZNQDQ3W30
Xn2fuVwk5YrpXI2dbTHXCQ4tujQf2mV/ZW5XdrD9FBWdtl+8lnhTRpgpUVd2hQ/9SmFxoTiBlKpn
Vo6SMTsgNON8dvGJsY0X6vOPyU0flinHM3ORnD91vNrn101mmt6q4X28bU1mBJfXZOxf7jOG6MuI
R+MqC41i7IYGU8HVCpRD2vph1aZsUQdEKOiNLh/LEahVVd/W3+4ru0e7CCIysAagNNpXRMaQhFut
Rmt6ajr6GPTeO1CKTlo4PnuRajVrCj7gR/V2sUIx7/zpzJu10vcfruqAaRx+Td1hwCVzhGw9Kftj
ohRzfqbubccf2rmbp63+MUeg7CxyhiZyDF4Kpzjd3VtyKIt8pq++je9KIaLtfdhjo6UUcpQmrJO2
1ZEKT+5DlB3fF5zpDYVEoyVGVqd3olXkSQjsmFwEovyX8FYBmIRFuhIafz1CXrg774hojsVHIaES
VSpxjVuru36VCV1VF/NAGDZx0kxc6bGIwh6T2Pa4kwJn6IjG+YLzTpgmXThMMduf6G0FrNt4fk7C
Pt+6VGNO1RAZUzETcUcDbmwc/r+LpbwjzOI5MhI0YYQt7lg248bxtQ+KKYL9H9xb5Is1YLIXP9jB
6+V0J7bBGX0ZvQTv7Uu5gtLVhEzBZLdt8pEUTf+2LmAfFcntJUVw2K8quAiVMp0pBUX7Q15tORzF
v0V1j9vzREr2QAyD5YT0f+2KjxyuC/MgxaUU+ArNGwbjOLiFZjA1sQ88tNTxt+AztbgIfsP9TYT3
aqw2J6FJ+GUWyrQH+/qRcVSGhoinD86be0NsPDk3eaC+/QgsFPivAZ6bNuteykg31IK5v12hIrh1
euPzjLM/2mSWRE8WS+uXgC+vFD3vuOCWY1HPMXU0NQmMRbYfIUQQ7s9AZxtLjEOvphIRDKS/jE9O
86qcupMfrcgxbXYrMrR7TmY9xo4ghvh3PWVDDy1YGEDxY4aqlWj4QZzKeL9ISdBQfRiZi7v2YP9Y
Ub8A+BGQtZ5egG5+A2Zi53XqKQ0q8aKIHWALLlrm/60lCI/OTVGlimRsxfQLitdreM8UKV0xHE+u
U0xYI+E9VmIwdpcxUFESFrp7FJTc3JW4X+UMXK6FawwY3ScqsMFMPHxMeNlhcUalA0wFhdVWEINe
9cRkKvpSrNau9KltuuB8HJfcEZpHgWeHHGswG9/uMJTtcMTIi0eApdoj1KvJgdrxRPc6lj9q16aR
9e4i7zJAzJgp9EJX6NoYaOnBdy3U/9Hnjkgjwh6Zn6a78ePbBcFJhD4pBt6m+l9VtHr+I3ww7E0O
D389RzDj6CzYtntHOYRZPJAcvThxdiKH3uWB7ZPCt8fwLo5SgXr0Vwyao248ldtjUScTqub6i4/y
N+zSZsIqnGB/bKWnY/4iSfgapLyRlLhxZAg7Un7JI4OCeF+18RqRmlr2kAPTtMx2PxaMwnnp7qDo
nZ0ho15EQ6xx5aXb6aC0Gi7NXArKIfvloUG2fuTI1LfspRUm0AWwAt4cWfjIaffxwtmbfIpnwsPx
VrB+/XhnwBfNKtcwPMSXApwhoPxnXiprWhJsRgGVTpCMH7JYdj6wwDn/XlAWxMLpwexLlsP02ZYo
9q1ehgVtYYomHjW2LOU0Jzjkhae1ZgQjDeSb9yogHXRE/SXIAQp/0oVmC1FAUodvHOPoNhv3Of3Y
3hM5zCsBJB1DfqV7jsree3SNPbCRmkzB+ro8zbBpcdCJukYY3Iamq7zUO8ls4Z7h0dN6+guQN7cv
wbuPVFXIgOqZdXAq1U7fh1eQvO+T0ErC5Uz57oh0TX6COMqowfLmIQvzmQG/9cFr8pKctnj4jsVU
E/JtATVO3+jESHiP5kHl9kzegcm+bJyfvFABIpaQYTwNjz9KMTVNYkT+irVFr5c/jn8OyjMBCCoy
8WMm4Ozag/aPHRlDtEQlqv+MUwAM4r00YbafLs5tBVSFTnA8l7cox+tsMHTiKnBUlCnxAMfJ/iUy
3xvxzyLxJ+CMqPr21PZSf31EgZTBwtTLbIZNk+XzuZADr7e/alwPrZLlRMI/+anjQg6zJIV8sSBq
Sh1O6kf9pdgUgTxOcZwi0K3zEOF5RbQpq2uQWw1EPqMxRqcEdqegeyIW8c/KG+Hxg+KVZdOs/qjz
B7YnAnkIHbODStJFm7l/EUl4KPB1Ku3R4UEvdWjpc6IHt/CKIEgaArQ6+g+Rd87GzEzhHY3RWKq4
76cKvefkpMOJ8RhBnjeeL2IYeCpAhVcquixbEW4bYNcNzcYPlNK9fYn9DlvS2byTlv/PVnvqQZ7A
8WX/alHenLSGTg/0ljPCNQN/ER0nL6RjvuCYbWj0POZJyShyQYHWXOKGHzO6aTmq4YBvHv3X36BD
go9iLhMnZ+ajaYvL4m3vaoHkNmxnW5agc+sR6+X+MPMFrrQCilt1IhCFv74BFGXbK0zZjp5w2826
oKEjwsVZvOysqZ9C/awtFxbuxhsFisigKvwnXRk7la5ynRD1KJw+OJ4GTVNwmt/kN0R8xGk3Zv6L
7dXlpufnlQCfsipD263NNDkH5F02HuMKQGR/7NoQffHLc5qyEKJRKuWLX1B15nAk7zei7HOGb5d9
7ehdkxlIYUDr7fLag4RdJQqi42LZAnSKoH80UopHCLZXO72qC51Rum8uVdPRmDonWwbZ7inCg8pX
Pd9tkDmbe3+/bgbfJ8bxS0ns5ZcEHcjWCq4Coj5r/iN98PxR/mUTGn9ttSeIXC8lFBZdViTGkJ1z
ZJ/WN7bDFT5q4T+vOav9pwDnQf+7lsGa2gYsXGpvrd9n/Gh7qTNrCmgDffFNvu55L4HNdu6yZY2f
ifa1rMARR/wUgSN257Batp8PTuvneZHXc/FkbzoZRuWhUtb09p0CuFfohp9kSQwknucHcgEy2EUY
AFpBHRIpAHfvWrsY2c6+ZzMRJ2ivO56/3MLDFkMfTQZPiqXHbh1hLmRWn8b1NlGrtmFhJz+dPTOU
tr26aCkdq5wUSNu9sDMdf2iP6c9mDNwnv1CZHMVVsdtHoD8CVyI66PP+2q71PiSmaMPeQvK+it1k
9wau4TN8QOAlX9NMVSHCF33Ec+oU/pc01d64FHR7xsY8Ts8pOB440M/a5qt2LHEkGwHwL9gbQv6o
ACuJxzv/gMaJe/rlI4lMwPc16s4OwIhtWT4j24S00uGpWbqVlngAX75cmO1OC/ZLc3eCt0qDtErO
8BDjWk4YciWEVFnM6/5zrHFdeAaV+6xBOM592RKKUQA4jWqvYfiqfihRz9jOUhNkEzZabelGa3Xq
7mnZCmClxTqjSyD/5rDLDAqsXfLgSXvxP85ZuKyYBG4erSlcO5qpFyiM2VGiCb5TJhw3vliZFM1l
5wpZF2QimuwTRFsbusqoFarTx5NVXMkI/PokvaUQaASSfcumSKDUh3R0bdOQKxwBoGqHNRp0ECYY
JLZnDA+zSWHJ4eXOBNB2Mug2xmgJBApcihsNFYrukWR2rVNKRL0HVYe4rTLPACv95uhtzTYY33yZ
wqJ7HK5BM42OSz4zPVa78D+6qtlXSnQmHkGrIE4DyRn5/7eaXfFBZkSA8MwsSbslgPrIGL0I2Dtl
x1xeLQU5kM3SozhEPlLQh2IC+YMfVpl3KebFSWpOzw6Jeu0iuze5j+EQ7SRQ4Joot10G00OC6u15
QBGuA3aug8fa37pqmdQAz7pQL9iAhGnZWgdV1KRzssr/HhARWQcmYo3IipX2kdr6PVvX3n/vY5AV
lyK6fHCspF6IJLz3c+adky1MsEgNAl96855Liy042UjQanIXXtxhDngg8TuMSu1LVyAY1p+BOUGO
HSZdnqsWbZZeYYHagYZsg2gJcZm6bXvSjTZB4mtzytC40NAdXsF5jwQyDgMitvhsYBkMJHKipcXT
jTl4aB1qWyH41OPaPZVV73I8lCmfsinVeLPYOOEciLzMJRTLkSyRdeINTwxIrBunJtHd123jrJKr
zCMVu9qSfhXNGSX+4cSxJuKoLPLLUw3onrNIayoHCD0WNG3qhA97nb/gNFWvzLib9+wbWMvEbCuV
Qdby6qOiRFlSgbVasxgo/3aNe0r3kgkgxmkwdtPHI2VcWqkLXevDxWniQ1EQLOYxSjmOaPfouSEm
XkDgP1DYThz+AceMIV0/q07n5qv2Uahbmms0vSexa8rAh1VyR/lo9bV/oK7Xju63U2L0xDgpikpZ
ql8BO7EtDtw3/MwGxbq+gBo2D8dVnM7UEys19Psm2RP+LFX/C4IoEXhq4PNdaGLOO90v09KL9Bco
MJZ/6Wis4tXRnMqhS/snk4pdk2u/sGv0F+4vNXQR+Qn2nRrnwxfvVTqRlvDR0L8LUn8Kqlfi6gaL
txVmRJNEKBdhwfyS43NE9fL1O0mIwSmcFrNqdv1oBgI3Yk5gbDsqMzG0nOFZ1tgcI6NITsw7v/Ga
V4WOMsy0trNfGRypAFqCxyky9bZt0ujWP6RLNG9YCNW6KDfd5dU6Al56nPlSfI1+ZdEdiDijBLAE
W1uj9YXk5qN/sr3fINgqyMjHMsZC3Yzwfg45VuayKlHjxNHa1vvaFVZDCvQPrvnfX0FTPTQcMffl
IH3mUxt3KCFjrrxL0KTv/dLYbAKmHbo0drDBuICOq3dLCSw95MZiS/rutr+lp7kupu/wMMP0h/rl
ZIQtcxm/8QKUQOIcNF86sCYSJYPNBV66njUEvAlhjsmr+wBGWm8dZPaK63rNBg/mrU1WCBuYjQ/E
syC3LygaLHS7VdoWCFMaYndBMdtoVHy8hIiGugIdobhoXam9KZDa/JAvv197ephGm3CNX3O6t81S
851nBz6Ieb7ccNI/yHGSeA6b29vNHLqTepcHYot4EcK+r4roV0JHDj8ohcU5ScjOiSkuGzf43nbP
rXdFP6G/7pC8k8461HvBHQGjEzaCt1+ERiFjT//1OKr6bwjwrzUsVe03rlTasK0mXJ/5YKywXUH3
gHGLvwTdRSsNst6inYYl1pIanf+q+wjSMUSSKP8fXAORIxgmBvYlqC/lI01gkHZ7lbb4POAsTwic
kiO+IGi5ZS6wCTfePaX4g/Su2h8yOtR2I4uAVU/2rOVBqdoiutHwZl/pUGPuJcF7G7IxGau5B1oC
XPI/IuRAH90Cir+JhVzgk09EMP+OoATDEuWA4SMT30CNklJ0XDn267+xf8g84kNSFh4NrKMWCBhk
Ayld4RCssVh+AB5gpJn0EVtn0stJ/cjkyaLmLY73SR2Q0bwq3jleRCC3YoU567opnXZrlXUiatPI
4qjtSoeispKMwApzMAEXnvH+KA9XSJiI+enVE/uJD7cPdItTBdsJ14QFkhETMzmHugjZ5eEbzPkM
ECtI7kX9PO1GnhyMiNTNXO1RFUUpDKxES1UGBSECkonh51YFMgPJHv/0P3mgabCf8l4MJ+mTWuGE
iaA0QKm+CPVqqKpWHu34rJIKegaZwRv850xuppTC08UvkdlOnAG1XQdrJPintfgDRr9Ygs2eZ8ls
+xaLAOIpTkUTfGD2GGxRcUJ4zAiDRbFCjBhsB/Le9bou5TNMFCD4bk8F/mqW9QaI6z0CVc7y0qlW
0GSqp4N8EpH5CGP7VMP4wwhVQVloIKh8jQiUH8vMbPbwYeQ3sVJAA7rHQpSJxnCF3gy9VfRtFRiW
m26KBR0F36kC3UoSlo6DWoV9pmzdGUDOVIw3GoLYnE1pU1y/IbRfngEAEa9EVauG1oebUv5dl7RM
YnAmDjlLaI8bd+tisGfH95GcWoSRtsO8klY5/YF3+zwdygCF5p4FI+dE5WA/VQvFJh1Srzw08cmE
GCuxuNFUX4iluTNsv56PQIXxHXEyQzDRrCMZJYIQ2Bcd9PB5nVtWbBB8UYF0/kwSwXus2MtF7t4s
AxnpcjP8rF7mHtiPD6lBfBjda5D/PQ/uI8hGCKcy/s6PaMvFrRt7f7Qj/O3/3ZSwnrmZQ8rRqGDk
E1C6Pr2L5eyINgg5jJ22ACdBUgURbru9eBS6eU5JxC36YVNdbntuL8/jcuHvhTZFQxk6giqvmYag
OH6+xDYom2HChP3iYO/LgGfvjuGdiv95+SExDjnL7cJpp0E5lg2g+WiO9qzR7g2Q5xEn3rVFOHX0
gmaBN6zYGzXtCkAmxz3SEOCgFssfQD1UjkBpbi6lHZo/ulMurhqDzHmezOF7oMDzkadiE2kOCMGs
tqAP5FJgIKg6XXfMvCoCXQyrCFO/ACPO0nmTbRpEHGkYY2MZrG4ByxUJbXNl7Yk5DcY6CqKg2bsa
37Ge55u3Vti2T3ig7kjFCu27+RmTpVoQYJDilZGm8tq1NHW+EsfEBvT2a0ZiGta6XqFkiKC8Rbrw
TGpYoOQrbH3h8kZfCTL8ut+Dqbu5m6GtoEjc7nafgL0r8MUUhiCBNmIOmuJB543NuN4offO89y1M
yfw49HN891lwE37LXa4d399Uj90A/vE1t/FQ/4PgXSaJe1TqCOn2N1CkUBMKwmfb1aQIdR/uUraI
vfOHlS4+CotMtEmJQ/YMUBlC4JMkCLe8c1iYDNnharPvrtX5d8clrIc4Jr5Bzrq8WEq5T4GY9xBa
N6NXJTYbNEpq8QjzUcIRDVVNcWQNe4x9Hg9ImVy5P3/U1xeR9AF3dYlCk9IT9s6z49atRANgwi0n
mRGU3f6hzgtynXixw4WcF4/3DdtGgO2fI9h2YWs+hn+v3rpKnxbfQ6nqQQdkXVWvgnE+x3Ntb1KU
RQ6/HuUh98RFYe2ilKCUYzSRYgEmtDtCN/vYJTBJ7fIA7QFnGIptFdrkcqsSafjUAUih0ry04Dpd
gragpktDyMiDTf++HN3jpmWQt6PzYedNlKp8FtQbNvQL+uB5c5nHepknlvWUX7VNkWfXKfA+63hC
6lPLnCj2NzsFaqf70bad+yjDFuUidHeZZ42Bio0wAOp6BNV6Ijti6GzRhaD3Ng7ASjMIdpPnL46T
VHBZtnxPUQt59J1IXo8SjlMcOOf9XVHAk3TJvlSBeKULSU9gc2GZFPpVtC3niUtXfh51kb85T+Su
fijP8eotEXUodCIAUG1cLTwe9wgra3Mgh/fkbTWdPAp1sJmiT7SUwQzI2Ah+XoB8MRJiqJjQpvbn
ukaYv2nYcaXAjJLtAaPN5221H9Vqt42tC+K0doFqdeFIoToiAkHyCveU5CUvkU1AJg5dMB2NnJHz
NCQR4hFov/kqmzK1u7o6Q46i3+L1Zb6Xl6FNACDrgenmNw4d2SVvYBHzEfKZbb9aGlTC6mV1B2sY
DmzAgc4qOY91slFTkpqCS+pd9NEaVX/Tstd731Vmlh/pV9lLZrEkoU39rKli4DxuPpXbaDNG4ze1
AzPxADOcItOK1BtD0FTzLejQAlEHYaVeIhMo/bfX714n+l9SVY5qo11xncepw1KykU2ahym3ab6I
OnJfZgxc2vJOD6Ldr1KmwKT9PLSGDAOKNNuL2gthhEh9HpLZu9Jz9nNLQDAydEpNusM8/FehHrK6
D+DYwBlV9Rd6DycoBvDlK93kFWrWc/4eFMqs9UJ7/nMtlAaOt3SFxqj6ZrRW2AYFngsQgr5twaJD
LUhS7IEf98czwC1m+lhflvWhDNrt5Hk9oiXI6viiJoMtzBaVCUaAQWD3dbqtiyBCfckP6lo3aS6T
G4Pywa0f6J+0NE/HFKwGhliT8DstEkftnaEzNVP1KUoH9o6mZfhTclfsBINLOyplfw8+yfAZr0g0
zFlfDg+CLRVrdwEcba5yTo0MW+Xc6/HdSAX2DSl3PES31cX7vJj1/ARJOaDuFYdExbuwtR6ayJfo
xZr9g2fK9rPkFCWj31iscWB9P5IyImEUDvhBt9+Qnq68CjLMfWzSgx7XIpC0KWBzWqGA6zNo5POl
2jKg3nr51U0V9bTV9AmelLIl1n1kMexOCm7aQY4iANayT4MuvoSUt5tFdfPgeHeIkMnoBcFGdzGr
iP81y2FxugFyIgsPlQkvbmlptMNulTYQlTuZRBn7TFXw2ODyY9BzN+qFMK5crzVV57GyxHUBieRW
g4DD7dXpPCWJOtrPY9nDMWWB0EfZAK7sYLQxZnrf0ae28YUdmcmeEb34ejBBZKysvnQfL4VvYba/
ymzJNTuXFXLgfpVoWPk/Y9san+bdr4QnCz+SuWCEl6SpOvk0LrpE9M3zHPRVD4ZkxYON8ISiDcE0
sa+QUzFvvSVebPXvalpIHuWfl+Gr7G0C1CEV5dzcnAFme1qAXQKRczTGXNuDmPBt2irQsl3jRw39
7pAFnd+E5q845skqMgCW+rDhFM/yEm/w7DkeXUrrl8m3HuoXLwUhJ3uOjmoZIWJn5I1YPiMk/QkP
w8hscCuT0vJlbpvEXm+qeeJsOCySecSSUC2UXU4WFlRMgdLPwBC+eT22HNnIJkOkhYCrwMhTo3Jh
git7SfJKQTrfvcJiOOOU9RGspBsG/9y8prTYly+O+eM1hfn87k50XXlKSnW772xkruz9ngNXnULp
bZ7EsG5i1hW9jcBiS5nLvcx+5drkHUSXzAF5S0hVLIcpxRGlpM/27NDvrnUZDTkggxJSzACcYS1F
EC84i9rf/oTdlPVr3Yj80byzDWm+xnv50qoOILe7LROljsDvYpq6Ymy+kkvIDoNRZ3a5lTHScWRl
DDn9Sx2GNtT5SigIV8YQuYpONc71kgSdcNIY57NUxKeHY7svskUG8HGP2V6IH1VpaGcxyH0BaMOf
zIAqMVUluYZJCbo9jZKSmMJ2bkCACeFUaHYhxeV22AtqUEYBL/HywsWm8y+YY4+nJnXKWQMPhrE0
AAAYDR/3EpIZnqwXbXwYrAEnTmDcelzfiK7qf0MBJCYSh7YcCAKXQE/avHHGaxhIeTwWtRoRbBhv
X/A2PxoQJIA88IDbRQatArw4JZQn8IPudA+wg1v+kiyMLCo871UPdtk3X81HYqW8XEc3qxwVe1HM
m4jjfz/ZD3D7y4NL9+4FYf4diUJV9iOD+gNG9JL44qWavmMNoYq2cs6yYhuHQH09kxfbPkXBtxzO
1TjtxoltqqsxfQ6AZH+HycXX+Jd+Sjva6MYlIvGpNeDpUGf6fQoy4cYGGSSyUAvsNX3UmOAIfyHk
fq66yr7FOCXU/1Xi3EfgLE77gBrZNUMpM3Op0TGZojHRDZlMUuMJlSFRc22WLctQz+YZMFaczeWg
puo7Sd65gUL6hVGIX5ySMVneY+4FugJidZ9/yelB4ROgNWNNMusEJypI7GOJPr5AV8NSMCiPdllY
W6W1W+EuHGlmJhKkGceiZHaaiHvN3nRyPXaCKvARCosft+dT41DypFLK5mTNwJNUBq5vmwenLYFD
L3ff9qOnyL7LQmkYUa0YMErEJPmFD5N2mhXSzg5h7iMzIqBTtZP8wFOyzqo8i/Fm+Cj20li3Fs2a
w66JIb38Bq3HGfq7L7sgxtcXOm7EPw1Vd6aTbyvoxjE4ztCanSAkSAdIirvJAL8tyBpmjB44kLII
gM9ZAys7YrilkFj310ld6YX9i5ZW1hRYurpkHBfqIYR3RqjtO8SyyN2lrTQYEmxTS5SRY55JJZZt
y3W5QFcG/KROBbBuGEZMaGf9AEWveI3QciWX/Y87fIdzeula3OGtUTuLF5TO34M1YGFQmLZR8t+z
d6duLCjJ2pW88RB1iYXolVtRKVxxt4MT3DKvhR03AcLSY/dI++jGSVZo6PSOiotQs06V9fNyrEsU
ggLXSSyrFTz96K8yV8LpbAdje+PA4jNAsl86t0xYHIvFk6atHIfmE8BG9yGPrerCln6t95mJNhqJ
1QkRJEkHuBu51/ZgQEgawbCKFtCd08ZcBOuPzblwT0r91D4gg0XIi8rsbn3CeRLshFsY1nJN+Ia7
dFER/n8OsdzePAUQF6mHEBsCNlSUkVtvBs0riq0dfNdgvYTVQhQ5jFup5lCathT17wIYDFxY5YZA
6zBLJ3DiqsjTjcx2vp7F6eT21a+Nu2+zRL+qsbUcYEjdJ7KqdgGhv17FsIMQmMsgGmK7KsfLZdmH
VkI3lFdEcNtKp4BfnrjfuSVc2uqbLAYgWfSnUfKWGTsWP8UqtOuZXA1QHXx1ATVCPpOBnVRRbk5w
Ag4g+wp9iQcW6EBYSxxxglha7RAOeas3ST1wG/XxCEyA1teqfTagnfwAMtY/qKDzst12/Fba6d2N
h904iZ9MhCbpklanIhEf64EqaY04BG7eh+nLIPEPMar8XDgD3O2Xk2A+G6T4Mp4Mld0d4tGzsYlf
xu/cwZnxptx7SCf0687Zl1Atym606qFJrbpQo8WavqnVNsrfS4lb7C/tK3NUUjOCUD89/1wF1SI6
vbGP1RnkbK7XxQFtK50Je7vTAI3k/GpscyNdve6jlz4a7yO9H0/D+ksp8ZtXBDU6W2fRun1/UAG0
prsuJRaL8GTnkSr+ZIR+gBq7kDnhO3Mv2davQ43xxzZ/kjnD4Yqui5fthORziQNNvguTqNP8t4OJ
GXwqc75vSf+0yUhX+dyfnHJSeuFUNFiFukDPgLtPoDNVAYCBBh/q5YL0a74SnC1HT9t5cSAJ+B3t
4gxvMcQxkvulvW09btDYOAvepDMaE9Lc9bpm0M2zodtCNPG/Fq6fSxME82VcgbQ7wBdb+wWiOvxU
WK9O16CSycU/+57CfkbE5kpruB/sDAcxHht8veeOKCiTx00tmV/tHWrjcdya1DLE/AHaVdG1s7ll
xuQM2YVsrbbWohLZVpZdY7n+NOPxdNbOXT/V5mRrSo9t6RDbobkcB1E5PZ/Juoi3tgCasXGowHOH
6KHV4516zjXzkgeyqPULRLnJP5IINuKVNW6jjZGwn8aZOXXxje8Nly7fbM7S6UkhWC3cDky4o2wj
79GZ0IXUVm6KnqQ4Wg+PXQ07T1xh0whtuKm8KyB2QyY5Ga8QmXQZ0wj4mzK/q679R76SE7Miv6R5
B3rdDnuyKEexjZNUjsZd84eYzO9XdvcxIDDatoLxgC4cJy8Lk1wqiIDDbZ38DMvXes48I7xXJGpo
ugVq/7E5OW1ifpBfiE6GNRZkkNlIhDS1Mo2RRew8Y3iJrr3ZBbYVDCGV36spzvQbLz8VHfqu43mU
E5d7f4laIDY71j5EniQ1S7qCc4rTIkug6xPPv5VVmG2xfA2rAs3g0m2spmGlCLWSTuLnxq5SzfPz
WKD9obsInfmkCGVwb7lzE07wHlxUenRYHqb90wmx/SgrRmp4MdGElKjqmV74zejiggZ86G8O3gL9
SrIdC/uy+gn3nvkyBkPimXvTaNnVy6DU8uVTUcVoI2fdzwcrz7nPyLLay4vO27nNZ8H9yytazayJ
5lN4ybbdKs199Iv81GUw5YdBM2eQxPDTaJi5VKeMcA+xcBc0bzy9Z7VollTZ2sj2U4mVfdzdaqRR
afyyTGCKCofsBO1agHZL2jzJMEOtk3mWT1MpkztWhMI/JVnpc84Fw2nlUimz6OAge/QpDpnERPXd
ZP4oTyo6Ck4kFHvP3z4zgbGdu27jLYAr1SMROl1lBvIZl2m1oM0wRjgMu6Be9IZxc0eew+MCMQtC
BS9S0oezYadqa2ouInZwLwlp6TDNHBgV9unoAh2ZdtrZ29aGa6847kl0083O1GneRZnZwgIXlTP5
RVhQPA4U8Vn3FxLwCl0opVwjvPWnvq3KBAivLEF5g+uZlHgMsUvdhN9Qi2U9mRYL/bTL6tumw/TT
d8+CH7uRnp6xqh+XEqomEgXcMalBsYhcr2QGX9co4o/BsU+3iJdMhtbyc1cGPdkcRtyjYNnmzZnT
0LzDJ4lMExBrCYzMKIEDDyY6aerGx2UiCR6VtVJRVMA8/qTohwEoEZUa+O9v8gpNcZJ0tdOFdEMu
JAoS110tETlF3OkYBHdnTZmx6dQp15CfqmcbJSI34ozJkmuGze+R+eGbWC5bwp+0QAyB9oWh6p9C
APHbkCs062/sjOO7VkyGuu3lUNcXwNQ4bjbjS9lDwuSVSgOYnyUHOFzW8a+Y/bJLADqHvwKLRj1S
JKg1kx6mjS/akqOulArlHZ/d+YQTrD/Ny6DbmHRGXzSLZGE0y4Kc0vvX7/mRspY37CivsEOT604c
n9hx+wtuREz+QapDLpyxIzrQ7/IHrgEimRJtD1GscJRrwhuXLuJH2Q6064++r37vN9XP5FZxQW38
l6drNkpKOgBQ+HlVkBWPbN4BV63QdtPLNqnzMTQYaGwHrE2SKeDmIe19/OdCFWPyfdKRnf7ZogW7
DIiSdOTOEQz5gTS8XVRPuLD92OTJkLpoMy7bBn3wltUXjPpCRi7GOet3DOFknEVvZToX3z8loGef
iMbPs0h+pAoVtxQEHg47gaHLe+hoeLcn6RD/GxdN6/uuS58tgvaG6svQwsC6pSdqE+O1xynt2p0N
v7vt2fUDfFT0PsOH8ETYJvwGh4UyrY6LDrQgB8XPFozjzKtPvbDNeHYdzy3qkuyuhR4wYmRJ+Pz/
/wnyc2IDYWG/AXNhywCuagaXusXif9XwiqTdAtGCS/Nfqw1a7f0GDlS+md3Mc5lqV9AS8mzEMCuh
Ko2ZRqqA+EMdrLXigSxWXYmvXk1/weG73zihQvnRZ9i7ePsymYqz+wBxzZ/0RIFve79ZCkHaOuzw
lFM7sVt3IfeexM+munTvpnvEJwL7dLdI5gaLnwAD76/MnB/xJWgy8thJ2s8rRfqiBNu0PuhJ/XXs
m/HWv+dqRjmPT4qm8VcA+4kZXIqyRh7/JcILaM4FrQypzr96GfGibXYKeFz9lFeYns5EAmtOwv0w
o3nthQ6MvlSyaxkV7K+ide3qgr3y7iYWiKTmIKqAj7qTrdlaUtmnvo46mBDhhppHB6RzlK+oS7co
qoZkseZ7q1PwMpXmyImeFB9k0zV/f9H7NWR4erakmvYf+ALnumbckP1/jAhO3wXN6Tc3NBCGnjcE
O6QC5th3c38lEN8PGntWUlQzootZ7b2zJPEeTD3Z6X70lsiOhl//ew0aCl7QxhBujtF+B72gCX6G
QYHz74J893H3ywpQXi481Et6dHbXMTuf/e9YB+/F8MUCk9Ufl4u/MJT8+Zukfd7NYp9LIO/nGdep
HWw1obmk+PKA1VZ200bw+bUL8YUjuC9AvWD/HZqnIcvOx18azGhThu911l35HQPoj6MutdE1WzSt
EM0v7nEwVGsXQ00DYqghLD6kaFighnIOt/b5dApxtr8D3peAGlKTFJ2Rl9znopCM5SWPH+4My5Ac
2y1f/1Q5rF8/CODGCb95GgsdrRWB2zUr4rQiir03ibEiKvT0J5vb1xNaSUJdIiElY4aZ6PQg/S+P
FylkNWU/sj1fhtEuQjuw56hO4M0+sz1HG8qB84Aa9Bs3nlxkUmt318Omq0lQcvVMqR/Ztp/Q08MB
HK8PEWiS5uJEamdiVCZcsNNuNo6R7aGjwrgn/AUl0SidVw/zmyR6rxPeUgVxDdPX5XX+7GlTdJ7Q
ElhrZCebLCfVdfQblye/+JUhQ/jETRABwa5K9jqco9bRV76wYeO+/bEZ8LXyb112VvfSWoTmCUYl
/hM7hLyACeKKXH0TbqGtu/ue+a5bCTPtNT13Jpm30GX5YCLPI495cNWDzIR4NyErVVTMi7UOp6vF
0TAz3cgSeguSTwfl+7+x7qI87RarFDKJYfFmRqEICJLMYN+2dm38qOEgEflbh4LWqpvbc5iPdbge
UwcfmSXcvEv/lfba/JXlw19eVKuHm0Kw2tlbVb7Ug3BpNGDWeoVc25rMZ7/Nqfp4x95/G7OXrok1
XnkcE2LVCBCgyh+kan9eRqKRmbM9Fbu1kAhuiH/ZXaG9afg0kdrQUXGjZ9vawojGebT6hca7ZvgB
oXAGN1xACHKz9iGNASAAMrYutYP/FlyvXWv91/r972FD+MO91ODzlgc7s2Eoz4alJFlW6+h+Evqd
OWYs05Crr9GuUsjDtGVUPa0fKasjICDHalwhcIQX7x+UiY2sNmc3TNhTSBE92m9iKWpcd+RQhxu5
Vjn+2JbGOz7mNPOPwsQ5ZvWSaFcng38ff3XaZyjmLIQgh7yAI0Q0G+gntmkJPIaySIEIsSO7iBJp
kNokI0NgKQkuDEZP5PdA0V9VdVH281TK0Ig1IgeKyBBuDgVGl6m6wSUPjSR2zA8MDWckRx8t2W9x
e230P4b+PhBQQbcvURnxKSejaPpheQN2PzFFocBWaqhxayJ0FFNkPRPOEUkftQz1qmicEmFa0RFq
aFo/xWItjreTKqEKg+Nd+3Dso7ek920mCNLO66pfgDxne3G1v63NGFFTI25esq8zYGeLjmeB5yWI
sxlTyq6BOiaqCgr8Iutvg0Ed2/qQzEwupfWKob7VbvoDmi1szwXnV1pWuwXUvLSG4Ajw22Me3Cui
iGQEbdmwRaafHNFRFCpXAz3f0RIEGQXUR9iFGTSdaifmw7rNbOiBRYvgJShF75CbV2cgp5zPDdjG
1cx+qdDTerkeKJbt53fglcDEJR/4wTs2BaEmoqpRyOnsbXTNH1hFc5Akcb6o2bljag9LFF9fMHbI
oT/HM31KOCwFE/CskFILQAf4FEfvt0CyJ4kVb5CVGgSXwyygTeE/6Zbidfw6qR/dYCUdLn+x65uJ
PqVD6sHF/yM739v9GQU5WIo3PJn2lq1CXT8HqYHoxkpakP7Q6lhZZY9D4pN3D++MLLpWEKXvIlQg
F7+2X60hgrTODI6FFF7YxhQHchwCgDyIBmc3fB7a6K5YlMaSq2JokuIhv2s4QecrO7zpLRgrzyCg
YVxFvOH91o74yKVp8X+hpTp15JM6pHiFPXbo63/eDxRgEj2UZ27dcjfuwF2EQ0a3zA+S1o8GW1cr
Sb7oReHYnbY/LN4kGbCx7mDZxrKKJHLfEitg1z4U2nb+LCe0XKhbl8x2AgB4p+4ufMnEmiRXIEAj
S2Cspir96Xc8vU1MoLqtBw0tyFNsBTPuW29kr0Tngtk3dSIz8IIxvodvxu0n7iqR8fKnxSj544xk
yaegHsYbvs7/si/mN1wd71emHSQ3fK83dF8pQ2wnay/eZrtNv8pjJHInbsUqztaSOK+KOTlTDy4l
rZJ6P/YtU6v9/6RvX9Tz/qLYGixHQm9fEaIGMr5/Z7suh0xGmVOj2y7f35prM7sgHXEg7WmXVixA
yTF2+z7jbCuesjqR+otwfXADU12h+qC4t78ebZaPrFGdRdtqHLLC729n9ZYNdKRbdmhK6u5O+ujz
9gQQosKGxLJ80ZsDFHEC5+C1E1DRBiTh9DdAXO+838W0UC6iIQ7hMElZwtbts4rR5RVaACNZ8yau
EaAsyCTw3dAHukrMTahr9HYOYIesCVCx8Jzvv/92uDDOZ0zR7EB7Ds9sr4wPspxljI1xMVZ+qmzC
wPk2mq98BILXWjpq9QBIaqPVw4WinhS+Ulx5SacQIHZzpx7f68KDJAiuigqBFnrPNuZHaVbouWuL
aOHAotEopPGp/3aQGA192OiFC6pM4W8QzjYmOFYuFxtbg/aqWwo/w5pcwRcD8309pt3L5tcNwQef
NIVENsMd2GytdmCvHQdUjB/aXRKsV1cc3Xb7mvKq61LUmj5OkKhUH56KfO+FGaCX5Psd40uqDp80
YWItleFtUVWhUXkNELOqE9wEixgcRfAZ81gE2IDT9VKNvLYSIUdmDerzFTjjA13wcBvCPs4fbOvM
4oTRGkBwo2NEzhgAy8+AdhG2NTSVd4BzxqMOEeVSGEoCLTisQLxzNTeCG1pfRJauHMO87n6SJltJ
QXzrA9mIkeTRbdoMpGd5Eq+ZXbMNmi2RG0WFCpF7KAuRzzEXG65Pgjga7ckaRSaI2q0pg1ZrpDij
+DdKlRPT00IV/S1KgSkl06vW2DM435T5ClPGaRwZbJ7HBcqXI2ggQTOHMKlBEKffe9GvMg0V01Ag
2nY1i0XGJdcIQCy6hPhP7aK1k9PJEEDS2B9mAawCfVCEXn+8wUWtTwc6I/fJy3l7DXpAvuS50mxi
eO9xWyL397SVwRr7exTWb4bL0h99N5LBI5NOzJ1w+nzt4Hvv6TBMKIslt0frbFW5tk9cFbOIIsKW
Z46dYftihaHImuuRZffW8DHU6Av3Zc7GKDXisvDVgC6uKI+E65LdJqTAbSBjaiNfxyC6k4sWRztU
Z/c4epr9q2p2DpWT5rBvHmiUzeLuQZg6INOv6JgIu19YLxK9b8KiWsZX8WbnhjQKNA0Cu29EGl5n
veKS1nLhjcin9WJ37yJHbMwdje7faXChACrX3TOuRVNUo3gezmkkQqu8NUL57huAYDd00CTC0Jm3
GRlcoHyu442PRMSmoy8ArxDsJOVt/H2+cVyeChdHMQzKZKRjEUiEupbTZEggQMVM1wdZInwNGbDr
w4JWLLYtjT8A1fkVvsWyppsVgxjByyzaSkaN/QzFd+DbJP/jNTmMkQ0vSua7mcM129XbOSb9Kd0a
RC+qS8cnfPwZWcJDRTEdnBu0FCSZGi5BktzX5iFjtaVK45rsA408iKdSNSquTS8DqdaE5upXO1ke
Qe11KhJg0sSuKbkXC2xbW1sSgR2rLEuyWXyH98HImaZKMMgHrCNiIy58ueRXVjaMq/bkdgYnJiPp
s1PS+OfH5Et5u+LdwpjskIhLHEE473lWlfsmnrX8cSdC2lnsuheC7LQDUzYY2cGCAX+aT1V/HSlG
1OA+jGAYe12uy+50kiDv1O2O32XK+07kp0dpCpTar4qhQda8APNzSuIVNPzmVAUlK4OjOpJDldT0
g+hwnLvp9qdhf5Lfg0ppOuc4o3QqckRhqWfJidt4uXIOXEbfhyzargaH9Zdi1w6f7agVaRJVat+r
pmFsE8hd/b1vdgd+bgHxjKZB01NjeoJGwbQOQAeGufOIJy2JER2M4JGGYz4n8J3UEjdPK8/PsmKt
2Sq8H4nbDRJT8SrIi26wPW1/EgWEBwzZmkhIuj29BvMj4dkHTi4zi4o4PBaZWrav0EFMDrxZl6Ne
XJzD1RJYkljNHs5AJjYnKfzgdToNRJgq62dPBKrOagmaojdV7Yjikp7+vPDYtw36FCUYAs8pMg+y
O2lKTY6DTP4sr2N29yeLVmGbyJHtaLTvRR6eRME0uLQsagkNkZzg65sQicEK0ks5WmD+SPvA9Fp3
bKYyKF46CiosHr4YU7KDy47NBq2num5KGAK8dW8bAMmU7FPiJ2SJ5TGwflxwXxAEYEtoXwKqnIzW
ek0O2sL4BJzrL8CJvvgBmRhjnlld3yIrU5ai1ED/Py1VtWE4uSCYKXWY3OZDmZsQOS6MF+P1wBf0
IdKWbxh4DHmkoUP2+l4R4H50tS+FkSvkQ+8WWQEjrRKoYPo7QDYIngUFH7wqHPxpIGQGjU3pP9YB
gkukrYTbmkZGIAujDO1GFa85lks7BPvqwV97/TQf7+DSD0AqzFRJTrd4VSv6HSbEocvg8caiB3mc
WdkKQwvj2BSuxlQ8tQ5bBy43TrZXQg3lvsD28/QcOkGK8cmPUQOlZdMr2y/erUTeSYGBvfEuEPfi
nhhU0CwpIjIt2BHuQLl/2Rs79KVkpl+fC4E4tKNV48CYygiCe2Ypr3G1e3v7A8hGiWJVNxdSlJJh
0EFmTd9sRWWQvuFoVZADWZQBgVA7b1BHWc28In+cgvA6H+JWJhsfA1jId8UKYFx08rNQAixRQBxq
BD/13AYdsXAeqxl/KA0sINIkbuoVsStqo2W15jE+Baw3FWq4s8RwrzBKTJFqjwmUuvACroUM8T88
lk/zAVP8taGzzXhVC31srlrla4WUXOhyiqlhzDr8XXs3zwCm1r9DMfXBtQF8flsn10AsQfts5rsd
DTrx2c1lvywJQT+Ooleb5AYEITLqtPbbnKQPd3LI2cxvkX4xO1nvVwq5ungBK9/uLLlHJBaNK57J
gzsHLg5ZmtK7eH500y6iZCC8T4o/iEt/y4j6yYtbMgi6+G4HE9pyHaaLSNCarjWHApAciQgfTu8e
qBIN3owyeR3S1EU/NGCueVNEgPHyv7yxc8VPQmJR7CmaWDBRTECiR3/vAydAza6imLGPCR0FNVBb
y1dbCsklTLqbFogWTlI+LEUScdSyTi+AMHn2FEwz1Kz4GSEj1fBO3YMc+F3M+K4j8NVJiV5bKCMi
8/8pvi6Eq+C8trGlRavrsftq9OQvj6G+5bQgPLZNg9na4wzFrhRvVp12jy4PPD0u7p67xy6Sqe/z
g7zYCY7EmtJ/Y97DjPFk/M+kypgINY0ABcEJGy/WkCAhvIywbz501xNncf1rIxvtbFHnLODgrs5y
eShjrXoQ/aXYEREaCPHIyGG8XKvgfaWt2B8bdeRLXm/a/dxkSaF52kZ6zekT3OtblkKtVbaPTzly
95vatyk0mLVJ6oPcgAJpO/99pvBSrxMYAaiEXybOymZ0rHx8K9EvtIfAP5xj6W4rfHDndUWPeRG1
nbiAV+Yn3c59xYHAvWv28Odpar+9Xr+SNvijQActoJANBOKoH0dZwHwB5efzSdvH070uToQBkYSo
mTXPR68wi7s5R4gulHONfUP9+RxozlqyXRm7rdlm6/mAFYxYKQTCcjKt7jxGHPyM7IAei4GxMvK4
SBTBpTlTV6prORSiRn3Cx0wLXduaFqilxaU5VRtZsOaKlIbdChWWW11GOBOYLvCwyaBbTxEt87Xg
CfDs8GH0QVlH3+iJwP61ZW03qF1c3kTlyozSDYrlzhrWBcQnmn9GlOnuN61f3i7nzHCRs45o4X6c
2VzZ3ZqMyvduf+RMUH+BtA9mZdM2cRW2DJV5XvPFAc0Z0WAfrKSIHOmsG4QBWluDHPo1xhWu72Wn
G+VO/fZsFVDn2lZYaFeLav9lJQdC5StHTzqd+oEk7U6r76n+63nhcG7a0HjbAmSw4vyvSSziqEzn
YSA2FuLHoSEWDXz3CDXZBpZR+10raaKlfJB+5X6dBCsDfs79fgXGABAyuyqYs2B0qWKbPyd1HIFd
dYvG+evA8jsW7dufCYAnKVyIK5/0yPRXvrnX5T4lhr/4oaBRROofCS037+4c6Q0uoY7hU6lYN58E
cGIjKXtHnnpLzwUowBKnJ7nC3A5RZGzvveyy2kFWj/I5KY8iHqK/c0nq5iFtDZDbo2FoNc6fd4Dm
LPGoL0dLGUtNP5nwGM346O9UoxKM1gjTxKoOO517aviVtYKpSlftLTfeXKCCwVm3OqhNAN5Mjfp1
G/4ItdvN4Wr+wK2QT8i+dOHL+cN6XpY0m2uK78BS6fgaqzigcqTn7O4Z8ZW889LG0pwIz0etf5Lu
7PaPilyOP0p3pmAotfHaPsC5pNuinZGXSgpR0hbveN4ZfmEaBn69+DzSEkIJ/hyTg4CalcKSN08l
8Q/QLlsrGHMpwSbgKp8HLobdXoKoccHuhkZt7rNOQab7SC+2RR6wMx3hG7jF5h+sOnM/PL0tslrq
z+lRtKitvEmpcGUQVvx3jmU8Gf4a3O2LxbHAC6LBIMUp7jORNDUcJ8swru+9BnqYyts1/L5npXMd
i4CDx80EoSUwOTYDbOkZfIJOoFLG6CmcsUEOcea9Yub8mlBC3hpPeXwFppHUvFGZezSgPrqv4uxi
IFpHFr1opLNWE6N0dXMPRceusPttaJmPlfp7ehQQEXOLPVRbDyVS4DhOS3hYcEmhu5mCaik/SfUP
OcnxrfRkLE2A3RqVp8VCKa7/XQcAvOuFN7B6H+qDrI7Y3wBa20HgcShVMmvEwFv27XzTHT7UN5H9
+t0ekca9ZcJtdTPNjI4chOarxvNrQb9KSeW8h9PkCgCwXGan+p1s5PoqvcbxVgX3pxlRAYJrgQPv
gO9sn5V3UjGCBG6mPhUbmYRTQ8kQVRktSRfJgKEcryaeEBnjJ8BKXH/gTeRo966+vfVZ2Wy3jmSD
Tc9YGlHazjW+zZL4YW8pJri/cG/Yiyk7rNea/Ka/JiDWEHc12n1YvzUwKAXMBXtpkFjNbY5ZvlNL
dqboSel2XINYl4Yv/+lxe5wRLvChZMxhFwBUvH19mVRtQGdjTEfEmx8tQwvF4uL03qM1v6qJ6Fjs
IJJoTpzs0NKHZqPEDBV9Tu/NjcTuIhBqKm3mvbxfgV5bvRN4CQhGXDY8dr3quOuFhxVgWbI+qj36
4KEHXonq7ih0b+ddf4OKf57ApbguuTeBYBep2djK3EcYVxBj/sE6XjcH8BMHM5wzWR3c9qXatpfw
Ah8mr0cmyYf7OeyuDFeTCC1vIpLz3ZN5GFJclyf3lXr/iUxIaOaQH4XVgZfiJjpf1zyzvHxPfsgU
KS0a5P23KOwtVrxBrQ8lQi9cYymwocb11f3ADHiv8hc6zCKFlstaGIH9PAWP9PQrOiZzYOy2nhIY
eEsTCYnRS7aF4jQDzApo4tl72a1tw40nZLvwrsK5pmSOMSAVl1cxHWmPWiqoLom2L3mZX21AqGo1
6UpQ3ylpLNRDt2RiGqUwyXVCm61Xem8vvhDOqMNoVdpbIg74Eotx4r9HWGRWZG6mCwgC3g1fEhBl
KX/t42IZzoYZdnr4t9M7U+z9ngCzd6/bjtjdHZ8OcezIpebXezaTJi2YFWKqVdJHIbbEKfS/fdEP
NYQoPgNy3Jrq5qBYQNu+Okif/xKCsafsOp8pXMPegM9nFkSZgq2+9gpjTeadNT5JcXZExaD7hWtL
PvTy0IO8HcLn3brDaRCrtYE4Kh/FTlCtLS8lUt48SOhBMP2NOBp05HQp8+rFpeiWa5IK70ylEn1x
f3zyf4Dopt93EVuQTHXDuXYVz8sFisEE0aklPbwvRj4HtjTdAFk7kc0dARTjFJzD8r7mceKdjmBj
6DrpPVJKp92MqTvIQ3nTBwjJ6nfpRDMOlUs2/BsJuGWgGO1Ija97s3V0Jwtry2JNDcx2kV9HxLbc
g6QosSFqlU4W5uPGAMTGf9i3z/8OPRnlphnaTTv1LFpg9c4K8em4E3E8zYKMVXizrcx1nvDEWLrX
5ngCuQQ1LMLRL7h6BDv0J+F39HZWyD8MT/7ex6mbCllG18EDOV98Gvf36iiUM/LFi3saFXQuOpBx
mhfeHTMtazrjjQ5JJ6usTW+XczpbF08uJi1zcIyHpCUM4ZmPTurdvtXoTRpvfjLnvU8I/tWJ7/eo
JddEVw0C71QS3JyyLoDKCuJaXfo4yGbZZijIwbq/lR5m+Mf2TVmRFcmpEaKu9dNit7Gnp4PN+foj
hjAw0Sb50kXWCWsRWmHu4u0N9BJQIIVq1/IVABKk9SJSjzNxiZWGMlxyuSTy7hO7j2nXuOoQdpLw
ZaaC2pLpQGkRo7ghIRvgYsSfCOONXMb/1ubky1KLgq/KxLELN+SDb1a3h9ppK/B45zQy5/4pWPP1
JZi2HL948nRAqPKpR4MnEWXMxuSeVwX1Bo4O6gsdv8y3/sezcQI9yC6PBjOELpCmq9KOFJ8FB0qb
GW3MBnE+E+DV8aLydwywwm8gJ3z04rECh8AwGopOOelC/DCvJyAaWK0MDD/J30vBqzHp2XVVmQt5
2N5sdOg6kvSbg/xwowEzeqX3ZqTc8HPATszFSh+gLVMWEAOLTuo5zatA7/wPF3hDgK+56XMIxDLa
CGASC5R443SD0UJdXNclBSJR3xxblFG1kZN9wfBjogcbymqJ8FODKxHwB7w+8EcJer8kTxyeG80d
U8HHnHkX/SrYIx4mIfPUPLdmioMwIjNP5wYBcW3/WSNF3rXid74saqmecCuw6uKn1jyydD+Zqy2J
6z5zgtYktI3jueeWVLMGhXik08YIM59ylJcleTAFD2McVa7IvvOsouOKLW/Zebk5PIgyVkUg+Gry
zoRnhtiEmbT3q7RCT25xuaaJeDrVSeOzD5qST3RfCXVNd9nLdiFCSk7DcaDlp1FWNdxlkRXKiBA2
2kJBZTNEpyQLfuddxW403OH+DT6ldGUoizNFc+mztHtpghLPO9Gxz8CUlCOTaGxadN5wkKhU0Og8
nclFAtbg3C0Blpb2l7mkYbZCFoYGZ2LzGo9jP3Cmtj+HKhEtlk+0B6nkYeNJ0HVQY5S+jUfqG0YB
g7WlMaTByYziJlEFFHh4KhXg7jvBU+srgA8uzh3drRxMlRYCDKMo4YgajXxDk4Z/fNCvij5potPx
GLwPxLobmgEnz3lWogfAFGRFLeKNt/zthnrK5p335AQmAGeArW33bwxUoIXMhuuxvViHpzwlhgMJ
5tDOuBui1iZZuNWp2eBh/fsZv8AvX+YzS6MZtDX9O1Vt8efQxIUAFuJ0paTBlmtVGI11HwV5eNeV
j2XXi6/POqUMyiytptbBJgcbSC1DSQsY9AcDnVgOVuCAOC0iHyXUZNuunRGDXBANP4JFDenh99qL
IurSQrLpr+oswFdbDbmn1LgoDbkjePTXo5hbUNhL711Q0sXevU2mlUp3/v+tGvesRDtY5ccB5mNH
qNMvXxUpP3otlH5p0ixYIEHeMcUMpPUmNwfRPSvz+9lNtek3PVdYVZpyUsROxrGjv6SAksr5zYey
aF9TAqm7Kcjqf3Oh0dh7Q935jS2fjMQUk+ie+/PGGCsIryAyXhIEgyj3nu369JDPgv23vr/JGwRj
+MrXuzStMb3+vvGIdNA//ypaRQ2mo7O2nRcQIUsuuq89fYhjkpMXIIPnf4cVcEiQUyeCaUZi0XLy
AH8/eZ9rRkT5Ev42im07NMWXaBKNAHmNsa7ZD4pozJmvKwLS2inm3xNDvCz529hjlf3x/vXHyIKa
n4X8ti6iHXbEVH9fQbIfIbxhu3tOQFvR7wniwSoCXRYVrkfXOYJWxtcK4ZIeq7J6SO5sA11Hz8pL
6ydgWX/9ZgVzuyS7RMtzSmxe9GWRsK1CLuNfDYlx21ksbj/U/VKjw2c6d/byU1jEKVDDKdhdJSbA
Y44rcu9Y0TkcZ+xOFcWAzQZckbpKWrO7HTptBZcQgtc9UM+T7/NljjMjFv+WLBR0v5nDDQmRus4w
tgPPRVUNRJrlnOttbS2PoavV2vgAQpwR81YllWyIu8yv6DyN5Mr/L/sVmLfAIKswsAQf4Km8GkYh
IzZm1cw2QtGdLWs2/BUPNA9urKT2N2z3oO4bvoEsnl+p1PM0X5RY7Y+ALa00ICyNIXzvEhoWlWN+
PSkb+bWunI5/eNjorOlicYMd+gcvgoNApRqvmN2vSzlothAvmSufmuw01SFMu2aXSCBbONjmzCvV
3th4Fg//bT+4U3zZF/CTVHKQL/7GuNHLci/sHi4vKeIGtlfOy2OP/8+bDP0bl/eAzwxp/0Tu1POM
Fvhp97nStiPnhZL0VFcaSsCabVIoC1/kjnf/vBpyrCm1OKaq3J4puWumxr7GItsuWnZ1o50RWsDD
5H/ytBLXkcjgljUWynUPq1In3oG+HFQQG1L1UMrlsXGE1+96JSLozihj61JHLtoPmRWI8WwzLZfq
mB/d96umQKpEZstfm/3ZCgixuu0fRFwV12oYpfKAcqbm4qHvM1LfGVk3JqBxJYtIraJXWvpDlQcB
aQSR4kThDANH/7E/5YTfr0h+CemhqSjaMUAVu8Pwld9EIYdyZ6UCyxqyultA7eglCRXrSUyHnG7m
0pF8xMssdX+ruuRxHpnSdHxrqGsu30119xkPoCPj4/+Dtyj+GnUH42XV2vZl4iZAPUOzq09inHES
a6qpS6dUie5iz/r5BA2+LAmalN3oSgieB4RdG4hTCo4/JbYrXWVMKQUlS29v3q7Q6IseuGzrXBo1
h/E5H0rTvKoGtcPz/+c1cii0ozRAMDq0uvImSncgm+k4o640DvjMTHHQoEjJsU2OJgYQ2r0XC2/4
MbkLN29pCD9PstSMDc4CcOqm69r7gomPL9/NkSn+G3WGxwC1V1rNgRQ3MjAhHfqNayXbDo4yC3fS
cnh8KN6tii2b3NmONdsLGXPbBE9QT9q4+Ny2P3LYeNDs0sogBFmltjfb52LW1qVhXU8xxWLtgmyg
npMRceYYpsLp2zSF2YJipyYRgRX14pD7IqR/48f3eGawBqFaUj0JnDjrFnkSNuW+a23uS9IUQA5C
z7oBme5mKg6QOycKBykCZjoDQf3jArpbIf1iPXx6s5CCtZ9MnhzhMhnFiQlIvJtoQpVHCytLQr/S
5KXQ3vEaXKS8IumK/xqYzxcF6BtfJhYhlkvelDHJAHhtuA87sPtiMpcGTYjwPNA8NFINYdB5itb4
H7v8JkB6LLNW0Wp0ONlXpFJSo5SL7AapFuXIIiJBClNo1PYhxlAUGAwwa0DNUH35eO4DjZZ6qaK9
OCppfXM9eSL4HwNiyNez4eyF0ylv9SUBq/2+FyKQbGV/9PqnBaapNYiOmrFbfaCijR0FbldVVumS
tEbuJk9ARqYpOM12f8FCK7SSk8L095Iw0XKK7GMeq7n0TPI4UwnnkdVSkXuMsxNtSHtyjtNKJC2X
+AfdOH621JGJdYZMtp7atkCBZ/7SXE8Ad2nZ29c9kCcYYq3pgt2Q3Xw2RmD7nDq0p1M93XzYso66
CJzwpU2JAI5P//o9jeIKCCedpfHgct5my6TM3tANuT464qNqMwJfrjBIi0TtBnVxKQKg8wCnyrMO
XSL4Jc1+c/r2jjm5WwGzhenME0miqPvAt0pM9yjjRMCq/RIu/EcQeWHXEA53GjxDIX6ulsm5WnOt
fj/JurBAbz+f3wcN9kjD/rCmGUqlBIHXKo4JOuBx3aYmNu+gH57T24NJdbfSoA9/tud71IhHq1DH
ovTKcLj7qn24M2MqKXTBTj8hXicxJW1At1rW1e0ACTU5Hfs03qSXtxHTk/Msa0yE6fuszpeTPxPR
rQF/SVY5RkQNxCLgzP54Yns5Csxb2mKD1aPLpsSlig2Pz1xiod/h4VD3GbQGKpHXuDtFz9nwp4XN
qotYCxD30oDY+2o58z/uHzyw1VlTw+QeqrGyWPjRoTVK6ry8icG1eW6VdWZGPbsIG+i2QMwBQmot
W+nFaWdVC38cFY59OQIXokinAUHpyovZnTn4j/Xr/DBIMWlFP3p1uyos3d6qeQSOmDrIVNjf4S6U
qNlMe/N9WS0oCOKpV7IE2//bLBYdM2WuZCt8PEkagTrYvKdw0ZRmCleuHDESxsYSXh13JT5F7ds+
UN+jVpGIp4ej2WCN16VAgIhVkmeydPZDIeAWXL9Z3TKpxlr8nYpkDlXG29L9eBUO51Oj/pHMtu36
SPn71XpjzFDXWufgmQs5bgMMOYyzKJynM628axRMdcBLhYUlxGZEza5Qf40lJKtA72paRHJFm7mY
tC8Uu2Qk1emk78kdwMwyfw5tC+ZVxhxfpbIwyQfQixNxTxNs1dYhSv0dCA/MtZgdLUHIP7W1FtjN
Zo3i/5+q8rVo0qSeEZWuxJttyO8iiuoAlW2kTY6i3M9T7EVfHvdpp2FLBMBMi5OC7uu8Cl4x3AFB
rK1qxcwFgUIwjaOG9Te/PVG1EYRgCHu1UcIkjVfuCBPuvrAuEDus7TBYlwKSGjscTNbgOjshdBAV
587RPadOPxhmFgByPGiVFhOYjA8W2nq67pLd4uA4ccRXznterbKzcBeD0SAL7FfRvXqI9c31lyg2
E+fDyzg+PQRhEg7IQ/Egt5qBTH6Gs36BampQJpmllAWSQu5pxoLF2+O9l8n6aFbXqjQBjkSQH6lR
nOBmnh3m/YZWEntyrK2zXYjMALF5iOpVtu9na/2LaAAg9lr6tAISAbd0/gIIT7rRKMGrMrw2/r6S
1uqDLYPfmUF8k88CDo9wmDUQAG+A6W3+Ik6xOGEwporumWFH/+9GMJmelAwWfRVf/zf9/WHfFpM9
a3OVTw1SlLyJlb/k14dbnKIXw1WKSblJ7UQERc9ILIJg9TECEOm0sZ77TLm+YnHwYDrfYZB0I3zh
z4XFmNeaZa9rDVBUG+3IgpUTK8AkHpQiZ9MXHEobBE+//zYAelsoIalVgrOrqWzGZyak/a7xgAZC
ErpPHiYGCmkx9povAzHll7KExeEX7z4jnsinV1iNHXXog+Zu0ddsx5HbLxWF4lbIwijMihV38uKq
bS3VrYhn0GAsubA7BYMb5W4GbJ1gJZCXsT8hrEHiJT5FFaPXhBHGf/uya6XUEys3hmAwQJFe341Y
fLwVu4l+qDL2NUS8D/hlD2QQ/LFAjN19/xYZZg1DlW9WkIzjs11Z3N4bTf1sOh4+VtNtMW4adhKp
PF6J+BDH6J0dkLFZCeOp7n0PTcxP3gfnjUhF/3jx7ikLo4rNCPig3gZcJBFKIihQ7lMRKK0qvgfC
51sOqYhLRleIh8Q4tS5rf5sS4diZ+LxhTf870woC8sz5XfAM1iYkjiRGn4UsrzOK4pzYRT5IZK5j
oyuH6clV60t06AobyxQUXw1yhVVzZi6V7MWD8UgVNH8jRmbF9xseiDDEgoOLJg7TokPE/3MXodTi
ARPFvgTKpWubdVlF93DB7QFIo9EBlUfHDGN0x47XzfGRGEX9g7Ia9i4rnPS/nVPmjvxGWCyts+j0
HG+KtvlKz+cNw2lUquBbl9Clq3irj4qcdR3iYxkMex0xTg4O8vZEUuoqzZl7almQJehWdgBKgARA
+TN37DaSR1ERfdgT8wc7EwuVAtM3KjLNB+Fx51gn8TdASjy1cvdK1vhrKeAChb67cscNo1pUkySw
hKMaZW3VaVotbZ+9f5P8nP9P5DFqPhhoS5dKDQgeEevPtiuzYw2M2dK17hwAUnp0Qre+gknhePYC
ZLxQiS1BPAr2RkkrGdtPaBZKBKgNueEDe6Pe9INtM4jyndcLalTj89eeZf8TLYUPGJMGAH7j+6V1
0Ikg+aFpaV5+TlGaRRBnPk/w6MtAMG5C66LI7V9WMCm6ATeIVTxChLGoGYXFE0eohanmq3VCZcgi
XTcC0TtNe9SgEuqSmIsYVnWFRA+6RPNWxjYEVy3GQmc0O6+bPlrqKsysOG8N4pKHYAOb2T98LlRv
c6tDwVpmJiAHBn6xjXyslZ7Nz8jmaZje/yN51AEhpNc25cYK2frEJcfOpxvV1SZu1fxyr6Kyks0u
QHvF18CJAgGdPqAvrbQ20uEWiS4SP6MwPY2Hp4C7P5QwwfnkfiDYJVlyeZxfOl4YX+rCb+xEJ0JF
eDbTVKXuEQsb2qq0PiOyUpa4RI2yvzCOBPLSOAw2c5sQVuHnclNzONadNXBYp+A36NW5vVh1MUW9
O6fczBa3FBRhP9Id+IJFjGbs/Ay2aJ+0L9ID38tIgH/o+DwboUqZpdsl4IR2ykQmrRfw2Hdjo1XI
sEolPyzG/mcKhAt7O711Ih6EZcQYJShtvyA5k/mqJ6ImeJhDLVolbgvoa+lEUbHiib++cchSx7iH
bSIoE5lSserwTwUTy5ws+LT1Jz1BZBQCsD4/+DI4i7fajIHf8Fk7KvvfF/Z92odj1h/vumhW6R6r
jzk8WBN7fBuiagwN0qwhLERXhf/UYaF5REsN//3MpoUul/ahp7JHlEWjKh5eC1RwBlv03+3cCg6/
8WMXN1YSNYHcpiLN8ypEMgkGjAvncz++nzgloOZrq1XOyZaB4v+H+ZPJ3cih5LIaYtFxhUC01rLO
JcIDePG8vGUFLNFrAySgtFvvammjbKrJPgpz9YMFe53GKgCqUPz5eAdyK837kI+Ml7Z6dMf9wUoo
fTc27KfTiPJp+yCIbUWZ+BeVBF8SIyiht9+eGZmGftnqfAR4DuH2XQg/kyhdqM6ZAnvxL3dVYXgV
QGwdnCdIIeYHOwa+A2WUqAWyGBMaJ2eivo6N9NQsWJmWaklc4IhyjPdOjafbVO7BMNnsVnj71ODr
zs4DP0CfGDOowAV97PKj/SH/gLEupjgJ+LqJ59H9cW8NREG9FICB+TPJMp4K/VSis7MIg/Upk2sb
ng7Xa/bLcPy4uBh26NLdmRleIAFq9/mnYWoReUT94ZTyhevTP2gze1EaCB7n1XeFyDbcezcwXd5c
WReV4Zz9NeEh4gp2YOY2ANTzykJzc1wmjuAcjSlwX41DZQDrOy3oXa0rFmAAhVwKTHfflxvfoI0B
Rtj/f4yJZQzS93x5ArteGeUkWcWKqGoEHkscsz3SNSJk+KYbFDLKYM9Zh9OveVoJXE0aIRpeV0s9
0RBWz82QBVDbPf1OEwmbgsnV3oqapr6gOINfZKYEp2CXRxmfb2N7Wt2JoYhxeNeSVGDN8BpBbRdO
zlh1esi7/MyWuktZ5/OZOeiTLBwP2/+HTN+ZQtvE2KjoDsVBRye/xbEbbtahIt5f4Fe8WMHDGGkK
QmiWFRE/WBHzyis/5DyXaMnlbkPJCc9Juz4qVWnP9O3SWArMHVHJz/3Sk2rqcoYaL5hdk4z0UynM
p64GTZKFAFPtwnP7dIVUqAYPjueID4+FGbLNCNIScp+JQwvzWzQjk/tcwA8Kp+bS451TPOM5SoBN
sh3Bj8K1q5xHHcziyotUExEJlQyLr4x8b9vTjsfhPOnmOZty5l6d3gyFbbJdDkUhyBZkr45qJ4eu
vrjrv6mgfe/RPrg4hD1QsCJIQovD0diaYR4wu+zd9w8upRhHVsFvpmJuvX8Ak1jQUs4U1L8xYD2m
23QNY0idGxY7atgDFJrp3ar5qRUOonI+7CvoeJZt/c9+n5olL7/U/8E4XDWkkqOc84jb1vZiTtfA
Za7bI8e/QhbtFHdO+bmmWpc71S+l41UPNpBtmDpIZSnFfwhBMoZUtLdvAKpICfyZxLyoHf5uO7Jy
UkQu5lXXOzMGWwL8xdplLakZpv0EsLNfosF5uGW+aecy64sud0+lQDDIH3T7pDi4T23ksNhAMPzn
vmES+l8htqzXyy+vJB8qoQe03COekFc0vfmoRsbXxr72G7AUUdLiB7gEbfJXFej9Fr4gp597rew1
u3rmhpx25yKozdamrgIKvSphRx++5LEsFNpacq66kTSEikmCmnk8gymIOV0Z0Pj8/S8OttaZvPQ0
SheLs6vFS53aMm/yTCX9dERL4lursL0X2GFSlD9rNqNTamPNXMT0fDiGz4A06N/rmrZlecrV5val
ljFav/Hk5GqUA+UdqGwTUDNpkwVugys52SpOdTWFuBoHWtddh16VEmXmp6AyCIR1OhP92yuiCxvW
Cwa6lTEB7Ul/n54zRsmkPmECr0dV1bbjkVOY3U7b72WnDYmwkPgvZZVS8qvmnzmjRwIJ65n+VJJa
m28rcPbiW2jZnu1fMpUMSfioaD25Q5dTykfUoZVkQkasn7rsQpQbhdUJjq+Lm+lbc8pIeHgoUFzw
RSKntsnINU78OUcabCXtXtosBLOQsU3D0IfMi5Gm5bNrSYkhIfYfDSRYAxtMdvKoTt2xkUTeUnBR
TKCDGXxZa7LFvWbaK03pGUsR2DqUB6T3g+OgXrMN5phUgyhJnKXUklSOih+SYRQTXLhP7s8XJASg
8hkPjeK8LSceev+TNZK8WaacLjlxq5hEn1+jr0hFeVzpfO4MBcBhRtsEIOAKLJOn1UwYvC9Qr5kS
+bZ2uzvUM/aEz+3ps/TXwIjJdEQA0tS8dXyN1OcG4vm9SAhsch7CvB1Zd0QzrLhVDHq4RpuJOZEB
/t8tnXzIxESv6sKrpuijHIgUaam5ZDag6BdCrlFIw7j7IZPV6soqHgzHXYU3mt1NEtWBlwGQOZfX
H/17UW0tn5H4zvo/+hPxrhVj23k5IGNCj/v37XkvJ5s+x476iAqYEi65oB72rxie25TLrhXKA0qD
+Qw9iag+qpS42CAukfI570eENF1lRwiOTyvZFAzZ60nkGdz7vvR/5bZZ5UTtmOehqyFs7HKcOqiQ
94IjbfTmNN6A4rrgX5KSe8aRVWATpq9OPItk2uvR3EcYKxsmLak/T29umvGuuZMGW/5fJaQBEkeL
F1mPtR8iANDXY16Pojcr/xPo8Z/Zwcg5Zvl2bwO9qdd2dq4ISkwwLyLJsft6yfbPdW3s5p8nwsr0
7a0CDl4KIY7OioGGGjDFHeTG/lYP8jZLEqr3WjTD0CsTpZS1rHA1Gyzm6tIDSsWe4934fXN3X0a9
o1+ZHmmS+VYhZ11fhuIT4beC0lkJJB0LZM7epJ5fb7mGU1gvgpqS84V5q7K3oSBp7jpHtqp6PnaA
L6lZBFCq6lGe6woV5UoIa8Loqu4rglkvW3bm10VswFmbPiBNAOH2Jb7ZFlWb2LrpzzlHqHNhKNnA
NyiXmshhsijbpLP7j1o5hCxdGVvdnuNggHwrnNxuJc5miKI+PU2Jxl6GSUGkQMRNSLLGez1GqFrp
0JC1bZm75zMuTHIXZA0p4+E6uKQoHt7AFYeUUKyJMowoJH8FqbxsGJ6ZWgP7KJ3bX6A/10p/F9q/
Ke4FmQP0Hu8x6xxuMxtvsUPac3nTFdQ0EwQUQuFKrdXVq9vl4XK+A8ltkLhHWPb5ttjrgyuLODIJ
Rtzw9z8eBsb9GzpiwiTB+lrB9PAafXIpJmlKlRJEWD9H+4Auel/2gCfr/99cBQ5JVwFckhuEnMlE
njL+SHkogGOu5gT5viej5l6+FGi/Dolw8GJSMtJNdHft1TVm5oTkMQfKPaXLtDhXPsF/TLdImuDR
b+oUx7XBFm08ZgpRtQIV7krfBgLUGs7Sv0xJ+8EVXOSTeaOgWjgeTzCijv1j+Bsg5wEk9HO1Hr+m
XAHFZtzMKhQ0OtQiJKlbhdAQ0eLHhdxePvZ8sL9TYgxLQs+O8Rzyiewj/1pclFFDXkWGydlzTL8P
xcJ5CQiubHxsUtNNlNlYdmtAjihNKgHeul74r6I0WT6jscS31sXDM/cJaWJH8ThgWmZC8Kr0Zhn+
uiRCTKNL0dP2ll9e6gxX2ZUPbn5HLug/Y8zJyTgy2HmOuD4H3KaJIP11H8kdOT6fSe/zHijd6k4f
pHbcMt/xVUPuvh5bydco0GECiLhvtpNgrAFN9iCamZq1AqJehfhi47uQZKmP7lHLD+SfN7NvPVTn
swPJivIlPTeT3mjDr/L6RBzLysmshqMTNjJF982HQAHfbU7zOUZg9mOjj+/oy0UWd1Yd+N7GT8hJ
ece2apdtJ3atq5ToU4lk/52bj4QBQ+XtAKL824XKAnafPj6r3xHPRVp2L7zX0e8xyAxDKnTFbFkd
jCbAbZeisEq+YJhPm4Q8ax3CbdpRX8OyQTXHyO0pbyOpC3s2BSRuj+xa/x11Qp4fGThO4Wr3q9Xa
zvd7P4e2ygookPfzf8ikIqpl6EH37RIAKghY+VrLUjgvEZJEnacMgCpX8DSxwK5VOEC4qzpINYYu
5/qbymwO+05rY3rfCWHPtFCVo1JXzS5cuWDo8smLmCvMqIQe7HB2wHl26w5QbKRf8kng29mdVZjz
tV4LZQ0WYF6mQ9HHdE5M99b1V7dj90jAI07+1/qbNEqMil7fDZujojKy5XgwGB9OQT8LwTHe3Wid
zMm9fKSIyGou2z5NRso4fwLW01OWZAlUs5DBZF3wLT4ZLryYa4WQuLkBxoFgINe56d2iKg6fSMac
A8DBmP8qSY8vu7jxlnuurLddsW5AbLEmqwZiR+3aX0oqs8HemlNI5nMAzaO8eKBIhLboYVJB7AG0
mqAmfH15Ju3jAHlgJYvVfWnDdTSvqI5KwuVQUACvbTPOIlsg2kG9WE/OVPfwUIdWQHPUA+e5Dw7R
2AsCtAp/CSbCh6s0Dcuh7wYJ3zCbXV7MSzVQQg59DoeJUq9m8ycMLhIRlQ5u0YCwyFskiNIYobca
R93/K01hlGyqJFox3Rux2EU/yi+UDa2CI8Yfcfm63aJFBT9sa68xetYbOANW6XQ7cH3f6bNsEKoc
zkp3LYBeGrmGoPYbVFJ+52JZK8EcXYjT1h/1zfnlBQ8OZYYGt6ZmWDcf6nplk9waTriwQHNIrP0T
EeWBU6q3d7l4PP19OoBrBx6b6aXYoSyJZGU4bQa3BzHn7FYuVv4eGW/r/A2AUjzoTahhdm6SjEfe
ajY862Rn1kbpBblr7J/la6aLHbVhkZ4z3XRFr3ng0stQICPoIIFTS5TQTSSS2pIa7r/ky7E5SvVq
FWx/N1c2g7WjkIsCS/kXyihJGn1Ia2Frxj0dozdStN/rui1AsxqJ9JZSSJvSlKVYqRQE1h17LG2s
Mht/7oMv22WPV+bo51dC3Rc2VqY+Rrn/i+2HcNjzPY//aLXt/o6nhKuKUx22t1w6FQcfHVotbvCj
uoOjFgCtyh7du+5H5LRajTEuPEj1UdYXQq+iIlWLPl0ATpsEVXodWn+UW0r80vM61dHsNDbH/2Fk
aNZBFlxK/l1OlkustNbWfrvxUKxsdDKxyJbjT/aQiT8zyJAaAtcXDkzFDj5qxIbTzY6cktrUobM0
pIkEhfUpe1x4RNR+yqpMnzDesa13Lmdefj4PZ8HxH/Y10yc2E2iqQ/+TCZ5wQcMFkPC2Ur0JXzyR
YljHsWEknTtf7DVPYxGIMARHryb/mGgy86FcKjXIG/CRypTcpwBe9QPjITFm4MWJQ97U2kxdXD5O
kxwIacGT4uM9S8u0Kv/hRKNBhBAvWnyqptGZ8XBC8SMoNDXWrf4qF8zyxqziMoeqzDL96/K6RnCQ
7jldI6cHB1VwnQOGj7azDXH+CTPfj26qS3LFGqtRSmya/h4TR4omoiWrhhNFOptC+/aaa4sj8Zzf
SmyoTUne1Kg7kpdJOFtwWppMlv3Ik7+os4wB4qANAQ3kIz5HiS0xsLUf/H663h+1RvWAj8gc6hJQ
B/vGznS4opIDMxQZY1ZQyY8nJFtscqAuz2lkWd+YTNX3yAw9MdO7AWdQ6iHjfchTRl8jx4qusjOp
8nTFdMyhQ4SRWe4hSE6EroP4+S0yVh3L4cVDklmwrpuucvKKdNuE3emP9/d8tswbrRgCV93nN7ar
J92FCDYAVo20NQELlZotai0/CzgnFDpxQXLbbdmju/6BGVx0XQktkWVA4xiGUh8n2Hicvw6ri0bi
8SGEX5I+gxx48usQsr4cxuNBlZ6bis5nh/fjyz3MLKf9t/f7vkyI/94zmjff49MJecs7lTfId5Ie
dPEbeIo1W641SBDt83+AtXGqWSKqifoTxhm2cUKTvk069WMhTTFwt0YtPlYt6wEEljEuvBoSlx0t
sJdIvZyRnUNLyuZ9NPAJcgQYm16PkbQ431EKP0GJcZZi+gedfIbw+cNBsH9sB2788M2b2YoVKwEV
e6NjT69r7yczCu8sxVHe0mT5XOhQCbPTycxyTtl2C6LDbMIfYrhXBHkzu7xsPtlskns77+JzpX37
07ptL36fz9Zo6zWh6m+mx+8NMNH8KYJDtt8HFtDQkG5rJAjP5Gt/ospVqwLS2KeT5rXkQqERnu2x
dGzSQj075y1vdQ7sVPPuwSupFd7S0JpZz1Y3WeafIW7puF7LHHiX8JENipSUWvRHRKgMT9p6SLm1
HxnMmYpS4Hdt6dQ3Cd9PQ9v7slArRRXhX/GdRpbKOPKpz1BSPpL5szlNKt+B62Xg8J9Ev7zDDbBe
4N9ICVjcC5xANeurx9G8RKUyVpgvuXSs8N/lDrCmu96FlcOzerougkFSiR2EgYF5t7+FcQzHanyL
S+oVTZ22z3iMUz5I2Oifgo5hLaNEZ6GtwGZOTnexkaQ5rvBrfkSARhbl0KXw1kw50BDFda4/6iXj
I5sV40R+hLmSNa8jvPK+dbeYXeHValK5Xh9OvD2y9e27q4VLf24MbvtNeaUCS8FZTKsyEsquTtrm
6yQz4f/VyJv+PYTmJnLznS/KDGO84t6IkX5qYaoFd7YryvXVuMx4qwPjHJ7oji6SQI82Z8vJIYrw
8EIkJCKznUkwmaZBdQQpO9K1kvBE00TousMYoU7qzP0FS5MtEW/1VRG9hPttJJToKo0RWugzXpyK
Dk3+HUEEUTaDnKjkO51pUY3Dpp1/tet1N9J7xoPp2PnGp0oHXDfmPoIyITV8zXkHo14Anjy9uMWM
lXxWeOf2dtEriQEzThcxKCrP1iabmHtpChOxCnaEbJGNosOApAsGZffWjngEBYYKWfry1l33Tsq1
l9jEAxdEpgB9I9Bs+WvNhMwmIvYkcnI8Jz7WkFvGx3Xgt0jCgEi2dGS7Pv07Z5NCWNHXSoXViQjk
qRkbIlf28lsYiluHHjrue9Abe/aIhuIWaaPDYmk2gNcLas7miFmlWcdBk2oPhpx1MzeW/ChEmW9y
YkbSU72Nfb+d5Uc+i6gUIS+2JNUqIY6kVvV2t3h/p6Yc5kHaxSPfHI4XjV4qYOLRSpNEm957LskW
AF2wEP0v8DYV1K0pVZDYZI3hYGEq5QsCUREpsYUJ98xLNUjKsD7ed/3jPMt8XgNreZx6bx40z0cC
6VZOJ6xoypy97JxW/Eq6n1vG3sKMEIhpDuBpmjswBza5KSnZXBBnZj/fnHjz2024unWUKE5yB4Or
XaEK92hoVbPWdv3Prk2ybzBRu2F56jpczLvPltzFWPaRVxFWtE2YN8GIIaiOH0fciugYVGScU+Cp
tebPtRJsvtGNXTSgBe6OedkzIk6wCwNrm0d6YdrUXy5OQ5fY+9ztNDhRHtQZdXAL1CbkKJQgD3q1
JeEh4DjaBB9iq03Vw8Q4Q9HAfun2huaBcO8tgpi+iV6jVZ0fwG22j3Pw+SCi/pI/6q7s0owUSxpK
JqZfG51VtnrvuVvAJ7A7u+M8S7Cjv3m6qNVrkpNzv1pGlbFFheG3t4OO2UJtOBI7bdoKDUE0P3WV
zl53wKYzkkbI18aoE5B4TjGk8NQG5hj//Qbsp52gjb91vGai7hzRFL0duZisdSGRsqelQmfXngFZ
nez6f1fIyu/Ow7Fx/U/G2WTI6HfYpEwCvSy2quFXI34Y054hYme4IbdYEY3TuXSjfAzd+77i2BAO
gVS7LgS8y7hRmj7YygR6UZW4jig3dixTbKcekaxupf6POCWC6XVUzP99ESgZFAoM0ye290tbITdx
PN70X8sNHfFe2ZXCL6CYZ87E++D8CKtS9Kbf1EcEN7oi3l39Mudg6OjZOHDvwiALmBmGGAZMVsGE
q3eqNld+WytJNz/56WNiGsVEp2rhA3JR2oTQWFUMdBhxxrAOsnQEiIG6EOHCquoI/rrsnZEVYkI7
x9WDrWA0LZTt71jderuIBaHFER5rONp1ivgam9wm2T7Um3U9smR+CRqYibcPNfFJhXYz+w4YClhu
l+RLKhyr7Vu58dtxuwKIikaPSRx5RMXGrFUSV7votZjrvzLPF63T8VSGH22/INwTx25i2uZciG5L
0kg9+Tqnily2XAsxR2EkupaF/rvU6HXig/bS8lT1immfy732ibHBNBHqKwevRunFmjigLclvK/Ye
r6XvzPBlRdO8T9dRphDWga9KiGOKAo9lLUSJbJ3gEjD+P+DJPMhqXyxB2uilrbi3dq0onkcMtJdj
UTfGOv+XynCcccEcmIlY+UXx4/jCD6hMNEN5owpVqBARN6NAMmGlZC+05CqvtyJGOTTvj/+uOpbj
KhXhICcPknafAQwpnLiPs7E4jOLZPqsxJwrIpK2yHW7/Kyqee7XMhWiJKLOrOBJHmGIXDu+pO3Yd
oDAz2IS0iLr4ekfFwMnnATGtGhWAYJX4ikLnR+sTcveHW/Et8fZEIX43un7nY+rIGNp2/JN4qHGo
oSx+SrtMoe3z4DDuXxH/0r7z2T1eVDZbIGXn4miN7bs929GZeZtMBWglcPcs8nLzujYZHLDoZhvb
LSC075apu4Za+jzoAZR50KbWLN0R5ovJMxE6uPd6BRQUQjUGdgXr4pyY5CrGkPOc7x32E1GySlIK
OmCNKWus1S2SeC6Hb9n9UiL3T7M3cRinFRlX9LDBV7F8QubQaCQfEhQK24ND/ykVJWqXemuXufWq
fNs8+suNVfODSVMwkclcizJh6QariDwR03XctFaH4wVdtAY+FGw204kVY0xp0XKiOwIBOHt4dOGd
O07rLCMsU9rBdywBQbcG7+XKvu1b1EOgDC3VNwptDKSS595mLOg3sjT7m213/IjTj2GzvAMQjx+6
ttvJMbk9JwAN7xEQsdYFtinvYB4TBRraSB/An87B1uHjnzbKykYgy6F9OES8BE8Ggpf6JNmPid3a
JkwqkKf/ye6QQdAtGL0K2wV60zrk4OtPdbOputlAJvR+Ej4v8ZKwwN2oTtYQDEiSvWmUwlKU5kOm
DEID46m7IYaLhqvvNLrwxmw6nYQ1sGWWaHOtgqD3mbt/Oc5v3A7hI8WboiqRZTW1AumUHu1s+Opq
Bm9Wd0td3A524G20gGK2d7EnI8QQxVdcL4K1tvKO0NPFE3q1ZhQO6qCnVJvKDqZY2OJOsEMODjZg
gXO/XFGT1CKO0VIkbebEzqo1XDEECzuyIrLqzsMnw+3602G7yZYXXjtjcu437uYu87Z8FJIlInXj
mYTpHI5JVc+xGsb44wxZ+6fXSeOZv9gSXgyIKTgtw9sCJOxPswDNd6aKC4XmTLmW6T3er3/dnsg/
E0cL9sdq2C2tf0MFb7BqTsoV7+Xu/nEzxYI1I4JOUaDiXcJScuNjYS8jhf4lV84YgguCJ8lC+rsI
v5UwOxo28ag1tl7ShPAkY7Vabzmx21pB0QNj2OJqTSkZZF15fMMEEpqBJFz1MVpmoTWVTNPZd+EH
5ypn7ZnkYOwhjwhFG8iv5oFrMMyDIVDRhhop8wIixQlBOftHedH0lpr2ci7d8XoLYLUJvJRhIQW2
HKBs2sefqonRD0omK36hjzSvMGkJcOeuk0Cnijd4pE32nE2r2u1Ir7WHXrsz1N5gYzbDqe+/eIPX
IoJdRN5tJsGCUnOwFVXwcv3yY//9aghHhCVSQt3QFal+J6TNKAherIG5WdQxo+AGJGI/1Nx+NLEl
xMf2ndxn5a4bHOSVL87nl4ZCYw8fia2Kgi4xk+J5VGbrOMMk0Vy0ZuSyxJMbGT/g+tsPGapjvzJJ
k6rm5/JyQ6hGDPJpcJ5zVUpgfhrSO9+T0ztCkrZCsEUl85Fl60tTXBcgZ2CWONL0bffJMcmMAC61
8Hdj5io/E7A4KbGIH8aMSIidHy5i8xLpCL7hhhzyLqeEGcq1VE/ruqKtmGlp0ydyrrtUQPMCY5sV
lEVxJytflluXxGuh4QhGOXGw4WXs6EhFOST6IRrNftmsJpsJlby6ZSTgQqHN9wo5qNfdomcUpXRN
Hh+JjzpRdwGsX35JDIy65uc2RcRuMLlaOkX+28IZJpbfGU/zrFcao3EwWIDTW3QGki4ey96JYwiU
BDFbabcyOb28/wNO43SYMqnxZZ6D0M2bLsHEP74Sp2oh/ohRWPXU1gYU/u0IYA0SrBYWKAGcTS7H
lzuz9VH4n9BiPIDyHzf6o1b1ozNIlVPRQGDxsYhLRgFiygBOwbF1LTbVEoteWxWYvmFlV5FA5Pw+
mdg1ep3adaFfHvVxxrpvLInoEprNawdUTX/7+eI2LB48j+JKhTgw9nOOSDSxJ8jf1V8RXqkdSjfR
QDDubRD6oZwIG/rjRvSgwzlizEIQ+GAXsBme4eHi7OBTCJX0yx4rUJZXTt/HLNXqig8cTBhMKEb4
0Ed7AMBQrMof7ryNfIsy1K6GbBx2BqNXffCNHpLGz6u6V7QCZdSYsyTNjLZ/Wl1ne44ceCIxFeAT
iNOBMSQYJCpZiHgjG3KbNFGiAvo1pbkOFFuptBJ90keFVQKvPQGYqrL97BM1VHnr1WEUoQ1DgjDS
Rz19uwcbei8DrmBbKvRV771C9Es24DqGQWyJK7KzTPVnP4452gO1631YLCcEvZqpztw6AE1DlblU
x20yM3P6cv/d18sB2tYSWk4WrydGJ8FSUC0uPVddOyjLJLljkn22Kv70mQ4xTBb92CJMeW/v+KZM
B9zmcsuqpSTpzug/GVlKYfjQ1fDzFjcFaQB705oyO1+TiuvFuNpmQXn03zZ5VWyjX3Ecb7NjH91D
Jyw6oISkO8WtgC5JqNkYsGWCFAbdWe7r/L3YW87l59XbjEtqgbt1cmDltv63OJKhzAZttFO5boOz
GvJjobi/dZRyVKsA2MCSrNcfIVBk4HVCabUOHM5ANtBzQl1a6u3OaVzq+aG3nKVLfRhT7CYVrMCs
PlT4OCg7uAhSlbbP2WHvlhTKz0Fp89BnsN8xUcAEeDd5VEP2VZZD8WTB4TQJYa4+EkR6ToBdNS+g
gjffadqRX5nkGAwqaQWagG+8LBmXZXPNLJuqa19Spz6qz6aJ1aafTXuQol7fCAp7teVj8Tsf240D
8Qg7a+Nz3VgQmdsiywS8/zuvA89t0Pxpf/45JlWYx71ML8XWD2dyQicLCygIoDyzpOfMvQbge77U
uXKQ3S/MfWuCzOfLjKS4kCUJcaiNF7lMfsksbEW2yUnk2weg3wYXailE0X+2vnximDy7nvEy82o2
Gfd0tX9Ely7LXqADDtZPKpq1ReqpBUOd5l50eTUd3bBuWtK4eTNN2EckpzuCFoXiLbKjtjmhjUWA
aib4vGtLx4vvm6Haw1WYmfppEwvcRhKbEkkihtSQ0+cPZ5ITUXzcRxdgGWOSMBSTgSeInYCJfVT2
Q8eOZNjgVrFcUHM79Tt/7Ojwjt0tZN2JliWnd/sCKxmCJMlUYbldhQEmyAeOc4uMCOdSh38n+mts
kb6ILraKbc3NKCQoQdzg6OY74rqxKLO+l6xVQMtEhoVN1XL3ndbtyEf2V+Pr/0vq63pW//y106EC
Kzi6iNTM6hCVSWN/XsGF5SGMtZwCf/KxJmw9BogxNjufBzU9P8950g+H0z9pCdrfKWMjsGlrHu3Y
Wo2f5Y+7rVpwg+LvmbRJ4SjLvSNtlesRZLj3v1WO8a4X8GqfzOxZLTZGRIABscovhG7r2ewRjBFK
8QC1Kc4BQ0XpmHDAdaRXtnqd5doX7JsLnq7L0XGaUS456k2n21yVuk58msQxRyatGLurdQUzgqcD
68qxRSCx6f0wvHBmUH+WFbrxCfHnfcYrrF50AQr+/ve85f4pRRMft5FX9F8m7DBwm8iPgtTuZRv9
d+F1Ys0eS6epaowg7A4EvJY/S6p5DMr5tuwHn0F9NhH+3J1tSuOAZJj60idm5RRPVC2W+6TN4Dww
vXjLmLDNw1VSIVmuIFceQaTwncagM73udBTgld/qAX0r2ehDoK/ieGdNtjdH+hPSXT/o/0427WvI
8kIHQ0AHrZqViZ735aZvAswwZ3+Og+EgGLZDGy7dEPDCi4gzNKhtsDCLFfLjhhjTrjjzmvuish0b
WUN3sdVGieEEehwr8QY9MO9+tDXaSm9F5JsuKiP/oj8W2mx8a8kMdoAf9tt0+ar2UhgkOZjPTBrc
+3EgyEVF2wyydVQ2LwOTY+D+AY9bAkMVZ0qq8Kaac5csVwQKRo+W7MwS45S5GcAPc40ZdYPpb9c9
Yku3kBSnZsqaPaAm1CtN2TqkiLIyH4wtoFA4FbAvjLRj6fDrW3FL4O9N6Z37X3qDMUYzeTpE76JJ
hPlWqNnj+z/M+dkelXAiHiUV8l+By/RaqJ/QoD5INWabsw0ZGI4Jfv0tAeUyO5pRy2vY0uUtoJcS
kwgLiICTJEI/wfO4nR+rhLWl3ZU5ENxN8sjMFnRHUekKWyHl4NlFKLY1pr20sZsg5p6zJaTB8CPQ
/iIkl+Zkn/fkvPejWbk54b/eZiOlY0LKIgVu8rYUwfdbgDzUcxmoqq8wDRmlsz4P5t4RP4uTZIQz
hXgVjgL4b8kir0859Z+FdGR9IoapRkKnsVy81n33H8lS0M6Vetb6D2ch+TrO201NGP3V4ZaRB2/W
hM5HCoOoAcA5NqW5/A/cvsMyt/3PmSar55b0jKzsMAlx+eEbzsMoZryhDaBGX1EuABcO7iZnJkx6
e8icWX/bgrCR/wC0AJRYe3g5IdIaOYAEwJio/zZ+4/MUVN4AH0NZXX05EWmmJLpcyPWoEIinSz8c
lu8lowog7atsYU9w4IagRsng++adIckD4fyMpfAXuXUgx/o8mkO2qyptHZhVcCZDFrO7/Ot9+w1P
LhBnQpzVFytnPudBlWcOIQohB5TjhXvuSSHui1CZrpayvP0MytyZNF7q9TpaWqRw+UGXtMr+XIdL
CetGH7PlwC0fyjaWeT45W8hYpGABqoy5Ku0npuFZcln9jIqWctqLuPLm3DBvA1jkKQkHLrRtXylx
2N4GXqBiUNP1OpCGylgl/RH7ceCNEM2jo6ux5Fe0h9m9mZEi6iRQ67W42e00QmPgAgC+dD27UFZm
5FccFt/hzquD3sxlQ8AOTK/AGQFErRhZZOROBv7nmQVta9Bpf6mtooO69zy3CRN4nHoyFSvGm5f0
k7z77cy1shA5EHj4xQVn9BTM9iV8am7kR7JVnSKHIRYbhWdqwONNiszhu3nKFIbnfxEuMmVF8CcT
jJasdXErOU4M4Gr1nNSGlTwbalWsis7HBBTnD3mnQ4uUxdjG5fP2WEndewCW1vEupnRCpgvQpMz1
fXM0lfqeD78diDsxLvEDg3ajpa3swgPquVx6L6fKREohRGBJONLPnre5FzcUlviKhjArlDckPayU
fJgse99TlF3nSCGYR3f6y9nk1ixMg6E6lsbdLFmn5ea9XZlkga1i0gSqCL/jx96VxYBEKSp0HcTP
2GPOYVA1XJ6wqrkRcE99xBld4z3OUGO/GWbO5krbpjKSFYWo4jcsSTeFMxIMwyQRoNVGjbKAwM8i
9mCbGzXrUMZI0ZgdUPkzFhwSstZJoJahEyRkasBAzACbDg/16LXzd0BQXWB7sXZxN4zVuQgacLA7
OHngpDWOaZXppLfqbDIyTOICFE1/6C/ghNOkG3/2b0jjkjyWylmcqcrxq+g3zsm5J4kRh5wi/gQ/
0uPSp87rmdyq6v9DDLWHqA+FT3KBc51I4gvG+M9IdK+PmuR5f7fCQmOfHw6nK8vYKEVaujNHe/Fj
xX5oA9wEYn3Tv2FKyyobD4hbjvVOvXwAFk5EhB7Te0nFjz4e/mjWvB0XZ1otxhBuXQ7EjD0dVpno
Vlu2WSEea+GVO03+cJ/nIGwR2GGHEg6TfCHu+LIhyndB8lUihgtc0dvOac/OdptZPcB7Xep8G8xZ
COqzjnE2I1gkSWzGEdfxAKQPbCUWoLaJMrz5nyvMcKuD13kn6qOmsS7lBKXIIt+LIzLEaXWk84C/
XzQN+RLrq5NAoDNixJBiNmFIh8ccRkhG0PUmkk4UDUeOXlMS/17Uxy0ahV+CUxyDpThr6ewNBjFz
svDSY+BZgKpfyrb6gDqQXj+J2mbUVRA7IAOn5nWKb769YEN4oK0cty0oy56oNGULeC2WWljAxLNT
2L3eZG9cYCicRcaItP8EVSxpt/DRqAsxaCtmQysXV4FndaxjMYO7G+LNFAEH088y81w+KwIx9UTO
0S1vOYileGFE1pvYLLyhFY/by67aqw3ILGEJy7q/8FlfIOUAZLHcS+FfGNVwS2JiIhheWDP3PGxR
3hx6NTTQtx8O17NC4vV7ejHMjdWpUEQTLFobBkV9IyV9T0G8g14+MHxL7sSvbnPzbwiqbek05prB
HLYGOxIKqIb3nC7SGZWjUY6a7VrhRva7QcYmvFwCoPRlnFYjQ0rKJfO02wKtOaws6d7pO5xLZJWw
l/RzUXhaW7LnxozUspByay1SHN1FoI1UjwTLdkYf+OUJ3aSlTSf558QHI6QmwFaenekPpHHv7IAK
btbf3ajAy1H0qMO5Okj+LteuR6KegfkOSMm25pDlF7iK7rK/5AfgMpTFREEs927XbLe98glE70R1
UfNHnCXg2DY0xEp4mZZNfD+Z026TV4aA1Gj2DvqBc0fIgZ8mSBipXAAWp3lxxwrtsaFrfz+u8+So
Or3SSlHABNw1b3Bzcu7myXktqDlQYuAei/wQfm2HYzZ+hVW87fLCvvfA2OmQXeoa0VW/yG74OzyP
E7MAYAgXuNPgGGNux9Bv7lbc8n+36sn+Yy4p1Kq5MWSAVBRox/W2M41hmJlph8bIf1420Yuk7r4N
mm1l0GoykUZFK+Nqw2n0CmJC1AK++ffCBFHEIOoEd1P9biFB3wtTbdmFw8z2DOFKGqwsP+x0degL
uk7CDbLh3QDwiN1d0VE4jXDvgtkGhCnVUjKXa13h691mp1sQFvEGmycS026vG1Orr2Xe8382ezsn
mCxMI40+/2gf5t1C/3eLKQ1vw6HWVot4RTrDqPuO0+wiOh42zob3jdKLlkIBYiB1VP/ulIntL5ol
7uCkXBeXwQGotDv1LVDpGhHTFlbN/SkNTzACmIyddWC2S+lD8MpW4OUlB7vdtnUYrTYsjHRa5fg5
oG8qr72B5OkWLn5xXCIqF6rYAMilXfLGUS6zeFlFHv4mtuqjRi0uZITw6kg3ANKdzTCWa7B3UuoC
57+vaHspZLXfhgGl6GLKMdZIAtqUDDQSdcQHPQePgW88Boo5z598ec70CATcyBhH4V522y/vQr2b
a8tCLCD++p4ICQF+EqoC/rap6ChCn63I1HAiGGbQw/RxVvgvzCgA2y/12M1igYu2sFEkDwnLvk7v
laz+Oid/8yI80Zyp3uQNylh9dnObxMsegp+bNQ91qs+pzRlHI+DD8GiRcieWULl0Ko8Z/Rar5A/F
JBIrxJIbWtvultsC4/Fww36RiUlFv3bMU+q/H7H5DC7vmiVaQM4lEE2Xi9zZp+OS6im4un0y53gh
ji18zBKOuddLm7ITd5IIHJKznllQaGDIF/I8k1hWr9v3b2ywrZycMpmFrhP/s9M4sTXl9n3ZeM04
sMxYhlzUmzwOrz4KiZtH70pf53HJNZv+ulgDfJLZrZZ1NEXrz/N6o10x/+ylZqJkQm0xBbkSWMIB
K6WL92rcMDFK7oasUtxEl6q1nvRkwai72LrM4QU75PLH3zkuiGMUWF3Kcve0AXRymZWSjCZntyI3
L6oCR1PSBDFFKZTD2d8xJkCOhT6O9yrOvAgi4w3zOR24vGrITtjSS6piJxgX0tWFJkZVYRhflq1m
367cJgweuSx2WIP6vWGpYxbGwZBq7CvCNYqO5ptVnVgga93Xn1Qa8UKB2O5uDOcwMF2aQkpfET6X
C3MUaTfNBAeF3/7803qRnq8F/a6Sm9Uok2+Y2JE2XPxqepUSZHW6I9YgN2a+BImPZsLwciUcjylF
7tb7/DsRD5OxPiX7zw4YOL+gjQQOAX8TnggKcSupeYiSrMtkGNJ9/If6s3xwFUmOSiJfOIqtNU8t
pu4dEOgZb41IaNC+08/OEBfDpLsKcXdbkKEwL4YTFvhT1aWSCuHF7OiHqsgiBm7ldViMQVvEhDlk
SEQMxrDyrrrh1LVPzfAkt+S/mB0Nr1d5oJCVv0lLCzGv7B/EbB0jwkCiTjd0HDZDNs4tiy/WZ7vF
S/76A1wwQS6y6OL5OepCddHDR/Wp0wPwZe5wGYyrNRJWC8N81H/tnB6ZE9efaIxJPvOgn5tChNNN
ZWXSvGB9Y1OAnDNjwiM6W0dvhAfkeuhmMYVXtLcZZPCa/C6GPJ43lysuwMWjUxs3T8ckcEm91U2Z
t8YEVNJFcSM9XUfO4RGULFnWitUm7hbyg0VxqHAZe7gM/ZU+WTfyh2w5Bu8UimqLoEwtgB2OkDxZ
AE5tCQIG5XZndvqDRVeWkY3AxLlsHdEY1QKGaQPmSVVFv/OKcihDo7PLPztoQmpRH3bXxrylcNy1
TiSTP78CwxZ2zcVgX1Bn4RZV5+0A/6gKRUqwE7wc8JFpmG6yYdUJMPfNgdkI7VVtl4l1F88mGjq7
4zywDdtO26Rx+xQeG+Q8ORfLS25IZRCZ2NUlDfQcmvwcwVhUO7h6GXG3t0LmZRKXSvJbgYITxU4o
Pfre2Jpv7rTzZ0a2We9twp43xMuRvRzQEJXsZUCP8/FffCFzmdgYcOV/S3GLVwav0jDeAhwDMc67
5VmIP5wf1lRNg4e1YhEFxHiG5s7wjQfLtxEvG6pbgp/QzyLkW6Fxwm3giHHy+RKwoLFVoiLGYvul
VA7yjZ+bFm4vzzziMFzSQsBD1Ecr8kcZ7aFOMQeNxpR3yloNxdfFm9Buci8v1fppx99GdRZ8rXP0
tBRgDQLGUeMDMwRMI4ccoG/U4NT+RQZzCJRdD8N/fdRKsPr0ygWHpdSR7hqgadZSIQfJLFiPpt8n
wMrUBfAGs72vJ/UTWoUiXpKOJRvRzhmDMy8+yTAz2pY731Dho7+iKWzKOhT7buuHkWp6R358fFMb
J7yrBvG7GEzVidW1Uw0v+3kpO9oC+nBudeB3rKbFfUQPsBR75SYzPurlu1HrO+Z5g1Eix0nvLvbi
RtKRvStk/lNYAhZdbeWnIlxCdjkrDIEoQu6aXZKgNfI7dxf6hz8d7iK3fTN9c8rxUIrYs8abUM/i
jpRmEQvTvvK33gL9G/mZgbNlbrBR1E7GP6C+4h3WRgLuQFt4qHdkl628yHEyOHmyntgXEu9chYbv
U0Jkqs6R0jgkWcilDTk1S/i4jAWqA5LPLqwgf9STREnQxCfrWxUlOHUjaC0EewrYB8SpqLOAF/eu
OYAFdj4NuNj3ObQSfd2lPgLEsUlOmKf+ow7sCRdzVwLHRBK8i4Y/KGgewHb42EoqPZ6nsRF8Zc0L
ORuq26KV9SuGASzQWJJl8+qmRdz9ZMUI7yYTABnH93d7bzxVElcYlUgg5jz2yckROB+CDUPHZbqH
HiOaWN8XUndnPCpMkvCM1i8tVmgpmUG0b+rwlm4RGFMUJdAm5/0RDWvjRxl4U/bvYzjh8IFJjYeq
hPO0MDx94fnZIXllWycxT3bAOOn1IbTVp6Ja8u2WFuV9siwjUbSxT0KCUGCpwgMJgeDvFDhtJhNd
bE7U8kK8oUaRbQWPMoz0AHdAtSmePnDJq1Wch4boVJVK04FEqvRVdF8zBeQq867123WSs3ntJETR
qi6FwRqs5DwVMgE9/2kImmwu3uqiPPm8hOzMgwOhxRw3YiGj5lFRA3fIblocuCQ67os/7OYZWWJ2
68JMFpfUH3PoXIboUMUsG/hbu5b/1eoDkIUgDQQEDo1amyUvmULQQUPH+2eqyD2UE0+ihMMS1cCY
+oEtGG6wwD1/S4+177AZdzW/GPt1q0v/89cpJ3I+rdyJMjtidDqR1svzFPFX9FyZmdqZmH58fzLy
8pwFtroGK8sSC+yIzCl29laZrSz4x32d5pVuOhYZd5+qMNxCae6gjCAF/TemWA48Qkulhmy0LZOu
CCUgj8HkzgdoSjWsaGHd6dbhPHStFcVi40FBk12PpJvv76EEO5kxtiafH5ophNHSBn+uL00781qP
5H1zdqydIGKlEiOjFtsUyTdLwDLjJkzqJ5EREgo88thcsmQN20ujUdkY8DYlJAVf5iuGObsh2JLA
7PykymLPz9065ESl+s2+UVox6zK54L1tw+4j10GUss32XJFQdBI5Fa5siGu3cnRFxc0DyC8CxjRq
BuSzUy4ECPw7JaA2blQJItzKXfbf5ATuaEhm9wWX48rrSl4HVkyH3jA0ZT/9Qe42xHPSlb4+4VLy
O40Q+gjoCGJyazikuUzKAYJdC4SRbLhhs+7Tf6RAMO40HMnRzafKUjyqeq1tJTSru0PxwHF6lruO
wcoASs2buaI4mbcEhIkZcA1YIdi6yIr1WEglxICKAxluk0Ecrg7ngXDtMTpjNIEGXG+UVDInOLW5
iHzUXH/BvzHI3pMzblVr6SlnvEwHz3J52ifAvbrIpjnqNg91JtLj+Ph1PJoPi6fS+izjOhiblcaq
1gbfUP8fSMm6/cjZUG2Nnn1wfKs+i0Bqqce3h0HdEEnL6a1ZQh12gPDGwmHq0o3WBcgPYGzPLicB
YrzG9E+NxZIp6EQucfbZhGCqJYoMIagqUZ1AtDRp9OLgizJmZqpqLlIZjHo/GTZLSTIHxw2NTsF8
ssLRWpzLxTVzAHPJNjW2bgR8fl7zY5vaGpwvn/Xx7aC9PyjIhCILSjymL7crMkGqfpCui5OYznFA
mltTbOQOAUznkY07Fy17MHh1cuIef6cwJatEGON/fUStVDImnJovuh4MCNfYwZSjyvkWJYyBaO68
DiKpXRmIt246x8JPc49zkonFYIIWTCOqsmnM9J52O2/04XQyjiCQ83zZmXrwsE1XIpxwooBRuMF8
iZdOJ+Ybu4yacRCNbKO2dFb9DbQxzic/vtUxYgaLIKRf94/M+vwGE9b+ZIopnq2SmRbn08KXsdeI
4dS2PLO1OYAwOYuwqR49hZGWyVCVmvHACJZMeAd1a/RNfY1Q129xWV7wvjYSWZ+yZ1Xj4di/3BfJ
2PTfklKwiHxVUctfSAmfdSDr7iYYzxWml/a+5uDW53Q0Hzba9oNmZA4bBwsxV8in0IqbbRisjd2G
77faT+z/tS2l8gs+o7Rd/t7TmkTSAlyZCsKLxGs+yNvZyBWWXlU5IaUXG1vb639FW/on4RhAf5L0
jaKuKtSOtNyOG84eDv2s1HTwP+KYY//Yyri211coCKPqd4yKZGcD5c2fIQBXNgjlhv2bwSrdFJir
/hZ3KH7AHK3h2u3y7CmMhuDUwmrcdSgGt02u9pxl8oLMZATN3TzTZLqd0Ay9Afm7JSXYgGP7A+ok
rxkRLwjPZAfYC92JZDwbsegY6y6saoOCxhE8n+zvvs2gHs81l8TvNg9wp2IuasqxunWDtr/HhL+r
6O6QRT5PRwkBZ5jzx379OPACH4Z2qpH0OXv2kC93FpkHNykGs6Qkxx2vnNHAOqE6zIARv3I7Eka4
wJLXllBd+ERVaitclREf5VxKZmkZZhxv3U/bg0Wm4BV7ypjEYAzf/kvg0Kfcd1jV7uVo8uF/PnQB
0Ny42eK8yMr9zp4Ij4eJs8svfiu9xZUK8cuWCWNBdoTrFyeCb0eTv4mJYtzwYu89hngU9Re6KFjN
j2F1ywhmapwT8GhnzIxDQ9Nizdg+QbVUfwJbsZ4herq7F8QJI9SnXoCcPab9tYAeIxbaBj1tIDPm
Fx5BaH1yMBUiLiPUYm89seyIkKpsK2lwdUVL7TFZKmfBGtrQ0EteMM83SWbEYAXHtTRpoFFDpbGh
4LdA31OcRbHGT6GXFwZ7W2wtnejR9qOW1zpKjIw54pi3w5DnB1T4++/1WBH4Otj+K8poAfu5Jro8
MBABb54jfPne9ahx4ZmreOegxdCfHZBsFhFJnc7mvYIyGCeqbpkrXAOxAsIEBX0Sagelsyuesab8
3E2v2T0PPEROLqrPD04uT50o5C5c9gGtBzQVhALAIJlgqZrM9jZuCM1cGoATZ4Vmuy4I2EmMDnDI
KrPWFeUbfR3+MH3iGmnE8+gRQrFQoYM++xwTar+KLq1MULmCwePuMfgP3PdP0wyveDJ+4MiBlLWy
wYTdSKxf48vEFAlQx8sE+CkCC5BRSbaWpiX2bJE5vlqbxj38YA0YwxaiZB3kKL1RJ1zXbDtYc/le
NzmprhZ8Gt9APCTXTFv5tGG1LngDurNGneUTDRnCi35fcBt6btnCZSLgYtCrER8VWwFgffslz9qe
KctwryKmR+XDTwXz3bmVNgexO2GoGrFuX+VUFDvX/sdLEzI2WMYYLEEbnzsb5dwl6EGRhMWzWlNu
7dZik9F0rejeInNZjDKr0wtPiYb1cPUclDjdIY6UTNh5zW/xRKQLVDQ9rjefti7Gxk39iehi8VdO
LrJaboxJfBgf7ZR5+p+qpzuRhFMyeYm+SQWMDMhjCVpeSdGPR8rSiDGfqdC46vVABJ4I8qb0kLI0
ITpbPnj1kIw++aE5loeEd6p9EiZd+06qhB+MuuGRB3LLTh5j8PqISmdVragu+cE7+c2qNVp9TFJQ
KLtY20bqBhfGWgRqx00/Ufd5VNrvmnrSLlzGsycwOM/Ybu0+zwKhQRboBoh6qM8Vi0bEF49Oo4Vu
OfjneAabaKKYWU3ElhcpwHmxeggsjqM2Uz974vX6fJIopRgSOzQ1dXUPPoEJg7wCstnMmHlKOG9b
03SmyHGVTaPUyUssVwC+ZGrYqhECH7eep8v6+Rq5UqvVL17OFlYCUpGYRdTmDiUFnOpuLvuuWIMO
HbAlUkg5e1cssgiDVE0jrJjsB5D50tQGOWCbPfM3bNwZ+rsmsTU1QuQebSP3VAC4pdX61DdrM5Pz
z9rlJs2aqHvS4GGecSHIJplxK4vUXTLyzfPWNFzgBw7Rhp24wxs6pkriaZjmBVYueeRI++v/tGkc
+9Cw/Ic0UOcuhpX7j6jbnLu7/ySNlk90tO19W+W1NxiWJGI0NkOwrtvFSNG68SESkcnX0D+1NahP
xWhvkcpDBWX1dX+82fSM7b9dLoggmtHKBbHKexr/R1X9kVyTmFH9YnX4P3c9LqnqXdmc1VYro+0i
5awrdcpZWhAnAta/m2ketWIA8yPrYgoVu4AIYYkW8a5KgYCpPkRyI6Aq61o4PByW2iD+ERlsd50/
LUWXU9aXPAcVcHh7DTUCdxfUqn5Tqm2I6nDAkm+E/si0yNwjDQFzLAAuf6FiUkI5ZlkVu2VJ9SM9
TGffqMiUZxFXQg2EQohFHZXMXj8OMQLdqF/XRhjhqFYUhGAzsGbw8RX76SWi613FSuRAFBD1A5Wn
l3Cdrc3kDrUymOl9omHYjTooUpJTjHOZt2HtCOED8Ef6i4imh3kvkyw6ygt/RwAx+3K79sPey9vD
wZLoCiVx1fuun4DqawQnGDO+a1XhPMAzai4wwjD8kNL4fu44MXmmZ5TE5/7xxmfO+yWsvdyl6y4Z
/WNN4DppzHOsODXmhIkbwD3HCOfQ4EjR5C9brI97ESRqfeqaNFUanfMnBj3LgkQ5j2bwkvmJgNhp
KfipYoIsxsl5EFlD6i1LZY68wT0Yme8qNcxCDq9fBPwrHqKidWfZ/ClzH7/5wt2+6M3eCIZkDYVy
lZPJEwhv5ZO1hLby5hdDJFNoThKb9CB3ouaThJXTPiewc8Yt8R1q8RT1BcWU6FZVDnUEGLp5L6ZK
GV7iMyImyGkRNJ0hcTOrUsOkFH3NpKF4PGmTd9O7ZOr/Ure0gJDezCLfzC+WapsrCkkfqKpZuBcK
hPFiI8dTtjGM//Ms24p+E9l7j+WM1BxRN/kdLdxxKoavpX4Z24TKQQaZPPYefxbR+x2Do7IQQZQ4
grwsWFSA0Fexf/mnQWbyZn+8iwCiOPsF12oMlLUWKll9gEZ+aNE+Bm/YuHRSR9eHgustT4HmUl34
ltlecCWB+DpbdXuJ1X/pZ7xrESNNTYmI67H6ihdBrbcUzV0JvUyWJB+i2GDmjzcirvrTfMI35H7S
jBul8+K2kdctqKL4+U29IHl2f6rwaBfp2NHUOYtEM5IrD/gPsIG0L1jRipnJ8mXJQ9X7j0K/CI1j
a3ZqfV+KScPfX4zO9LsBQcb1hftGS5Fc4ctH8vpIE0fNtR+NXGJh2XuHLnmD+MYH2Jx6oK3Npzaj
RphMm9T6rCkbjZrEsFkljDBJxoAyPwvEz790TLtZ07txmxCqVq308PwEvkoBj3rj4a4g2JZBLhDn
hc47DMmBU/VgMpEq+hijqu2cR1LmKLkhLLnqLhNo4ULBlRxhs6FQ7gJlaq38GIjtFxcAWgDDVSWg
TJHAcqC7Hz3aik3XAFuHE0UhVdkDXtz8B6j6NmKQ0PcMRWCugJUgGFcHldA0FLhbKl6zDzuevdq2
vmsa62tf5i6WfiJF4CsW6gDYPWDnSclXm1pxjNroPVLW2/v0yWmm2dw9Ewga/phc7ZNKVR5N247K
KlMVABF7mNzapDZdGoPIPGRbOH4JbDB8KLGeu8njLInLDBLFOKMG2wmENs3FRIj4AY8omnWmJTpy
EnCAHR0kqbJuMg6IQe0rILxcONEIr71Q5OFGK0YgzJqMNxnwPzfz34AjF0u0y/B6bMxVwz5BbJf1
qOcb7Y8c6JMU2T6Ywv3QpQ41rIvlFmC3TL4i8opUScYDozqfH2EUAMqxtXVwQUVb7n+0Qwvc+OjB
e3KfzILKPy1lNtgckQtwlvoWIu3NS/6I4yXBvQMAxVf659vshGYma4XTaDbXwNi52IDvp4p56WOO
mbM6fEvnz6TIUjGf+Vm69dWczcBitgbFMDDMPoqdlIxLg2xCT5YG4ucQUXBqOn5xibO0LIWrl9pm
mUprmwHzB2o/Bkjz3+p85qWPPGH9PhUeCAUmk/fTlaX8902llYDTlKTtbpJsoO+3AZ2jbjWWjsh5
cUPJ6iNNjIIQvGrglHmMze3niUahEHlNHwlQmQBVI66WJ+nGo1X8hegyb/3Ap6AMCHSdubHZS//d
v/1gWJFSCDOGdiUrTBo3VOb2l2eVTFw7kaXnSIy2bENdTUOIzcJA7OyOJIF1bbifjrxhWQb4iJtx
N06hiVc8ntlwUfeofOCCyKtNjHGHWz+xCBxJFaVUuM8Q1cCe4ODpdmMMqvjIe/XEyfdQJFSFt0Mi
YUpxxzHn8AlfyiRKZ8HS2BhrM1Nv0AJ2S3pXo/OmjXYM5jwHwqymUQ5LGtt5CvYwEVnbO01A88NC
XifPV20plM7KcHVFw3KCohwYxV2fzWS2AFZQ328+MhKj7QyeNcoh72R6zoGg2gSOuZl3xgVxlvt0
1629/F3ULqfYn+1M1rnzst3TOGlR+3h19Wx+Q5QS+YrHNQQXhJ7CF4sajxKlnIF6BrXuXsV4kxPj
FUc7XivfNUU6cxZSHlL2ckQWbL2zrjl6QI2x7p0BX019GMS+PrXWYi5mn1YDDQPavPnFj7kM2WoJ
BIr1F3P2MN9DHccVHWakzscVqGxOME7ZcoOk/p9CdfzZ29v4KsA01IgjdL0ciZCYQIxV26s3B1z/
ata7007WKDGS+mug3j+0KqvP9OQHy9TSIXW3Uv2C6+BQ/MpKYp89hvP9C61ApWzwtIwFjo39AVz4
GY8rGnADlfnR2F8cJF+JyPJYLS1m1OnzhD/dNFRAgW+MAsUiyQIXGEOwm6rtJbo5woBeegv/O8Ue
Gcfovi4OVD1SIjirpitV2DaQKxvtt6XK6o7b/ufecNoRNc9Q029jxuOvuR28p79ahMe+smWx0Iw5
/1uuGKqlBigWdtVyTv/hsoAos/FIVyI2s37E0duVldAiTXeP/L42k7GntrPbTbMLK+y/4p/Q74MD
ocVeX1zbj49n9OM758f938LPdLVISY530OgaDnIeISkJTT9w8uUAr2oUeQF7Mm/XKnz7tZNIXyHb
WSdf0GrANRNXsKRwwnmdvddS0arssq8sfs/k92FDz6cI88HiO9ju40+ejJQHAersMQo88ytzabW0
qD8T6sQCtkfUo+GiW+QVFBBddEZHEkz6w27XFkxjYU3CwH0BryIUacOS5NAMVVveHPhmINOIrX4f
0tiVAGf+vKg9+YbA6d7qmiYxAzHNXSVL5LYchevVhBgT2OsyEt3UBINXSjKa1L9JI/TpTQpGLYKr
eU0pj+AOSnZTA83KE1sMJhTCLnCxtxYNyMhkICOkB0C6lJ/Fh+IfjyY8WeGw72y92crA+G2dmMe5
dr/Kwaa4hConhlaU5w7AB48wpz8vsQI1Ro/ntI4c76+AdVzK4mbYMwh0XtZ7bMB4sbCqtBAshXJX
KS4/EoTK4xbLxxkCvo+5LvIATMNZwLnujyHQr31ozWdMc+gvUThTstkft7xPmYk7zi5LETvXLQ6I
ykFK9ydQC4Od0e/7SfFpTLoqdJKUc3DoAYw9Nc5Uwv6aC0h2vCZeVgd76AQBn9ir4s+LCGftE31K
UFEefCnZwCwbCnnXCsYEnqXSG/UsUGutcTDD3MtKEpnet09HAne4H1zVSqVz6FCXTeNvHyuoGQox
7/1KFGjJu3ylC63y1cvDrtJNF1Cc+p9rVWjD7f6ItCE24DZc8XzoMHKGKMCIWpnGNtHn6jTLz6aG
nSRpMay7kNF0Ht2CfRBjzzVB/45aKsZQ3zmTxEj3VXh3wXJqJR0EVazpf4zdQ51wXdWua6yxe3vr
tmyqfvxSuMKufVNMrm7+aqPYPy4Cq9j0fbp5rxP1NxpT4Qrx8XG1his7/K7b23rzro4G+gHzYC10
7qZ7EUjUd9T6KU5wy8nFGjbgjfmCB3EC8RDr1eWwVT+yZRjMUfzG3iB0GvkJpw8/BWRZ5GdVACd0
vL1h17hj5CiFar1hlkPWGKsXPZeBZsQZp1dyNq3mtuIic3X3yn2ea599ny5UU6K0wE2M4im5Uh1k
b/f6ap31FNSUf6W2ztnBEBxF83K9g6ME5wugLaGT6pxGXUIpdQtcbqWqOQreFD/y+NtaK0y4ksFi
+wRrQumhi5CwqcJNvYTZh+pwN3OFAsicVjvw7Q+/OVBhssLI4K+gbj0Gem8dTwaLISwJlLX9g6d3
CHUQqbkRmlYv8OhLI3twhby+PKFRcFjrWxanJ1MLvW5fW8RdAnMrgGXb+tOwEdLXusX3gMnqBVqD
/ZW9aOByAa+M9vFvgHNPuRHWtqB/gKCSfQiTWHkdmzHe9GH6CEcP0DM751gGzqHbVou/7OWFL1N8
DmM4Z3vKorXrzyyN/zyvKESidBvZoORKnpSibRa7QqtXsCyeBuoaop3kD7s9SpY97+g9xWn/eeP9
ZyfOezQLTaUfMz+uZgldpcGwTUlykPUodr2U9kUODQjn4x3TeKwQROXwT4STZyAnNT2dLspi2Xpy
zlLROgPkw3lEfa25Lc/6pt9I5yXL2dJBAVLe7nCThuA+9wSZ+bZB8gg5w3RMQ+zn/qRIC1iW2IHL
Z5KdVydc6SwwR/RXjTXgHpho4pRMSMjbSB5X1mXd/ysTr7vlQGap2HLFfIuOTPr4lnPyId8cV1+9
N8imhrablNZTlxGcFg5D2szRjhZz/uIbUIJrRddHh/3d0HawW0AgGB5yqbpXlu9XfzpADaLlASOq
2q1twt9P+e19bmqfHUMphACxqkrBA/dfEyJoFI3qk6soqAtZq9qqBiCjUAuBGCo5AREUgDuNWShG
FY4xjH4b7SWtucFZFCbFKgXJiLwCRGkGuib8eK2GGC15klCoo3fmJFymD4w8KTE7xuZAtFh8mBNH
zvR86T6YZg2zPACQOmpUUb9DJCq3ElcwT8AK9MP/gFMqi2z4HsmkNN5Yz/W6cPPya0w7L3jW1yFh
UiFCvA67KayPnWthtmu/mqJ6DKAhPeonTFNHCUwxiawrv0EreKi4m4ofMqy2wa/e1dRPSjaSv0b2
SSkJSjDUGKeEX/POC9NrwH6u+5MKxfJxiy/tCDKu/3+j6L7WxBQKwYIRgFBYQlWxeSKTd5UTvR1m
bqLGrIaSmfVNuSHzb0TSRLL/nHzmIYsIUr4rR0Eu2Fc5fB5YF4crlJ8JxGIeVRfgwznQiYsvS9O6
vFSAy0QTxUOYbH6y2xu3y6tT3vOUSyO2Awlp0C5C70mUI3pOSN1ZvHmScYR7/szHhp9sMzS6PulG
QI2aYMezNMCmeLFdnItY2QkdEd/au4XHm3PhSTl0RSU7rSHwA9DY8VK9MFtdP1jDCsve+GiWkJeb
r71KmR52BUdloRYnjeXKMC8IPZEbxVKbbEa93QWrwntehdEBVzmO90AXX+qEV2TF35f9J8j99dcT
DkUNPWoHfGgOWB/4sBXMcFNAxCpUhCP6sCs/n4FRPsnzYOf4j4KLjHX88W2dIoWttmvOx+t+I10W
bDWW681S12aA3nh3wkiQaB/dQJXCpykHHTjaPv/mUsI1OEg9I7FHC2MVo5rrxlz6VRfkz1x9gc9X
GkAqazz24hSrLhPDeMmauLaFdYP6iGJG+4wLaqa/v4HfCSQr7Z29iFWquKxpZddgLEYR5nmJ7rMf
9y/A2BYlGH7e9ceBYlSgDVqeSqg7685W4NvF4nxC7J4m6s9poZPXwbbP7MfNdazNiqN/E6IPcp66
/TxRpYm8VD0gHhxy9cK+Orx+koQsEqXqAo0fJe0X42ThYhbB5TDW5qFRp1SBBx1KdYJ4x8/Je6wH
Hv95DsIqg5syiLYM3ZSqNsmaby6yVvfO1PPEU7F7U4NwKroqUmn4q8wngBV1UzoiAEyBRFnTiXAT
pC8bwyNgH4D6sjaxddoDodPU2w5I4kaQoOYXRTxhYz8I2XABqzMDate6tKwdluqS+Glf2MJuI9+R
tXKRhA78c/M2k3B8zaTaeBrFySQRMza4gBHi8KQSrmUZNj8kayAgjRQRAKTePsmXW2x3GkIRJcQt
FqvDpLyFhOdMcnNBhbS5MP6rbj6q6OcyDYhr681PpN32vrYkekdwElagLR0EjJEXvGflME2YIAJJ
aS9ncJeMAJ74Ayf2GcrLn6l+bGK/f22R+UsxnMeYbUjOZzcbRk817MPdEjNxWTPtM4A0itMaP7Bh
uhpco13uLDvBpe9z8h/bPmPhrsZq00oZqUngphxfiEAXfjtH1eAkmH/+dL/N9wfnuBF6um1uF//u
Aa8rCyCqiz35p5ejvsBeLRx38tTEN/Nd/1zkGzsSr6EyXpnOKCx7M236klC0Pks+EiTTcF1hQ4wR
5ZxPk7ZffoqwoZk8+vcz/qREMku4eRFVs5OoDWfFHibXudGPIs2M8Mi8JhQH0pGsW9wBshWZfYQL
X0diTc/Ql7uJ5ieB/7ng/f3HFZqKMZ+F2RlbN++3WJGflkUd4fLRIj4LL0gAdp09uGB/jwTYdAna
ITFvNN8jFiIMu6WcuOILjVqRIgsKZRVaVyWTJk37kVHt1uOOjCXiCBR67UsT/xbN+d+PQGD+jf3W
vgS8Kr33hvgo/pIwdp+B5yV8ZcqanK/4zIlwAfiISTW1XCsCsD7haQ6a/X7HMYwVAgE9m285s8IP
30OddSYLLBfEn67ws0muYYisAm9ENmSlQCjfkL+OZJonnMM918asD9srmYMNvT4vLHJxRpFaL+Fy
B8BWbjr5Ntw58BG2Je/E+71lVh87AbFL1qZW4WwhzT6uyiusjkqptaTdEd4NES7u1g5fgZffAfwX
D8ONhWNjffFhVCC/DHujSlmSZifw4ElA56GfBBA6gK4LD150Ts28eiDCJfZ23vN7VU0zZ8UNP6sA
t1xCz9pBow30qiJk1Pksf90UOQpjWOJX4kM2r44tkUsochjsVhQGdyqdYLaf2ihO1ft/jdVfT47h
BML0plxkoxi1p95Eysy3a+Jc3N7cYrV29JP9jR7B/HvzLyVM5sq8uXyjVqO/2K632Ql53lALY5CF
vJlhTwrh/tS7g17aSy13oTqCIJWBupwZgd517MEcNnDL3wpn+C1CGAR4rmlHMoywXg1iL/ooIyot
qks6sB2ev0oG50g9HRja6nHWfDVnHOA9yOAiD9keLd0Z7o4k5ADWKE7bbL8+7IC3yPw+p8K0dTan
PSOTvc/+Bw9hluMoCNR01HuQv4O0CaOOm49RzW9B9SfUngdgY8cPLoypxGU24Y4lTsLdxeG9QsxX
vLizUSfR0hyjIckFt6STFrrvqlyMos5HcDjsXFMGYefVczTEAvuCIvL7X1AK680HHo+bUlci7sLK
gPkjRDLbCt51Gam/y5aPuu8HP8EvlpWlj5pKvHjw0ANP5FvfpHM6wSfh+8tf0D3ZdTsZfDXiG73n
GFvo1ZJrINP/VqSkEzF4O1PcgteteGCKOCslLNYu1IfyxacXWof7D8OX1s0J8VQ5L67YcWCwmgaC
TBPbSwVM0Hfs/z8RRBHkqVd4HTyzHmXBGt4UkU8dXYA+a3EniHvzfJbi1WQRLF0wST9c4xlCz4R8
T4O7RrmqB12PuhfmPBjaXUWQl4gKfSuY5PHCNal0JKrzBqm6A/b9MqxQo8d+TT9szpL6EZpejoS5
K9I5J9orZXSryzOXcfy0zfANb7/KISugrdK8lGm8eLauW+ixrLAeaO3VvRtEBn+fFu9KJSCtvm/u
Upir9lBSLbGQGXb8Xr96P3naJTr/ldWySv3a8agKfi3uyk9jH2B8dNcd44u0pVMCInwIvG65VPan
DwPAK3p282zYNUU8rKzopRubyca20+ondB/TPSBPtPOY1+sDfnbuYw+Vubbg6N15irExuzNNWGHV
dekQ65RZCHhYQLmeHXDmyHt/leO97zw/Kqhyak2UBwoXpgrPveuc7iwKIX+FkhnmfflC70IpSadr
uOD1MFbPo9R3kRRFRtIIh4Q2EOy/j9W6HQPnxN9COzZigeBWghZ4fmugZ4MPBtuZoD2wGzQ2nHe0
84WI6TfBSaRtL98C7S2a4u24fvMMQ8+F73DzHeylkAm/0UxlGrf1lfeTL4U/IYbXgF8fpDGapjzI
X+Gug3iP7iw/RJ6JJlboDI5soizK8dPhYnSf+ppf+g6gjUTxzbZmzMP4fWvk7KI8EngqClIl2sg3
fi6HHj3lmS3y3d23r2VVBDzX43g8lCPKR9S63qjZeI0pjMeEldiw+WZhQwuONAMxhy2Uj5nRQQDN
S7/DRJXMJRoWdwBw3eSRSlIl1Fi29MhcGS6qsvGkJYuaWxTZSqZoSmTqvjKVrzAA1/hHTomoNM4B
rmyaZz3p1x1NYbwj/uEaUOrj4pl0ynFefVjf51nWwT43XJXi1eVF4TBN4i8wx948x4YKbuLtAewQ
+CMfhBIdUfdS4/y3rEWxF8hasqUnmON3GvXoi3pgHXWCqoKYfnyEzZ29nz54GDc5ZYrCNGLUcZr/
dG4+3FyCwl+Dxsuy9ZJQ+S3tDX41gnKIumgeTFmlz4/QPyMX3KhZ6Bysk/mXkYYG1kLIPimTehaw
CFzjRgWyYFhC5Mr5bhlhVrbJ+Y1a1CS4kMvFoNvXTrUXLMyGZ1g646oL3Sk3JjIdP9GvVXDChi1j
pLwd4qR/6qU5/OOAc0YT0H2E9Fka86EBSZ3tAqsQ7PGstaoFE0TUGNsobYjILcK3Wz/6OOqw4SZJ
nViQigCskR27bnSQKRNOHuOZH3jqEs4WFrjmg9+BEJFnM4OmLylnxr2KlAt8GXFDlG1+t/K+CUij
WUi+VSMequPXRrAhLd5C0K1XKcy2jE1ojtHQbXaG0ZMTo7yM/GN4dBDFsGYFQz+njB7eaZK23t7p
g33QxXSsummPXceTkTvMbaRfJ1w2qzcboAKaU6iL0avTJGUTtQIc/R0gzBgyJZ9hQYO1oJzbTLHl
jZNmASUzN7QCPU07OJO2M3K4p1P3xGK92385kroJYXrjxc2GQwOkUnEGipqf9k3xwpcmnG57ZYFb
bc0XVOm6mUVgduZHSwOP/Eu8kQ8atvzD+eGzxOf8+xoTbE8kcB3dgfvmDRQWqakCuSvI+TyG8VAn
QX1KMBCfKtAjU2Q5x8fy0opmpnT3ILWkexwjzN6wklfzPLmg7+KgYUVW4R4SQazlnqxMtPyNYHdi
fX7sL9gESlYGprkxvKM24B/rvdbQSHn7LrKK3R2b4jOJg1IKPXAOGC/hAL9FY6tMh7KdEIR/Yccy
TFlVoIxf8KGUvFozqG3EqgxMyDqzoSO635tUyy6Sx5sZL2R8hHeksX+NiCMoYUNKjinxx46VFk0d
nDRJlnxZcdRRMIlV+UJ/o+OvU928HcLg0V3Hn7n63U/iXsFrkMd14w2N59MbzEHKsziEJ3Y1GUOA
QFQ1M55ADI6HcD/g2qWHdMfW8S0bUlAwhvOkAuVqhrDm3Q3pquUFm6PjwDqr3RXswl+BIhZYh3HP
zFsxhbFRnYRKBjLwT7mCdnzA/rNxVj3BbXenac2Rzv7wOjxSC+Abr7XhXprolmePqNLM9Uy3Jfwo
D+l2FlDc5zx9o9cSQ9VLCxM+a/V5P9Fjbc3HzX7biMpl15Bq86AVdhJv4fC7O53jkhCMoJPG+uZd
xqSnnrWKHAaVWNWbKytwVeLYzMqx8iwEvo5d49Qf7fQMUc0tO4JlY8BK40iIKB1O/N4loKCp3HxB
tVJAK+xRKgZLCt+6wXp0orSZbbDI2YlQJJaIn2arPil34xQByypzjsZNq8ltYr+R6K9sy4eI07QE
OhAwlzSgTr4Ope0qNe9EafMQ8jSc2WI7QJXeYDWiPbgLuOzbU87U+6yRogUfuVN89+t5u+JwqyA2
97YVrZScWcGztP7frzUOZ3opjHwo2CvlHHlECzqBEee9EOtxnXN9F8yFnh+Ml83xbJOIRyTsbqyO
+effPSicJs+WOMcwd6ufa2MDvg3uM5ACMvNtQk4aB+ham1Zed9AQMpFD+HvBkr9jzeiVHZ38be4c
rKtx5mq1MMkgKcMrTE32AorWaQdiL3x3T5/3S3ZUNY2wu5+MJjKJnqvMmef/2KVLFZ2lHiGXHpWM
cO9QE1+39iN/O21sf3ed/pPZ2dqfloukKMIr1ewezEdx+2+bqrcoZTPs6UPlGuPBcQJD5I4joP9z
42boDHMHgAFipb/LDcRSEBvnBcvQnx7rmi+kVZGUNqneG6EcuusH0tfES8ZBqOQ4fY1Ta5DFKfhc
LDMZsI+zzjbaeitA81uSDoTL83LScXK+7dKUazxXvN/UwBXQGWXqb7cD8G2qNEP537AvIilfuTp1
kVQSOZewMJtTMY8ICdQn3wd5UrfVjNDkfXtwnwQdGW2E/f+HwPraefREb/qOQ0QvyAIrv8v7H8g2
/GcCDL+6miJgGfY29QUTTgBaJFs0EBozCMAjgSxc+u2s/m7Y6kNVdHlJdwDs3Kv2sCjQJZWvK8K+
aiJ5OCpydpvJeZzLJIAQCPinAXrrBUrSajFJYVKm2di0z2cQzVwu2HhkbYMvaFdGvjcGQ78QjGVU
l6Nn1EnELHcX+nz+DPZon67z4mnLmjs/m92eI9ZWsGXMvMeavovbv9rpOrTubCSgRZWK6xXs4S5n
rBevSa+Ti/SEDxfhTJe/DKIDnGPCL3+YlxGk7SmKJsXfNotsHCrNqAR0JczjJUWDudmHwYaosAYs
flxM5q3Zv9sQiYnbxwwhVs+KhnQ7PVUyhvBRWr99509VHSTPlFdUlPd0XOthC4sB5/9GuhHOwcdT
AsjHAsSjQP/QQH3ZLVfA6jhuN96H272tdx9U/RKO2RhLWiQAhEM6YUtEuc1kUM69YncqmQX/ZUFS
zHRzCHWnVzk5g+n2Onlz7uz9f1I/gvwHeBjj7PTguzn84ySIoRVbYnm018naBgS47PPVz6UKvXa0
7VncgK1iTpW5QtLaE2t/pyHiefN/vwqCMOtXz2jDDe4G1XNn/0erx7qHSaKSN5aMO+BdwVldfftu
NRX8ZMSij5CX3Cz0DUIJxkh7xBex4ujq0Qd9Czyuyr7kOCkM5SFNfFGtHZX9ppv0wqLAa+M+w612
BzxDYj1Um1BFCx1aNBJnjSdNzlUDW0msRmYBcRZWqgBPt9mfdND2Sg+bCOFqfqGq8FId9zx7fMvp
A5C4rSWgV1XOW2rpFiRMxTtSh1A9yOA9IQGrB/c+YnkXUIXjpvOIHqkteGOf5r5AAYtT4uIJrSF/
kXJT3TxVmD2a3K/8M6a2XOId1L6QGjtkepAv6RoKuwYA/n4D+eS4xMtIlN1QwN4ThodM0Cd0COW1
cmGXm/ovuODor9bVGu08H+2SUmO//s4XVJjOD0NqLH2hGEBbJHerIwDViKRUTNwo/LyJU01J10aA
jw3gitf51+iiVN3cvfdGE+85hfclLJPjDV1kq6b7naaj5SLGds1LHNx52zHnIUPv4TsDk8F4t1Z4
GpN7jUI7XDkmjfO+rjAq3iFGvPbBs4AZOLMvzOd5hB46b+wG/808bFxhyQjRx27ebeLf3DzMq349
g18eXh0zqUfBsDyjwEkNVqr901hL52kIugZZGfqm/hB0tdkO3wXS9zCVZN3Ea296rJX+gel805P4
xCSRH01sZxw04GxpsQmsRZZFZPVnhSFj8NfJMul6XBPayJdF1mhu6FYCdLAnFXsv++DeOkrGRjTk
BvssMVJeQDoMHSJob+giggC1Bd8/RGy3GjI9o373Vu50HUHxgKWjTrYLeaVfFCXZ+cP2IysGzfr7
bGQ98FeEXPFz0FrJISNct60JgT+IM70b3p1Xqm7ocHjcBSTNlCr3MQxRwDvqzY0b2t9QOpA2+HMj
CYLpLsyVcZY+mhN4FsUQBX66YSyhFVOM1WOcZ7yh7LQ9cbbEkCGqHV1I2a4XR4qT+mj/6gRIFaYc
VLLILaMC68vT6A9gOa19GEgfftcBIFzDuY7EwAvn51ONDLhzsssLyvop5ejm8IPmYnD0GK4sRy14
BYZahbVargPdpOXi/NcSfa/3qbRESm1YfDMNW2rcUhketsGKgF6+vV1FGGVEDj3DUIeWcaCpIPFF
5H/aVcbV7705LLX6jw5VooeovZh46nieiJu6rfCvZnTxihJPMab5HZsGAzoFw8L4RSuWQoGuAyIX
FgwpU56B5O/QjJGtMtAFqequd7Kx6OFrc1z397gpMcB9sbG2tm1nc/XUaCmsU8baeSo4enm45JES
HHkbHhZvMowzKW7wOcnY7uQ3vlLKFLujFUKRwprq/5VX1W+/HQGoaLq4sB+EUVjDI5T68ZyL3X62
cUbUN4x8HWWxAbui9CJVsjKsqXjiGBaoQ3dvt4ek1nvQfKVCkxqBTRxIHc/10kAxHZhW08q+1DG7
YIZo33NFKNBoxuXWJwDn8gLLExwKxpM3uB7HfYb14vgORtVtQfavFDW0iJ7qHNmPgpVQxQBCaZMh
MTjiHwL2cmYsTIJ71Nhh00V1xPjwuTNU201Io2ErWlGM4PUE0vzuyulDRarwAfeVlvjlZeqhB66E
teIqQtwwUo3ELa1/AhjfyJTr2/hsA031XzFxOGLyz+t47xIEXpXay1yImz/tXGchIvX50c9P73Dj
0dR+5qt2apJ8P1+eqepbwlWuLTkCtKszdjCVMK9cGPQlFBEVpeG3hsvjEIDiAtMhEdVd0oXHvB1i
9DEivhC3fe0/qX9NaU7rl20KMv4jEPiruRSYthVEuCaGvypI8CN1/croa24ThY2okQ5mrEzuszqf
N/J6CdVuczglEqzHKe7f5SXFh77hqaDVj27obXzzqZ0E3ZmgtxsqVF+ZbRTO1YJh2YB0vN6MyfGp
1In6C/8icW+s9tC0RJJI/bvIU31n5VXxtXbBO9Y0Rsi9LMeGwX+LsiYJs58iGtK4RE9RF5dMFryF
3j3gDEc/rGZGDB+a6V5Rg3Jyj1otqA0T2MrUGKHhCsHySslrkctpZE1+YhGO60A5X/mMO7QM06Qr
qiFSV17uun9ZzUp5rgwq2/tkhNvDdLeVCj78ZWfOnc5JnHSSVdF8VWRbTIR1S3Q0Xg29zkUNlxDt
aJdDw2H+nw3wkCKhBmbURn4tloUBXun0mzOetcvw5otoXBdk7oSj+ueHCPd4ouEqThOb38PCqYeb
YUIFTHYNdYHMC6rRS4Uzpq8GEbwuyNUesyMJbn9GYBXY0nClNpXxwBF1wAymY+mqdMTmeris05Uc
HWzkOPksNv6PzuVDo1vqZ6GI7nI7BnqpYebG79O6mhqsMHHzuLYekiXKybq+OD0laSK0kx0urwhL
q3Z0Z7duTR4wGjfqrR7IUQXE7kebOKcEuyQA79h5QyaWdbvQ3QiNwFdwx/+qm6tGqcJwALeOSmVG
eFEqwbQrsJ5XHhjagyfeM4P7vEmuWmoen/PEEenWsDilPqg+OUdGTBDJ0rGWVpaA9+hFoGxm2EQt
haljQ4Qr2iY3CWmi92II0c2SfKPgBQOJmrSa2LtxbbK1O0j+WBTN0V+Eks1/I/Rl4TSzarCJN0QZ
pvazxxwkUrQuSaN0pk5JVv7wVV4fYhPZSB+8b9aUkH4+rJj5g7S0pniGYPA03h5gBGAZifxPhb9X
lOVG7NjredS8A7gEIdwrOY+N7eDQnxgjUycCAUu0DFaweExyNhJ22iQLhgCW3ftSAWy66tKsfGeW
zFsKUXMmde1eYSgWXDslOUj3UHTnb1uOVSLda7wXCgbGdzTouPthD1Z18eJiNa7svMn/df3MOCiB
SvlZ8wKcgFArBjaDCrWQyi2OYvuo5sONmxuAs3Dpb0mT7NlOKxa97WIxtpttNLkzxejdmr0qbbb4
usHu2QGbmYLsXWOODZ8Vi5keJZ0oPW9W80zBMAea1qE2uUdmBS+SKN1JSWBnk43ZyTmz7bSYd853
t4CaqZvnJXYm5q0csgeHKOllc0K1DCGOKMQfJLehLMH0C4l0ibL/d/13aPSqcGyu/m0f9d5vZ6M9
QdrM90GZ60jN50huCprq/fc4rHI52GJ6AySTzd4bWtDfcrh9L6K9G8SFMZP5voMP2MTR62KthMqg
sR+niVbENBuSob+AndOLgA8UbIepjshVWMju/FTwvx+le8dbxb/MBGoFPLxCuDD2n/SDUPVDSY0G
j4v0OWG5v8JDrDWVfi2DF9qTGBXKSkljCGHwScaHW8lXvevUPd1S0LdNFO/hXkSU9K+Q0CLo6NND
KWrbpN4ASCKbF5jJObqQSAcwNyywNr8nwbPjTKt8RhJMNjP9PNxz8MMgOfGaTIx+JIvXxqYPQwdn
hVkS4nW4uTg8z/SbMbGm1w557l2Ckz5+UkGNUhdBHE9LT84gfy/zIKLQdc7JIZzqVL3omiybeWMH
98wPEUYDP6PR3KQmj5tDKX3/WHJ+61upiYrI5PPg3UjgUiPqQuRPEpAqUt+nr1774CkxfRFMcITb
39jxLdpcMVv70kX0aIoag8K+2eDK1EEZpG7CfnxVCkRwoZ4UKdPyycAs3lnQsSuZ9MGmWoeAgVxE
z4pWhlp2yNRA1jk0DTm2ASMCKsG8SHQ9vup6Bec1ha86k/+U7C3PZTpjBONiidD4dF6K1sP1P7/Y
LWJEAzhZbc9FQiyRFm1E4o4m6I1uiEFqSPRzkT5ugN4l+7HIDXZOgWW+RAbDdwLU6e53SOtlzOlP
7AWbs5C+QdIzQnybL8t9RC5OfiN6a2fxaQu8k0pKug+hsFfP13LR2BaDQumf4m3YgZcUdA3i39yZ
9S5q1knnOdBGpKu7VgwZvl1XSE4dx8TZ+eDP/R+ybL99DN5nlvsdnxuIJHpCUo3xdg/ulxLSxUuv
lz8Pd1w+pz6OtDEGLu0J4Sexn0ak0FhV3YzPntEgpU9vi50tLbVysFGrWx0sUFzqKULM7WbqPjbD
4BSBLd32Zoxp/giW62WqOHDoTgYlrVQw3lHJX+MUUldxghSVPzbjhH2hzbxNonrq65blAVTX1jHN
asqKIY80xQ66JsbcfxM6i6bqKOwqhiPkhSBW4qtqaeL6lz5FNZhGjp5cwdUGcL2wVkNxe0NEivW3
D0+L6HxCLNwylywi6CXd3u2GKxKOcg0lVGPhKfipZtXwn1lDMs8a2hE0GhsuxdER5Pgb2fkxKNxJ
FQkq9sqHAH4gUr10v2nkE2Tp8YRt+bLp9ZnF4wAVLrf75YRhq2bxIqXReNXK+JtQ1RXkgcNTKodU
MgM4GKdW1ZpIKKgrz4u0gJcHpan5JE2tnYCjsl1e4EwJGJqNZ6QQJ7205bRwu2nOd9dCp9ew3rCF
OoLJav8J505j8EwaLHmBO2O1iF0TufLZomd8XCdjR8sUBCco63CcbiS7SckTMpMj+jAFV8cIpkQc
NXZtatLBTfKX9ICxMSmuy5NFGrqS+wZW6vI/RUrV/jjYZL2ggzJ+6nDaNJEE3Q9MfHvSeAgLqXyC
YmVb/xOtKhFi8hWpnDeaEjVbaEVgxQaS6oM04cZsFLCmS9l+F71EMP3fLTb3TOZN9cKoqz04JbwD
UxHhpCnmRJEMuzILwxdbxWkbyLPdiC64NriASfQAfcbjAxcmoXaMbM/ihW0MQZDaRlaDD/mN2FvO
kWeARtendBWgO26MEfEeix8ko6IAVZKeq4aNkwnbAJriG34Q9nxvV2Yu6aH/IXfkYF2NDRU/NJYN
qFdmM6UCKVKT0tVBeqWXETXMyd/2N+/XbJuAyT8Dp7OaNDaj9jpTROBHxwTYTFeKAAdI/VTZja1t
3E4dCxhO781bIZoHb/tqBjd0GoShxm1vcQ4BN8BAdKArMh+46i8u9nk15Cm574X4CevpqpRAMhVC
M8hACE94JRTZ+UVnlB+XY2yihPOX2VBN3ZtXR4obY/1jDvM2mcJh6+ZzYjgEzucpqMSlhv58bLy8
fYb0+TSEpuXEYgfjgfjfQHdVS0RyghqlZqCrcwZ5gPV1icz7yHcx5PVM+Xarre9HhtqxJZmfxGWA
iUkZ64a6UhJEV1smbfrfXcU9VTTk/NgwZhwhBeMcy2JK1pxTur4MXbjj9OQdXTB0VlKRgFjuBDQy
gfKbgWU+QbB3k94sx+Uk934fPQtdROsrqhPbR2koy4ljeU72sCb9oHks5yuD070S0/tVjf9U6J5A
nYJUewN+pLytc4x3MMTqp+QL3Wv+7LGNZr1WU8xwC9QZ2RORzaAjmvq8aA1bT9TKXALquwOCmbIa
MtRvpL8eRD6EL+cYypt3enZ4eWDGWQ4FIJjtL1q3kekqc7+XNiDX+tV9j1aJTWYpHjSBj6JIiYYm
+vj8MPoiQ+uH2/ZrPt0gtyjipcBUvEigIdGA4YxqDYz4A3KBjUiPDG6kDGSjCQYHRsRSFI5k1zGK
/RmppiddifJVmZ4qXZP/gwNU9ctTHoVMglPx4lysuJ2UrV3fqTS1dCm21QyFh4TZ/yVjFpmLWIH8
ryaxeQIyVwfID5MXeSZaehE3QRqP1cihHyD3R7n4qwQuhfyD3XMasSCZmXIrYPbg9y5dN317joKv
uQgyzEl738n+Xrf+is1OVYpbjNuXMrmamD2wqpSwR+3/E06+94pw7ZSOEofZu5tp3lxMY+cQADVR
/O3AANUvsG8vc6CnmlgpVMWdWFPU6GQGXwciDwPSXpPSavAhjccidfR4LqbHHMjv5UEU0g3KE6n+
XKFplgGQkp9tXLpIPN925g2gGbSfISS0qkVhHNj7OtyspZtJrTIOXOxNg9wNnSU7ApNLoJz5tP3h
3qqQiMPocw6bKye+hV5E7X5umFShvQvkGQQ8RfbU1I3Wba/TQoUlHDxMTTNfpvJq1cE+0LB12Qb5
NaWlXqvZN6js1q9nJe9DfB6ueVGAXY9IboH2gy/trCHCMWrjwSJiyNQkmcDv15v7sTMRLKooAtVm
acjYVLQnBOseKB3gsfZijU6p7chJ1tjlsHetHR4dlj7+fh8A8Kbxb7/D0b2jWAjNxmod6fClk6rQ
t/AmShOZPpozX9xn08r1psBb3hKPxJl181qNLJv9NmoYQpWCF+FnD33ITa+7ErkbAjAMLd1BfU1p
WBz8v3O/H1EIo8Le6je+ZrL3Kr5cbIRjQ+AVPNvs3BA/2kSGIYi8Af1GFwvY2iaDgEouRWCsqDDv
rEY6FhD0WKlTOgtNpv4NkxYRo09ai9fMIA8Q/4G6qlYGHwdT2PrFoGV3EdfN14pMjhaObP1o7LFe
iZXD2nyVUT5C2bbSKmY4PVWv8nbz4ERaraqVtihv9dAczQ+XGx3ORCHxj6y+2835Mje9Yk1olXzK
CKp4LXbvkhh88WpX2wnWhE9Rrbj4zloYeL/Mc9KF4O9naWDdpn4YYrwTsrpjySYYMFxg622AZdNr
bBqXDRh6JTOHMmb4G0N9paacf62h404grRSoPYRko/UONJKVU/mpua7wFwRPIQVZf3sZSGopZKUU
0azL4ujiEJlGTZNYHWvQSwcIxvHP1SPi/bQknWiGAGep54I+GZ4rz0ygwwoTnRZTUl5HOQ5diJDe
upufCB613dfpEzbsCWZ91k1QKWKrsbe485MqZa3XhJ4P+GvPtph9S6FZvXJjmcTKJMuDrL+JOcwA
noXNfGOptsFggr2npENIdXVZyFK5kLQmxAP52O41B/YpctOIQN5T7d5y4U9FQzDk5CZeA6IZeljA
H4rq+aufAVKVt5AJNOrbsG0LtCtiGwEIixfsaGcUnMJrVlegohiv8czjEBVyz7z7EgDBEbqlNTzS
igwTeNVShGlxB4R6nlJjjWR/lYi6cmgKOW4IvKCYypHykWXTTfuKZ7+J7N8GIND15iGyi1qLweKV
9MOOX0KEdGeTmPZBXg3vfmzco36oIWNBxRhrQ4FGrKzV+IkEM+iyQOKuNu5qRz3ZACjBbjQkg/Tv
+H13I4k7s76eiJO2ROso2HBIHyoyMD04QoAQVgJeoO0AmSdTgmY0bKyErv0lqXh9erjX69yZRdIl
wiF4M14iAeKITu8uIZi9JzU25OYfWmP0Lgi4+znhklvoCJt0SVucEgtRJdfqfLfzcrcD4iX24SUm
uTQKZsvQjn4F+EJx6D464I1pTnmVs/fC6Rlbr8wGPK2jIolWBslq0dd2f1P16bk10+im8+LW8FAC
iQeDmSvTTi5YsUJQ+mWQJd9O7uJCRzIq5bhp5k7x7ep7GYr5Hc5GFnM62LRoM8hdX+Tm6KUNgTPI
EUNNsKuZdWKHVCAt1vPg+xdcjdiRuC552m5Z/pbS8+q5HHLWBLrN4NERrOjA/k2d9BnKf13FLIY7
vn1kUMBuijb9wUOusfWEDbhC7DDNdMsPiZ2rpbm6IBbyFa/xUqHB8BSqvJNHlWHqpMlmZW20G3Cn
epK9YMnn+yLEHS5OdW2hh1+7xl4YDxMsq9kv2HzC1bKEus0Kk2BkBY4w7LcF+u1nxbvsRc26XfCj
JC4TWfPIAO7yROYkYkqF4YJolhMJSPpxKVDDoyaAuRUUn4iEAa1aoa83U2qzo9xWLHMPgzgL6g/M
ss9z4I+MyHVI7jg1pnVtZJ+391uwiq1BQAItJBWnwO4MF1qTsdBLnXDh7gZQ9KMvxT/2YazGp7jc
rwl/5LF+WSP+4VALKf6fU5FnrBwGOC+CR89Lsg9OJdpZDCvgc7t0zd5WfErlKzgw68dFbVP7ADQj
KVOiEG3MP//fjXq3lwCPl//QPX1J9tDJO0Nf2Fwcq/M2viSa+UdFBsN66LyKWawefOrg9AepbDYc
WshEmnLchqTCJTc0xic0KLteAdFL30PEEBO0LhwZRs6Jcf5auQeYxrtKj5134rJbhaK2woMtFjix
C/w3RZ+wvKc4VIuf2vTMdS4IoZjCz2KL93LHGX4nL+b20f4nX45V1au0Ym4sYWXwPr8u0fty9snF
iayjlHzQ0bCgCMfMIPAgUKtLG1ZX5vOzo3kYsUolcUZS+Wjmm03+ZckcrevYoVwnpx6jn8pkNLoI
rrJoKfr2KTZwlRR7Spp2sZB+dyIid6CcTJm6lvtQvDOt5dZUEXFHfi/r5HJ4O6TZo5+qgvUkD+/l
+KoWXeA9Th4vAPeRRibbQFXcW+bf0WFVSFie1TXYF4wO5xS3JQDnxjX7LWw9iLs30Yg/pa4m7iSM
EDBgFGJRdcXpryorvJzopcgbxepr4lAzBK5owncL9zGPunmtXSpUD/ncHs7dIeXhvX9cDBI+ldRy
cFT124pkGo01sorOqWRQyu0kAAvq6ppLXKJRW1xS9fY3Xzlysbbbat9ToCmeXT3L47vvE/sGA46u
XnjTo0FFaewR6LxULFO/76/ZTOC96fEQl0kmdnJMMocfCBAYjarqL3q+wfPPwoo0FZQnQAh4WoV5
lETbC069NArmOv9Er20OR35b/G4TCeJipTqaZBTawWHkF6dkXGslWx0TlvokLxh/jr9M9RxU6+Bi
MwlKZiBG0BsotMelYXiBCY9fMvrcnzhI5Y9Yp5D2+Rlp34CKAn0Qlibq+HXeqOKJrr29Nj7vJPm2
4R3AWuf1s16sW4BdFo+awJQRpmk0XZ1HDR1wQqtmQSH1aFC+fHcm0wH90X508UU8wkDLqbZ2wrzv
uruN1EF707zYHagsh1482ojLvmPdTxLfXz+1yEn0RUczUbj5xwgC8t4v8ckMul+upjabjI6VIGdD
74Hc4KN/IiDaYgsf9w34qrOnFnDRLcRyA0SujpB6FMNUpREDIUYODGLzYQlN/ulFkBGQzueo6CRv
Zm+72g43XhHJyLoMCQ0Ig5GpzKeG8/AJl0+9oYLNcrI1VFS4z+8CDgzysoTmc+kwIz9iIhCmb91R
O8lPbBVXkHhv/P9WFj4jafGLjwZocigvIV8WKVjENlEHr+k28iy4M0n8hFqnJI4mztLMUD+4Qve3
KddN7asYfn8tRDUJpwXAYNgkWObWQZlkCcFBaaA6iHJUD4UmMj40D8FQwJgRu1Keo7v2vZpTBMFH
m+jhc9XT/r88/z6PoCTjnEzW7copmXu/fIUh9ghpDw88ZzI30IPxX/GJDriXFNn49x+3vBJDrDCX
c1VehseV/JArpwCMqe8SDg+oJyEKrDXwC7E6nCDTP+qRwGNQf/6CycLZPoYlkWflDlmxVvVyED1L
eRxNl8Cz5T6QjkiQ2JcVjdg9IMFXnJBWEN9HU4fVWAKKcHrujh5ouM1dZKHsYyaXCmwNPV+uhzxh
v4r9l9HfxmC2hY+H5wCitrEf8bnlBoWiu/MHNgMmS1q38L3zRdRgIG5ESrAMikW5TwngrjpB0dDW
DxZQALOu91W3PHxZ7+83TFVwL8i6HLOjpPwauYG4emIgefJHHzRb7XbkDtSt4s2EjZn/q/Wokq8S
9VVGjHbGXDYpMg5B7ZZYpfg/PDL+aVQ2gheqS6+7rxtS9yMAQK/SjLwgli8pFDhApDdFWlJdR4k6
jBYMjRPVlYSAnhMlNUVV6N8cWnXi28QKVfcwtpHqs5kMR3IPzrEDSqXuMB9+SKSZmMRCZch+9OdR
lTn8wLCQZHVR25+Ho/yE0+bAJW2ZsYllsuWypW3cW3VdlxhhkP2vyOq2KcNqUn9KRHRFMPOtOm1l
dPQEQc+s2831qTDRQaPW4Wq7xTQDm92gP+ciQSkGFvj49HnI4Xr2rba+bzxXGOEFtvYir/XyIwuo
qULjQ15o5ngD2qa0IYIZaCbpx8Bff8yjNismjej2HpT7DP1mq/FyB/7hEevS8WaWcCJQLyGw9jzt
rS0SKs9rrOakHs+iR8GErM8uTWPOeSSLQ1oPBb9t34ZosL/erPqsYF4KCCR5VTRVBTj8EL41d51K
85S24R3XHX3LejwTX9auxwdAMtE6wctNYIZfy3ZyxTsrHTFEgZx/1PkbrniE7Szn9Um3YV7bZZCB
qeik5MmZO103P9HmgnUPH9Rg+yX+zOWrWQRVPuypfY/7FoUb3vv5Qt0jn3GPGvmu4q8sBDRNtimZ
DRD8ASn3SUSuwxIsK9gnP9rmlAuVRU+Xz8lgwsq0X7hoMy4pRFVMSJ4d+m9xvWdY8q6DuB1KXMEH
aCL1mcN1rrLjAugziwqPmkq6eWhCrzxcTXZL0MJJUktM0L8LWBuJ+B6vMm51sXoMndHvw/3hY40n
t6TXl8NYL5MIa9j+SPE2UpnGcCfbCLYrIGbv1TOdjvz+Dr9g+rFaTQNBuzt8bT5G76N0lrT6Ek8T
AXM2FRjSuCzoTbwpuaVZ15UAEMjlbGEXee1EsbNLs8Ur3Veq2pGkpT8EDyGWCLxk725F8Imtv1OS
W84e9dLMZulUZNzNoLJkfvXWt4aTjnqRDHm6oWWvuAQrYwh9Jry52MwMrOBVraVhyEJpUu/qW5tk
8H9ev3H5doq9E4IMu9SPrRA5sQMnJPlyp7WTI15eH9340pE3OoIPL2kVnCAKeDa8RTEltpwJQzEr
mPT/oSgq766VZIkEl+jdZhnQ5SgXBXeQ7z36BuHttFEKV+xd7zU2x0zrj734P9vZsLMwXX2ppJM0
noMkHruegFiW8jl+3z4ogGD/rqYVjLhDb7uI6Wkv4wWWiXOpm+cCrg0ZoM28sRP6pifCxLy+B4Fe
Wdm+vuUlkYbTNdO0incnCvgDQBfCHG/BhwtvllnsBstnXCOrLPjNpzghavKb+HYDSGldIBO3JKvP
zn+IYlUSdyHEIDNU5DO6y/4cFM+ee4CyAkvki3R7Z6MbAoxyAYinAAnnQuCLR4oFSpTVZhLtUpFm
GoBiE8aNXlx9TMyC2WBAFJ3ZyD5r2V1cWJfPyW8Qpwt2nWAzZw2vmRJxx4L1FaGB/7SXw6o4tvFQ
QWgFxrK4rC9cVBUSZD23ZiEagvnXp2vCKuOX1Sn9bJnLduwpxTpOLtO8ICHUdWYuYWKjkbAsGrH/
5WyUusDWcO3lsv0Of/cDyn7NTYQqY09ldmWNaoErp5V99HdUzicONi129aFQDCzeBeRsAzLn6XK6
AYQ2malwrHFENjKPjOySVbqVP3zuniZ0kTITljCdMOQoKQb88avIRJA9RN2qT/GtTJLwyRzqZaQD
moc0bMfIGU0b5GfmaVNuyQrnrwZjINRYvLx0uTHNFfAyEZscN9hB2jQP1wThxaKswneYA5xJgwXk
4HO16FPTEMWBPPH2lXLLKPlYkSt7j8ID2+XoWAFK9MzxvH6itaqEd7cjrwBP8T3bZD1AAxHhJ2bQ
iW8ILmjh+9dHPH9kd44mDK5uHNRGICMj4DzfGIZwv5BjczRyogjBHGkiKtadF6jikM8cuaq6T+Tc
wWXQdS3y/PxWXurIgwMmpKSGkMKiYASD5D4RSlo+zmZKbKAMjzK4zadtrPYDD68NqNW9hTNLUI4r
lObph3imZsFWaKrLH+Y+ybnJ8O8EbAgtgDesvdfdPLmgkqozG8xGDhdlzO39tD5qp4APKoWiNcRE
EGBJPwZgqJjCGYOuk2kA0Nygai9/Lj7lBvI7be/RuhY/EZD4R8xBcX9q7mLOFLRl8NoTlRGjJWTZ
Bi1ru6SJglKKojOp/YBliGALAvjsPoNgNO9M2jjaZ6IOCwAOdg2ZefS+UUki1ZtEw9jD4UXJEqJd
/A7CPyg7zO43I7M0rp8UeQx4pkCV2uOpaPUalaR683pWjidwg6Sm3q9skQDWU9rEsk7AIvZlK+Mo
p1Hip/qdAYEAkPUBY+tEgVGy1sEgQfYSnuCMNM1XoKF1x0v1kGikc0XYW12OlBhU9phDzhp7HI+k
kMwdzwy+lWvt1Wlp4OCLzlO90Hkyt3KwttsHXI03+SaGaVJURB/NZboJ8f1+biCGSvBabVxHKDF4
EqQr7vNxafuM37o64lsQOyQwkpVFyh+iH3cParppZMk3orRKztuQtzfA6WNNs71NAHXUJ8LjZXv9
34szGRpQpztUy7DiXHkYgsKIAhd51PlmnkFLm+rK+sy6TKuvJjfwqUXFXMzrPNo4if2B7KphssPF
iIJeSomrtqQ9TDuPmeO+rEpmMAnUSkDtW20NBFIfifIigzYuFJP7ISEZAS7E+lXeI4XkfAi0pVaS
0lapnpEABe4kyKO+FEBaZUybi+BMPXroFZuhIllFoMIa+9JF0y2hz+9RKfVXAH6T3kV+t1ByE4Xl
XR7wbh96DerwFbJPt8rq2BoRpS+OJrdqarolABwhSkqZ42ZUu6+l7e/Mh8OJ0sMDm4v7tsu6NnGm
vQFSo5b5mjLOu5f2QCKSoGDt4JuDk3tEhgK0yqKK0zNap/OIwf1NuKoFBVE2Xsx4VhNVvm/WL+pN
eeiDJwm43NARGv65gQq/NVJIpeqzYkqMwzTvZKyJy8yvp9NEJGVn4vlzMDKPDDq8Yk1zncZkvBtV
yH0DsNpC6J8C2Fz3eNrvsmEq/xYIcyKwz9Sb3pFF0lvRVGTd7xCvX+NJy5yDCuHwViRhyJt+nPE2
ESOmd+X2pMYdMzEIgDwUlfKgYOR0uJtNQI4grZ9n6yEnyMPllLV9yuZ1+Qp7GHx/8VWjuNzjPt8c
3aktSiCb29XQECw+UDaJ0H5EhjDBKwRfCiOQr3jJmVl5t5a/y0IhcMcrfWl9xP6Yldytl3MRdQgN
jXxJBPgHRPizVEmLZJz5ZCGoWhdlFrlXlZNfKcGGmDGksxKP4C+NMEG/YqrSwfkG/DXvlranNWsB
lzbN7P32WxV41edrxwH6apX4KWbP9KVTD0+7a3Epnv55rfbkzxfLpEqEaoYMX7X1jDbS8sruEPG9
lu7EUi5kyXQ3L0zUwqrUU/ATE352x1u+7t7WVzJLrYthQbwBKGUXpmrf9ovrjNvqTVhiZKrhR5yq
wD+Gf/2ttuk4z3hqg+38iYsvSFJUG8wCHrlK4D+WohJ0RTLowesTiPxCatr290qEmE1WL9e7mXfh
Wsqx+p3Gu544leZ8ZVba4HmitQw8O43RMMIIdEIBfNGffPdZD2DXbNK+M2t8auI8tmuOqLkqzFpb
uA1D72GeIfrl0g0bJKfqK4y6PbHYyiUj9wdMMIepvba5C4cYAng6ScYHe7s0lFC1iDvpFpNifop5
nuWsbDxCTOvJG0ZCMEZCDDj8eeRDmwbNmJylu2VM6xJ2RlwTgXtHwE9aK5afrqUIHjBWcSNYDw0S
Qck5Cz1Pi5jK3Y9+asvChFLooMZUSfkjF6ZZPXRd9heomLllLRhMT7fse3z6+bHaJOIBLzaD1+m9
X7Fmm2hcrnhquvGyUSn1zMZQfnKy+aF8GvzjF72IfEf549WQRkopNq96hWjVKMjYDlpinSdQW4Jz
ggdEc/BxFN7gaZ8lT56IQV4ZaLJcrGcj3I3veX+KUxPQBPoZT8whcqgurzXqBsC5l04upTusCTdj
brYwoyNpRE/jgf/sxT0fVC/SnsY1Av5SaDYOuoxvLYTJnuGFGxoX1aYQI9nbDYuRJYKZD9D9IVUC
MYcx+e4eLH5bmexNEJy/k3qBNnqOamXo1tN9w34lOKSvQ6eCjmuflHV3/gxRQIYXx7HJtMMrOtYH
8W6sUCm6QIyCD8gtXwzX1zNvg+/Iz5Y+zx6A+ZQshnsSm9dqZxlVP0gtfbiG2Ls5HgELr9kcY6Co
5mPlEwUAra7udHJ6ZJDN52KOC8Y1pDF8+Fr21wKu4y1KFOhqIhM3A/AzOC4rewtigCpYLnZF0AGV
TshU9dEmKgkOzheEOBBXFRi52D26VeG5zH8VqVSJ5OLFVK1DLzTovhQ4Xb3tjtVgaNCmchS10AUs
KezHY8s1pDYtmO/P1ACdx+kq/+oNdAmSf/HxWZV+oXWrSo8XRoSYdnB0gpRNSUKcaWr4ycq470PV
GgphmfkKnp2p70WyF8wShUxac+/p4hUb5CQBXV1vqXJuHIjqjAIXibOM9CHv++VHAq3lSeOlO1Hu
wIpnkOWDtPlXzePuqqbkXcnkGf+WA4izTMUuRMJojyXZ7ebsI2IkxRA7NXcw45pOgbdkPPFCtGI1
kmPkFynUXGa0CwbHeyQctyrSNEyGhTP7/U16OvRLs5BMqAy72iJ6i2qtfHwwuhqEjhKxk8XDQcP1
DCV9P68bOKnv4Jlu8gRsPSaonvvoMUTpUN30rj3iOiPynFfT0p9t3QyF/GaQ2F8JnDAKM90I1pN1
wOt8eF9wJhpM99ARbHJSW/z2pSiRZWI3n3wShwHbExpMO2imhr1qb90fizP3S1dCgnW9IE1xXQl+
FEhHN5mufGiJYAuab4mZ/jTZmlCB75OSROnZSJ2rIg54fAceN8nOGO5uffBaHfKd6uVZRkQ0G9kf
DZ6MipniE8UonthG+OCPawcdPAqAwZ9fZiZXy4/OfJW/AYEcUfICuO29wa3sGcI3OisqJ4PJqcdQ
2YRzyD/2pcVETTi0ZzANStJnTUByVTpPM3QsvUxr3q3N02NSGVur74jFqqB8wYIWtLQRLE8bFrSg
mPsJ5Bc4x0ubciXuiLWbzdJ/12QUY37H5d/1U+g3U76HsQfNBsUoDfYcmqPXLoPLcfFgk50xdtbd
sBwKXt1JX7JN0CxOi2263InIn9okykR+6L3ZE1O8rWzGOMkHEogiMh64Sh/ROtAFB7IXcebXaukz
NEIztyRyTpH8gxDvfYb7LXETNFX+HA+OwFTWkdzLmqCdPXvVu/8IKK+DHLUmwiqT0gOmn0tP3Ym0
ZpN8GTW9I0c7j7sAIL429sFVeS9PvA2zCQ8BxNa3l6A1RoIKoN+k8rXC3YebxtiGDiDJc/eBC5X1
dFLiP4/1++5ml6ZeF7DjiyEPunIoO1raGaP4u0ZN+CSnomjkbuG8QxQfQzixFpN8HRv+BROQ1bwW
fUZtg+uBTEJEOZ8zw7ufcH8PugXL1/vSibSvScpnY1YS6it5UHv0+K9NWbzIkFauaGYZTpZYHg4e
XF6sWZyTfQc/9yAx8eIlvh7GWF6UXljBCgn424tscVC1KgdgDQ/BJ39p3H7RhZqMgsslXxFYX3Jw
/O/9l2qQ9jHTqpvQdsEPQJwsFq6P7LxbEEJ7pdzOsWaItW3LCd9UUdqcdJIpBKkfYdZZn7iCBFm6
4NHjvsZp8JHiEuT5nODG1HLUpGryjjT1VB/P1vQyL0nR/W4xNihuiuW+ZuvR9lMAO/BIwDdAsNaQ
+ql5vOV9rUNLTLUiabbCKucImiN7Xv0Wd1rcVAKCd4wrt34F/aXopr85hCjRJ+Xo5PXd8vmyhoPm
klCMAYB8/mKxXIpgKebm+Nlpc3JkFzDkNKxrKFwU2nYDByBJBd7t0+0YDWaOBaQ+ZYRSRjLnT1r+
KdtiG1H0SNJnv1+urEyP2CANfPyxvK5oOLFtSFr2mnH76meYLf+X7fSplxSS62yKTy4epR3QIzOm
HgIXPGkVo/z8FCsTpI8FAk78QsrTFVL87B2GLNOp+jxF1zaZM62UnC9ydLLDVsq/QR2xC46r1Fn/
ARSJPij908VIgGN/BPDmI/o47meaAa48RAVD50S9fjhNIRLe1jGZoaR0Foi1ltyd7HaQHlZ/MW4G
0YCp81Xac67CYZ4+uScu9jncaEwQYvn3Ak28zTG4njzLvJdbq0QMUdVPlzfSJ+IU7n2UchUZS9U+
j7Pz520wN0f4WDuq1xNl+ft7vCryatNS+Hd3j1I+Fb2LrbXYpAj0u6HctxaMdGVwr7rrZP55SKSX
dSr7OkU4T4LjZcGEHO/i4mI0QgOd9efFliJMZxM52Tnc7duTYDZXVj3JaLDjZFnVusCTCgr+faJe
U4AOU3lRdREcahG7DOqp18hpyuvigaHO/tX+EEMs8F6KDSqcBBSlGJZUMtS5LaECSooRUclZiSnR
YAf8p3HaEW1XM7wEQhcbWhRrNpLZ7KpuMarzg5kxY7icikPZmlBQMIinbzPcDHzxrpn/kGJr1D+u
cdC7J2vzGMO07HdciodSVKaXqIQBUQJCHgU5Mkn78ticGGr0wTe3/lRrY+948vt2l/BZo4z1TM6s
Ea/vP++B5SbMyM0dKZDch62Gk4ILrsDNWUYdUuuKt1hqZQZ/lVfS59GF+xnWqY/d5MfBcptqrD6W
vJxor5nVHBtCD9wwyqPL5tJVFAkiiZmTrXdemialT9Inqq5UgkbbyVw0l3Bdp7LjiRwHOGtqex1n
hNO2w26czIAbMB1FbRIer4rjp9B3M2/5aYiqXUXoWQ7Rb/Qycfdl/Ur4RALxiHiXa8kYpfCxCyer
C1suQeaFYQBuumwM5+F0LTBB4c6Q/jnCVSzVFm1rMx/wLDYdEclHL6ndZhAbBO4D0Jp/yVaCRdz7
tVK1mnRjeN2ksroZQ4yg1nc90BRdgEMpkig5w0S1mQo47jc52D7gmhj08M1YS+ISQPUZz8sWUr1v
w5aQKxVZpWor+aX522GH8U1+2OdlAI9mowcl1gcVnjspcPfCM5Wr/18TSZxnB+1KRS3UzTV+zS8/
iO3HH2ieYh4JEqJN5IS7H/+2SnQn6C58jTWMzxCmoFAjcHJ/P93AyP0btpNgtSxb24dW4pnem4us
nSRAItp5Yvzzi6aTifU3vFlRzJaOVr+f7Bnmp6VKNMVxh3MLx8oHCFpNmrstDWyDsL37e8SvWohG
z0Qrh8fVEX8tdPuGOhx861Ytw6eonHwk5NV1nSMW3EgEe06SXA7CU+b8TzNAH/kFKNBwwCRCpYOP
lsQHuCMdkf2IFxwM/WBkBBNvr1tiLRR8vYIap7llGjzlFRwpubKQ9Jw2IRcXRoHKjB4ULvcyCEQQ
A85HJ0YY62ZpdkCnLnaqC0Jih30oA180Umbb0mzv9mBr1uzVm8ljGGZC7h0WyHgXeaFxFsvOcuan
8IUkFKQJO/ZRRdNTJNmA6QX0dZDMmoQbg49CiAuY73gNSGmI3GbY+xV63JinR3FRoeivZYIRFEJC
OSxUu59VMIvxWEZ16+jWEdA+h4o7yET9Drlf5agA4EoIA5KpC1HOSrT8ZQynkax2ww5h+lzBcm0X
orGN6GHjZ8WNEKEMZzZ2pM8Br5a6z9TLz36ZIbKJYPd0H4j7ae6+d4yvRx/1N0rMObOxN/c94+g3
4Z5Rk4dhESdzryfbftU8LZNPmn15WwXnmlvysZx8jNa3hRaJvN07tiJ4Vnr3Pj2Q/g1gx8Fj46sI
3cxgNGp/ME9JeuXklHX/lzSRw+IOhlt2jqRMWAXlqbBaB3bY1Oh8npJX8OlF4hNxfhxXP99ZTTMF
Zm+iRcpHSRkJYRs1fNulV2lRnasBkuhaAwMZYBAVSw3TtHGrcXjmlBUHLzln98jTnnEmW9cuKQIr
GxuOWeQtL8UNZ4Q6F9tRU5EVsiIv6kqzLpxIU9lrjIq/DUzKmIXuRNMWKXlqsZmXhg45ftY6I45o
yL1EMHakY0UioF7CEe1TZIlHoeU+wiGFTx7cQYRxrWRCLQbBgIpe1thetucYkUTORR6oQ8oeWP06
QUa7O2BVrnmUgxV2InZ5qQLHGqndr/fsDW2rtcxBkzaAXxbVoBC1Wg3RF/UcGl+sKiZKMSFaHFWO
RR+FEYxi0cESHz+ok2nZeM8ly+d6d7Qt3XJMalbUeWe1MA3FReH+618a+RpPNBynhU4g2YjhEj1D
1CrcaFLZ5zO7NwYdGQk0AQslK34+mdPyxfGbD6dzmtak9LFGgCq+fJf/XIMYBxDXMrCQsV/L8Gli
n6ar7YoUrIGYPlLQxqRqAEjpXLscCN/AllzlfcNqigBfqjmPs2tPNdEenhpmHgmC4jwJC49GvHbz
+N1i2aNIP0yfqJ88zR3avziDb8smRYxEs2FbDgW2AH2e/cdDBLAaBTo14B/4nU9a4jvPNAdUuv37
xOfl2kEfrWHq3ttCa3kjtfUX09Dv4mAquUnkH5DqJf0/srgm7d+3IGV6XpC3mN6Mb5ipdCD0Fpfv
Ge1gvYQm/XeKca5f0Pl6RCUG+Rh1u4Lz1nKkhsyrHvv1b5QZq5AcV4MfhO6tdiKLqo2XGp7oN1Nn
OWs2MwU0sUpDGEuKVOHABeJ6lH/fcqN4gxKuouEXbHzaSb+wltJMiNVRd5lEZU4hlYxKihkTRxgb
Q1gfKpvGUKMFkXFWO09g+6WwSIXIHp1jaP+4AZax44nSmKN9gGnpcJ+M0TXicZ6FLFgjSo/dTriR
LiFna/ou3xGRc9n37j0hfNAEYM4kesf48JGt4/Skm1n4roE++GZUMjbq66XnuWXF71WrK/sKb1d7
HeE/EeUsM4plPMa3XGHHi/ei8cYyfdjVOpUG992lZjampwNIVghYDz0lL4xGnYku5R8xZatz0EVC
s3osK9atha1t2TQbZOu9mY9bojsSoO1fFd0O7f8rjNM7ooWgAuYR1LXwukHHXQTZ7Txw/FmH7IeJ
y6A7bCVdtDkNpNb77/Q8ENxLuAMVbXwVNXQdHoac5L5iCrGnWHcEQAEu1DWg1vEjzuW5lH+dFCFS
szw0yodiMWgNFqgczrcTGGSMWPRJkq9ZUGdo4VUIcllmsByNCeRBaRMRjV2fLzXVR6ZQGWdkboPA
nXrwLuQFsnG/A85yrhs+3iYfDAf+zuq0ZEXReFX32wQbMuB7ZlVUshoXwZiCO+/ur3hjvQa4Ec7k
V4FD45vKRzxXwAm8M/XLyF03lZq0ZXQWydWdwg1bv5n4tAN7yetjPjffZjSKHFs2vr7pSKVB5iR4
gE/ZMxTnSvWF6i/r/AIHVeQAnq6E6SU9VsmKmVOQ7805Mz/cm3s8u4Tud2rBfj4Uvj9XtVFNs6/g
30lg9tmi+nojVDqX/1D+yTEoZBuSo0gUpkEBUJ08oU9EvWWNJW1RKO4QVjxS+XOuNO7Ace1VkXKz
1fYlafmMrJ8HoA71nAvKIo5U224sSbow0aBcp9i8l9r2E0C3y0roe/VpXgbnvRPt3j/tOQE3wdqM
7FNPu/9EH9736v0zQAbdm6rNGB419e+a2+5Yl/5KWDeJtlOeRvy0NcV9Wr/qro4TMOHLvtjMh4pW
vzyZ4p5kbbqyaWr01+mKMYY1kDrZ+oC3xLdAAzmbXMaXrXUP4tx5i6AMF0/S421qdVe3BqnGc7jt
uQVWjjMWTPKxckXTOEI/x90AFBbeyA6z6zzXSQT1phRd8CXgTiOZctZgFm5fqDX26iMtnnKLar60
uvpd22CSmlmtUK+7i2MlzGJV7dvJ11N59Mc4l6W+YMmTEB+ZW8VbBtwcIfQqdUqbCoYmaBw1FfnH
v/OWZYQ289GzXSmwhZCBBAMIE2Uoyw1NOEiWCp/7/mRm1ljubhj/syu2wnnxsk83ObKuJoYTNRag
95XLnAN6MsnJ3Xg83Ir6qAlS2uugeJwT5CpNPUE3HmoU52LRnC2AsGVjacxiFdCrrtOOucmhhogN
1FuYC0/NDMHEtudeohkcc35d9edn9CNdblOsKsMWR1ET9cB1nueI9l3eSUBHQGFty7O671M8S3D6
u6Je08KQ56rh/Be1TS9VG134R2i/qShx3X6SoxfW6a58v0wQDe3wetd3dTsapCj2CKzPjMJTfPAs
stIHvNK9EYdKZZSjXpJPShQI4+qN6WM2TUk2nUpfmNf009E1j+4BJwXP8gX/lcuRT6T2SFaWWDdv
hPyIHpCvhcQHnJJ7K0ENhv2hJfApxoSmMgBkxi+9BusL1Q5YUwT7kGjWHUK31ljm41Sbk+jVkMCJ
b3yWJclfelt6e7HaCQf798QuOeOVKBleYqDrkqrgKw24Jiy3KD5NtymkfmoQqOlVfIHKM3tyzYKM
OU+SX3r9tRKNP77wtS0ri8N/VcwW/dQ3VmrNpjppbMKT501/O9tv8cpLfit30K23cJ2p42ZWC/sy
ByslwaJIzDxeLMpNa3UQCyRyXEkU798isCR7WToh6be8ht6/EfbQemuxs3ynlYvazB+89wlv9a0m
Jxsi4JiIdpmpeOR7Kk7EW1aeZh3ndqldSPFNmShgbRPU+Dly84ySY9eS7bB+2rIXzTy3si2RCzqQ
sP44xminf25izArkM/0Wc+1pIgZe5Gf3nbj6SgIzjE3ZK0ApZWtypoddDD+1MOabR7duS5ctmh68
PVaq0PaRb44KHS7bzrtkqCkY/zKc/8xEHEvsL7CS+kgiPDYOA/0LXxx0UY9LR58mJNX74K5YL+o7
Yrqu3eNDWmrqpxC424vd63RXVab/M6prBnZsfC/UEJkJeyDaH7Nt26B2wlNDo/H/oXq2K0L82pUW
V47+99g3+dYgQYkGcHGymXxuk2sk6TI01eK8HO9CjxJwD5jqjypCTSbNyCuMFLdvc4ou28FCFlvh
QdvvzsujD6me9yby+NXxvvAO9zK+2PZ0q9nC/2p5fMxAaQGyNalg9Z9BbvaFEGq1IsLHQAswicP6
c0sJBzSJxQ37izgcmcJmFqh5igxZpwOgxC4TPaOvsrofb0Zhclga58Jz9jKSC+dnINnpYVSsy9R/
zJIxJrYp+y/SxyBPsY3cwQu5WsGvxSsrQ1HyeAC1Dshy+V8ucGELYJ8LmXm0SQn4ziIZAQfO5cQ5
+LKWvqQUQkQ+QZl1zYyUWtoVGLNvs57NqIr9q5QdAc3rjB8bX+MJZEwNM2R4IDcnL3Z3tjOpKeU8
onJFrgsxwkImTFE67WuFJXsucMfYXvZF3/CoPaMW9tS/Kdf44RFYse8CZNIXtoYGr+ASnVLLhEtV
kOsR//PuiiH7PX8CAFrSYpY6altLkwDpIss3ep1zk1/YPUMtNIiM4CpqWqdOGsX8Z7ZW52HmUVA0
giHwhqONZpqsiyE/MTynKA2NyxgADWw/doMGYOPsiZHvCcTRkpx5gHapTmbr3zmW3DZbjr1zQeeA
CpwagLuNunyCD3R5P2ukO5tGoHphto5p46839QawWBl9BMfFToxd4tSag5FBeHrHru8zqHhQ21xn
VbvTp+kzPDghItIehwdRkElUWZSePkO/4Eir0DQrz2jkjIf2Lz90SM4MQSyMma6kfDTweHc/35P8
CkCyF80EC/fowhW7GSDlMmrUDrJTw7zInDQARkcKO4tCI6txOSCBTbJbPK5aXnjCjIlwaZgAoUZZ
GDqnYabp6hPdTxjF7Tdb5F+Bg9VBhap0lKFlnA7+9l8gRpjwfZx528QssCoRRX6xzmZddiiv6cWF
H6Av60LrVJcosu/qHOWJXsOXcsL9AFv4756r/tEWCu0dCHzLW1kXt3nw5ppXiKFUQZBpOo3JQn9f
AW/mW4Cpz76L1ORZo3QPG7bwtThdhj0kix9eb4Oa0zcFNQgHb+W8LiFZNtvvFNt0mMIVwxmtTagJ
9BoAsT8RoUewc/25up6oI1DUUgrrXe1Kj20nF2hqM/4bP1jN7bZWyl0r1vm/lZAvD6cf/6uXJ38y
7KguvYDBPWaCRwnoh4zT6i273at0vix3K0lr3qJfklDEA3b9tyS6CVDsFPcKwtQ463kcFbS7S0CS
MBIJ0KbdaG5GfyU4zfeMxyagaCOMW9kw21R9xNCEqH5bs+LMMWRSkpjZ5dSeYAcoZZmNcgwoyzSi
HP3g+LLoTfTmqbdhMRlabfi68tIF7uBmQiASLh7vcpUTUajk/RMp9V5ltZIgNHEwsu2D0Q46r7n3
6+KBLZkFzHyKZ8sZSH5BMgEbmp4fWVPEXMedwGl3PILnONNd46ZSO8BPA0Ah2180wfJRFx3J7Xof
Mc4cm1l+JiSa5fR0MqBvOhT7G2sTlnNUurXO1YQQsaYtLSHQ+DjinV5/JUSEyYZKPa9OHO4pkKHi
8yg8uC02CuQnxOwyowSwygVzrCleFsZk2ZfStDBEv5ysuFTvIebKVKZTir8yL1mZ/4gSaM73XYAg
99IIq8uYxp7/r9puKSvndgdo5R0UJB5kYbTvuXkLrRjxeftQlYtEk47HeqOCTmlx1StfH0Ppdwm4
WYTQrCam7L/Y8cBH+OIMKLmk2SczgdNOfAeC+t7TOOSX4l7393YLTry33iiYoNUg7FcbInaSJJBz
POqpHiPT/484M9BnPJDOEPR1RgMACk2qrbLQkrs2cdJePT3o02vjYhJo4RLgAlqNjIrzXAhcFMby
+RHcnB83/gyUSDsj8eRVEOTNcvS4IP5XgdwZ/Tltoyq52a6ggw7x+0pzgkPo0CVgYYXyPDwsVENF
tfinSDaC5N3u5AgxGOgAtJo+ZwCGXQT0Kc6uAaSZSGynuZoSn0WQCriiCFqTzxj2wEpGq0d0f58b
ythXM7fTe/BtuMnvPIhDk8RyIpvHIH0e4mkHdvuljZH8Z6Pc7HR2gMzUYQxjNcY63T2rObJ9uc96
FeEVeJ5FvauXEPyw9TJMXspGY6MLADbzZLuZZt5iy7pEjKdyAK/+PGGRkByDskUrOz05502kT0Wg
Aio0oEqj4e3dDCRMlyaz0SuXKl/XPEvl7VB+aOfaEDFtlklYmqt9RAvd2WnRtkaAT4WwFGAYqc75
OR/4TkuRYB6wXs5mWS0UOsgkakPw2GUEUfZwtm2M6Gx5s55cskKAnrozjAupgiKeGqJevuvBIMJI
AQlnJ3DQ08Dh4sg8xU06Ku1rPxdpU5bak/s1e/gAjOiBd7kJsRydvpGaaRpdZvSE7WL4uWnbQlP4
HHcGedDX246rFmPNfeqyfFtAkQFh1zLVzqPk+5f7BbXXrxITeWrF/F18p0O4mubz+F+2Ir1dDhsc
QLPKE9JZscZhqzdOtgC2DIQru98OKdwAv9OjM+FSU2K+9cR2+hPWVYTUXawyIFFyueUKf894JA0c
KcRxIpOkEOPJhMAtDAzM+qEuB5V2vQ6CroTdlIZrsseqog/p2YU8DDL4jgcv5d/QPeBXOkPStnEg
Yrh339xC5E7vAmLNUpHKTTS1yj/CHw6glVHIhFTN30tIedwNMjuQjnsBwDKBfZR7NW5b0ganPUrw
vj5dNqy7Wbi4TNHUNuyvJK5SVQS15CuqkNvsVAJ89VyXtWGDzR+SC3DfLhWCS2dcUf5KZh7vh88t
YyJtCf35BFIGlNCChKHgS6Hex80u+Ief3ql6w0JyQtOcr8oz9mKgzhRZrALnBw0sgtaShR+da2lb
riGPQiQN84vnDQQ19AEUtnG2nuXyrEwriYEJbhsEoCRKr6zIsffJ+EOhU7KnHE6If0vjBBv+NEEM
t8yzoxA0/O3wqO4yI3uWT11ZXvaCKve8ecM/WlgEK2hWqQohoYw0dsYl/2rfKg7tA6ngmRqEi5xm
rDngIxaHLVS8q7VDuRKGam8pvKCrDK1WCHUgxr/8VhF5UMl6Bw++ijJozBOOYfit0aMyCWpfurJC
4y1iHonX2FljI2aEK47aDD1sSNMJXR5F9Czz3TYZqhKyHmtDRpEE8ckAfRiZzEdkH8oDrAcgFiIu
yydAo48omsDE9vX/JuxwdpD/ivZ82avGw4aY74FPLOecFTO/fvumuxrtDG55tYpCkM40c811LJcn
e5YKwQfotZIc6pP+oFBIkR2do5xqsJIcafpfJfzv0qi+I/rmI9fZtJJ6FTUsvOJTio9ab+jEwqbu
cSBL/xA6JHhj8sSG8FSnnUptBvX6tsLijEJORConieyXjyVYEvjyLp9vRimpQzbKEc57q7kj4U2k
anY8S40WvgiTYf51Mk0cAeZ86lswlf4zHLsyAxs6WT/927gtENi/5wGt29Ir3r67OVsDFD6vaofQ
LTpbc+UTGAe/u46Xjx7608K/tS8fSlFXvwBE1PTq1QY5rF9DCfhSbRYuG/AHw5LgIgXW+p7Izcki
qtJDqpB1xxFkCjHjNh7SL3iOxWD/0DKv2AhE0kRxn5GK+2JQu8OsLCf+rOaFW2HeCk9HBc1/iVqh
xHNz4ajHfKPvJeu8Js5Y1aUKFrXHpFL6hAOjSLZU6dFxTKXjfSAh2AZ8x9w5hBU5WYMfrBqp/Zmb
A4HriuJogTGHKXP6eOZVVGtCbZhPMwNBDQ0HWCT1Lifz2LI3MhafIs27vRSgJFp9vya1JR4GLVOA
TlR3U5fSnCoRKSF73n6rm0EreuSO+/PFhpv5omUtskAk2vSFZOM7yNWlfcIisEtjlC+8J8zuCWqy
TyV0ePXHp5kdywNp09uRIXTnN/fj6A09kvwjBu1fdjaL/IxG0PueBoGp8avPLLK96YCCYysU1PKR
A6D5QukmxIeOK+WdhLdp9Lbhx2JZVhxGJfKmlMTDc0n76kwraZKKDT/Jy81lnpW/anpayTLT+akq
hgZcacj4V7q1G0v/w+3qB+naZVbA0VnMQLmTi2t8wZz/76hwfpQ9POBUQSArgWWkvfYOFM9hj2Nl
mZgbtLxf1pbQCMdsjIn2lOPaScg2JBRpuN2v3M8+9NqvpEiROVQYEPbIq1Wbqs3UVnHaYBDxijFX
MWeXYG11iLTqi0vGLhccA4H1m7iDh4KJxOaInI7LUXywsujSxdEc1M09BbrI9gUz6dsngSHwgiCg
sywsOf4xe8SaEW65UxkAcYJlShOsqLnG0sB51f/auGX9yUG9joWn1wIKE6FNlu+fnVm/8quQcsXJ
O/prEy41pioBXHX4zpCaizrliT6r8DcvrWh17miRmMSGTBjAae0pP0PaOOo7VWjMUCTKnE8mYC/6
66k93jRc6u790hsdXeYUYimFUj4I/idbgIks+2mJTdHZiHvHKqUTTEXXivW7NBicgztApieI8+Bi
BRC87VEaX99xndFPSuf1ENzvW1zhZEAAiVy7QycNLLrJzS4ZEdHBTZZvHj25r+Ir3j0L0S8vpxhr
WMcn/Z5XwlsCQqF/Gfn7C+YvXAfOka59dYmbuH0q+tCTDhECgSx83oVJazarooG7/FA4Xka6sqqe
WWFzVo00u3q6g+D9UtkJcSi3KrQQZNhffk+wOLVFMR2WdzAyJGaUTEBzG2zz+lYtFzKj4QUuJcaO
bZaOIJg3q6dTuaa4EL7URrnCRW/TxZtKkQxMaM+gzL7KjQvWGN7EaBKeHqPAv2NFsGKcykUE55IH
kixFoXR5qTTHIvmOsXldWzivxlIBr3JQEhurIaDiprxVSEXY/U5i/Q8w9VqXJvKkO077ZVhoCrm4
F1b4Go7fTU65/TER5wBIRog7c4rs7KqBComB07IpfCTBFTyWeEnj4fz7rdqjQIJwnSN+he7txjkt
TTLpyCGdWD+Kd8ZTj6Am3nuwcOAs1XXmvBFMgPuWdLNS/ZZwWlfMzM4luwjLEFIatiDjSEQPaQjv
t7Z64Wba2S/traFMUoTeuvY1o7H0IkwnMViv8pkIU0eOZ+J8gNvCzqOqsKBXethOjTX8PzPa0Bpt
rueufLvZTXKk4kGR4Q0ZWkySb1i60zKRHrNRwJKijI64I344Br29eOUFUnSagia6KHiz+g2R1lKz
cR9GjJD5vL8hkvMLvRnwr6SwK22y8R/xSt25HpcTD6KFZVYMOM2H8uJfSo2xH3QROyx06O673q3w
J0vyo+k7qiIo1DXNvB8iDqRJz+B2qoUOiiGcVPjeqYb6o/8MgE9bm4K62FRSHKQtN9DYvHpxo6Wh
aN9B7ZlmFSFc2vUAqnEDI0RSK2GB91Co6l4ANHA2OIkeBuPK/Rp2L3Mk0Ev/DgCzZeogVvHTshwQ
exdp60j2HYTM4Yjm8gWnruVfzlXKpvXp/A33UEJDBI3QW0ClCi0nSVunLpiW8n3TVT63Htrso+ff
vsTBJprFDclRMClw/48E2XV/qwH5GZBE0V4NocBNy2Nm67rlQLqgnwXKOUWpP03mVQcSAtq9WdQg
zYIvaQMUFmIV7tG1xFn1LpSUz5x2XJlgAXxVY/J0S5bxkr7JJ4CiTyhDRq8PY4Ppl6ptRbsRh0Ap
zR5QCl+pd9LcNICvSq4KiD65+p5CE4pWBJ+gm1EifB8ZBS9u0YgSWnMwVx/I13DDOE7EnaKd97lX
cGGL296jBZ5BNxJBePaELBuOVyyPRdqVZsW7JevqxNBX6M4YdcuA/PYziU8cfld9B5HHda16F9n8
ewLvECD9DXmFc80keRMl6r5admqMX9EPtlptoisWnf95sflQ2eAgxLhPCdTNdrqNoORetuyrDp2P
rtj9wnswFhRodBdC9zvlni7cGH2Qw9Po9vK/0tsCxWzIi5mKwGEv2wEZ1HPNh0uwyBhiZxeDPBAQ
iXCyrbHHvyeKjwtlZPhSoDIBZlcidAq+hefUvhMOUDBAG6IKu+a42alhi+akT2sjGmACtEvnOBPI
otQDDiPmSc0KkXiI05hhj3STPovMFpay0/sD47CyWev1LuBVdlBGkcdHkyKzxpa6rrFi4tMaOdOH
278Qar35uCqpxK9/CxJ6xUEbVrwbj7ahpVlwfBh3S6/SpC2I5eY1N+FGcdmpaUzliDEkV1mdUc3K
/h0PJn07+K2rZxwGie2kOzsv3DxoKPQdyNrLS9vtzfxUiO4woBGhDEsnLQEwxc2jvhtVfa7PzsKp
yurIOYS4RHEW5GP7bVzLiPkFB6VUzZzEktVZko30R3K43uFP/9sXdzRaChNyJzvr0U/acsnPQlj7
95fIq0zQ9fi+DSUoRsVWipnbMla8UGbMAmu3KZjzrkw9bL0Xx3QYXBflNwcqimqRMdDYtM/j7mCw
1trzsU2v5PuhifQHEsaHJvGaB5Hg+UoMViwqJDghXZmUWGP1KLddwEiOQB49Km2doRyuZMHECxRP
nheCpWqoR+FQAuoZldxnKqZA8Whv6GjpFAzeCiuMHxmknVQv5PeLOy9sSZFXiBMtKE6YxwvKJo4z
u8aGy6FbWSFvOoszeTOaK8f+9U/nvZaiZlRX+9hCwECx63iCg/rpV35C+u+6FWcIPfQ4wfRYziPp
gKHTpSImU79PhZqfy3cokedUQWYi+DL/bbwchW1aUK1TM6N9340oAhZv9+jKHFeMdvSstG+toXsM
s+kW3ZsRk1mKMqxGOW/EJHXUe3dN+Qwz6e8arD/NDyaWx9pFE/SFzbY4cN1JPWjyBQmwEbvVJDtn
hUSY0M9h1/cgUolYEBP02sJsAj4T5RWjJH/ltTLPbEoOojSWr/ftCAn/qqwpUw9vsKeAwfcpwUzx
1RIoUmtBtyMc89ZNlTSopzRJKcdEKlU2G+TS8dcYOJ+HaNnxiZr4hjrBh/TEUtb0s3AzKUJR+LIq
R6TbFZ8nyz32C5GLv3/jTW5nnnNLaACye5C7RT+mJo5wPN2PU33SEWD157T2OEBliMs4HWrERfJR
/LJ1wOAtW3ANUxZciomEFNPAeLr9h5vPUstpQhipdV4noCHRA7fTFPCNFWSCjYkuspMXZMlDCyMI
hRjrTvoULijqv9MJErq5NJRvd+HxvnUMWrCjc379Fx9QcHN/tQJ2+ivW6UzMYP5QeTHumnO6rgEc
89XUXkjTh16pd/nWGaOdeJOuITXvYkrSm4TOpa5XaZPS6/16ojvui0KxWlOl/FpXX9jldaktPl8H
K/lqqTWcLAgbZR1ct0sR9DKF39Yu6QXc8nMzi6hWVp1Uj0bt1SSdGEKvDy1N5UkRTzkm97EIFzNf
6lXX72QA7N6sYNvA9YO8PE6RcqrpYN68icmPk1GW9P0JEdfnv/TQYWgTuoR3Kz6keUREpQiIXfv0
cag0mmU12U+sf3etpnmhgJ3PNiTzuxfrAYL8xdj8S9qDWbbbCpvLvy6Zf8bvpUvC9f9dK+rU0tY7
eaYgqfPnK4JkFps2wuH7BJ7RCIoCDxgabF7B5LmqdikbaihK6YZGi3A0HaHjLGOD80eGSVPWcOjn
2oBHOnFfAD07TWurgYYqNJHP1FbyOfN+asCZ3ML8p3wuGD8nSt2sRsAHrzSyczYQru4U1x//jDgg
ORirGVRcF0gzriQz+H9i9xsagvf/0oVAflD/En/VbnpOm/LAGRDkyXtEOgISAFxhUk8xjT5oNIWo
rA4CRM7xELXYi8rwDTL4bUqFB4dWqtswvtd2QDUgESJXeIKAgWhu57A4BD7DHKwvinvOz696LT/2
nG3izqU0eySDxdweLBdQoruywBivk5C9868IFlqrF1rwkuloYAjpAA2DScl4WGWhchIDW/abwfQS
MmB7D+qbRT4fKwtqnRt/0abXEtC4nVKCa8cnDPpGOsBFU+E1G5w6sYiJVEO5QDr0/FfOwKPvxGNF
Y7Mj8iUXZtWekAuDXRhCNcPUcMnlclCqMk06oZXDADQK1LMdoG/3vCg9gKIDub7F27EE23GRr2Ws
6ox84m6CdB5Yz5QJcowzCHPkKmfMRB+9CtDhhq7hzQoelDPQaHQ3TQriAWV10RXDdpfsQIv8vJch
exUk1onueDBcwJPD9mQvBg7H7FJ2HxCsV7I2uOyb+kQs2irBP6D/qyQDiUEbsSoLkJ/tdVObCSoI
R1xuTgWGsMvq69D45EqV3r9MmVWge9tWM9kJi3Pprl4k3qEOuiNxUUyDnO/05YisE9To8YtyZbCz
KJWuSHcouiwzYp46KBqaZxRomTlnMTEVKU/cbxCuyRwYpVzqFshTBps6YXxlfVfH3eqQat2Qn4JG
6pF+4BBIlAh/bY9fI95YggJ/25F57u3qYK4Mt/GcvJomRTLAoyRGaESvvWK0Z4zfz97iaTlmko43
Vi46QxCJAdz+PM3RMe1okHqcYop9e7PCXtW4HzzKENKBHrD2JOvT9h77hR+7orO2hLwF9qpVcCyg
ogvNfrpH4sanumBeHrAT3z1Nt+oCLgTkzfuE4n/HUtBpeApUyPJao1erns0ZLxYuPMVNfgkjIao4
AuJ4yuAAqtMEKA07UGtwQu3cvuGLSH6Fu0eWyl0Q4gqDLyTC2awNuhvxl+zMg5NxpCFnCL1EKix+
mTXp5nE42gYJpYKmIYI8k9YP+Oe6tOvY1gWD+Cspx3mUbHp4wMZ/1PYXoB+rUWPFR+Tjl9eJR5T+
q+pIFhcPnk5QjqUFY21sEJaXWgqmzwWAjPojzUx85kEeUFjE1m0znxrvxcR0DqzawIW6fzeBhee+
DTyUsitSdJCKCBevEqiDIdafexEvw8R0/CnLbL6D9eINweILIMtHswZogve3jTmM/Z+e8npVoEAH
/kf+Dv7/+lwTNmN1tTeZ1nKzZBttBUwEWLg6vx8482J0mQubqRi6UjxRR2JS7vYXgswhJd8fdo5k
WNCkpC6e7wwWL7JacSiznB9Zqfo26mnfFxv/c88bApVp1SkaDEAoiNjvC5wmWsHdc5HoxAl/SNTb
C9zG12TjPyRagKxf98zu+JUKe/x43VmQYoRhBiMgz05IwbQvRuOyc7YJAIb5uKQm5Va51o/zU9Kb
mqNIcaFlAPjdAeyzeupGBSN63BLeL/5tqVBuF+7v3vs0+E14olPXm7a9ry9iKOjEHixlm9TCOuhq
z3YZjrRPKCwyC1EYlHVLcfWIqOEUQZqxDgg823mbMIZBtBUPl3okLnwbrx5M0Cx+ZIYA0RSh7VUa
BnKSy8FKBJt1MU25g6SXR4cxQEVw4EGCoUaGj8nqu1EqDVGx1wduyu/DtnNpHXQL8YRNKVxKM7Er
O6FOz8tTWQouibJCwDSCz/WNA4KsYGPWbu93IxusGMGoL43OAabEqHgVSWN91UWD2iRVZiaNIRaC
CTzHDPVLsLuzzUpo6ACqmhQ4TJNy6N5yCesIN2aOJwo/XkXL+6PgiPOssBrTuEqe+OQozPAMNJBh
50nJZOzsHAXDcKNmLEmbvEQ+R4on21Zeg5qwVseM4dRXUwlF4O/uB6lXah4Jn7C+xEyjES/GDH0B
+tegILPGM6vmjJyb54x/pJpmQlQPDiVg5HM4kW40YrZ2ApkDVutFRfyBlvX7KDxFi9JIDz1gtcrd
Kw6ebippKPlMUmx2MaK2qZ/Km7VOvHxx1K9jSg78qp/ESxT7RdbYP5hU9gopbSK0uSt8efqwIS4v
STGoSjtV1VBVprzZdAwaubOc13HZi1kcSye+1VeeQ8kZACLrmqc3f7nM03EO6ixpLs+9/GbVnLnJ
n4IVXmiscLHS9Qie2B9q7Up/K2JfqJyJAJtsqbVa60A6XNr9gwCyNKj52P3Tw4g9NTH83p6T6vhH
g1WXclkSoBheQuRg6hsZTeCDBZQDee8H77suVEk1EtFTKQGsXw73klBT74h2TovS3rG5s5QU37EK
XT35zBHqpz/3M2yrcRs6H6Je8lrzqVCzwvZps8BqtKeSFpYTC0BhJ1PIbOAomJsyPRi4NazYtMcg
8FT7g3cmbmoAuAOUxCnYZl6ZMcX7XSfQ9o1heEjgRGpoZx3oo9T+WLC2Avs0WX+KcTLYK0DNk8of
46FNBBCItfaEJ4Z2m35pmA+ghxPfpBEtHuiel+qj/e9MZVG0YYlxnNHx2JSVwY0fcsmWEzZb3vSn
34jL3uKA8HxZ3isu8swqxBRB3qSVgI2PxqADDvHe5ludGQFORrNFZcQ5QmmSSxPKVux6K8JGaIvK
rqy7WrCECUql/7IUF3DdL+QgXpGciRE88ejsY+CTe3Qjm7nWj7RL0/2p+pUqyoFAHIM/W5N5IexJ
iIuG0wUJOkPPRBLC8rKeusJ0GeXyqW7yw5DYpgomEmdcWJ8JGqZM1Pw3xv4KUkay4aGenY7+SaUb
uhupn5LE4LmksmktwasDMzVX8p5f4X0lbesHjt+1nbmdu+pFkNNn6yzg1K4FW8BiLfs13rtIIdiW
/QbSbes2u2pXZLMVddJhLDNkqnrz1xu1LmEEXJOP7w/RPunwBstALG+upjuL6WAsm33KDL6AtIU3
P6Ibt3K1dTPAu5vHM8tUhSm51eQ0uu5KcyZOGJHFmedKNdn0dZiA6WYVsNcESpBhjy4O22j4Ef1N
JU9jbbfwVozFAh+CHfYIZ5C99RHdo3cXU8yE92L3PYpCKdxKx1X7LzGcyGtCGWY/H8jAUBHiGHoS
rse2Ay0hjggyr44FeB3F/iDQenA46azUgNO8BrYbC0hTROKPqhwCYHb/sH4UK4lcBOstubw1ZJbn
eCL+NQGZ6Z9NbG8X2zGPkC/gN9lVE5vDChdZp6fxsb2Q0G+CLpu2dBtI3eU0JF2wrXzoIsDZ9W86
uEU6+/z9Vm/+cNJv+AN/zzrUV3DkrDwiG3iybyzmlY2iq/hgPZoOaovTztZP4ejkNFGKYg2eNFcF
BKL1fAabSOWOX0M7qON29x8Rjivu8CU+f+ROOu8gxxA9pI/FofMpv9PlDoTgOvZGGoq2XmiWoZZp
ln2Oi8pX2WgWHablCWt4Lh0rKLXtdCPZzcXXzNo3715mv5rugQCEj7RiPr8v4tqN95vzP4BM0MTf
NuEUPAK+V3aCrVrVcmRCQvi3//Oyp6XRRNY+3ko8WCBNMObNVlI5WSinmAnzxa5qlQ8IRe6SVNUf
kvLbg6uFQ9I08k4Mz65nZbE/n48klD+bk/kmG+zn2GKGchhQjITDKaLqW+6bJLhP8+jNGzGPGEgO
+RtHViicmfXl1q/YpUdEe9/C+VFFY7OgxD8ZZ+dGgEH1Nu5sSZOZyg3/xdL4M4LQyUNDPiy94cAk
Pa9M1IEmYaZ3VbmRii4LUURp08PF6JcIogmT4G/beSCAoe0qT+U+2voefS3MtJPA7d2eKHpSr6Nn
pP5K50SeMLRbFQnkzDakbkVbEEwyihXzckygsWmp7K7o6eu/lmHOXBcCobkAxSORdpybwGzwdw25
GQ9Vb1zJJukwJdNU5aytRB2CEQD0ArQtciZasYWEW99O7WEvjPMabtjnnWpbYnlXYtI1HZTEQsbj
gl+Ae9ppPecfG+9mbJrbIEeLOw6FYdPkKdENbXbOrLmQbWGUv4xJUiFqBvA/SmRDzVrtmhMOxtwG
KMI1yILOQn5grTEBBfE4vQ8+RbftCZEhIBAblPhv4k8yAgU5m6QZAFynv7hysuy6hMDUQQWJQER4
JX8vash1C78DkS/dFBsAIWm1PQXfb7EMKgJQLgW4VY6eozMAcOAy5RSLv8mOolts8xvLm5DnJO15
EAPru9TRZPT+jVQUMA2K4tpJV75Zw20n7YSIUSbL9EqGIBqknSy2GQtWRnbriVhZO7nXVkIrBMWg
dcI47c+HdCt5ztxD1gqAutrOyDd2U/2WoMzNKiEWCNLcNauByK6rFWbB/u9oSlgPf0PPsbl/WeF0
p8h3IE5olSIqM1UV0zs8CQqA9FBW4c04WyBeI3dpSuNLMn/PpJEYhtFgTbq1D5QbG6ny1eQhQ9AJ
CPE0aldrWRN/Zu5PBVfnYsVjZAN7QIkS7XWXa/s9Ds7ox6x1pimFZzbJYgskq/MCrz5wII1zjPvI
Cjpsnc/gq7Sp+khtcE8PmVBLGhieVMeVyQouyMFYjEBQB49EDr3Z0sLe4eZQy72WxprfWjV3OJ3H
5D/ojYWhvMZlpNsJM60OXtXkQxaCjduV9hY8ZaZC3JBwR3mSWRwlhfcMr7VefDhUK3OCKWS9VTA9
JwivYfLH9Hpa/ZdPxvu8FfJhXvsKHy+FpLy9/MGHbgtJXpHXkXH7LH9FLDuLOionR4rhLsaD9V0L
ENQEljsk3vKp9yS/LdfNrrMn3Gt2MepBco2nqSgnFN92tob7hgqcBBZeMkeKdv1WO2Ohdc8wz95f
D4WZYknRtqpwjNO/irWmlYFbMliFOSFzWievtOkvfXrVyCFRnFGTVmX/DQkbi1v5oSP0Zqxkfjep
AodpqNhHwYP2S7KenI0un8O7uSWcJObhZS4DcNjB3KmHRN99sg6PqFt4ai0KIOFOhYBv0IZkwdZz
7qJX7KHu+JbE3ONq8QzG/vNaRwl6X7ZJdZCAOYZ7HXuW3OicEjpVEN3Irgn0AAzvid6Td+PuXFFs
0lM6+TBCGQWzS9x2KdbZsTZLk9dwPqy9zqYCfGaleCBKMvUwbsfTgJn7jCQDtnzil0mlWTAHcFy8
+BXpBqNMVfmXdpw16TSNxkaAV1v1JsTY8JQcJY8jPfNxEmZ5YeDSV5FPX1eClzyOdcUabTRhKES3
jzTxsYWMuwCLt8gsPyCGLyxM4cvb8exh6R25WTxDVvSH7961TaVzhcUuxM/fQAJAgL2gEY7E1nbn
/nnd1FFOhWnXdANZu4D1bjig7+ceMv0wbxigAOfjo0864b4isZc7T2x/riw0CbYIL7WguvmN2EYD
LN+yNZAruDw7Vnwh3dBhljeaqayyRjtViBKS/URc6rYNd2eY7utNxmeaNeM7F6cTaq1308lZqEcZ
4jFS3aoSipJer47wnWvAJhU9f4wGXW0mD8tdriN0RisyJoqh5EK7aCqvlsjIN3m9KoIpnXtS2zet
5PmEiJdnqtKRHT7avx7LqooNeEgY7e/tGX6VOQ7Ukejoznj6EbwAwzYWJ0sTBw35PNPYC29GRJZL
xTZaytkImzM/p9VjVHofJC1v+x6imb20v/wpjcz5gH/Y2gFJSk7DgCeKOFymBw1VvGuyvj5xWu3t
EEqPK5KU/rtz/PCsGB+A/jhGp6d7ujw9k+d4X3C2WIpvmp1CHGnitSc4LtueLM1cEgEWWBf7GhUp
37EIEty3J/sVIunDccU2HCPjLoBR28HvKPsr+3DeFeG+L2aCjFDweUFtfzztRL6A2m7ApkxgqMGE
vNwFrL1hv3y3wdfFcmpz2B045ELwxX7QjPGIaYuadyU3Rd7W3yHpmEYJk+ekmSJgRK5iQl5RK3pX
Vx9yFQJt84gIvSjOtNbPCIfffz0L5FMUR2ZeE5nWUk5EPQwXt829R7SSR5rPYfYriEmrrqSw2SFf
hKYBJD6YRRvR9uDb1+z1wPfqV031MmE6WOH3eKw10ZawM+RHW9qFjjVPadD8Rj1VsJikvVn311MH
hPjkT9xFFiK56hXs/9RA7miqloNiKvwjWHwm43NEdXT/bMBnohGfoYJIfD/W0+0p+zE+tYnWF0mG
mSYX/n6Y72ctcFWcV9H7OrGJwHbreWyafxqyLXQ3lwUW5mLp9IyhSDXNu5cWUwfn/iVkUeAPL7N7
2ttUz9ADQYMaIuBMr1nLUjhT8n9j2hyBvrk7JTIf4dMfkkmcCJFloRcnmDYm9nhgNnv3MXwC7B5h
eWimj8FvWg2webiSZOpVQJZ83DedbPk6iK9Ws5qnE7Y1UF93788udvc6IN6v+ouhsV4EwZigiNu2
SAIIpHyc6GNGV1ex10CuygYqehu/eTWOTDbwnb2eU24NUKCF0GfT+ttyc9v/pHecC3/DGuwrekj0
l7L9JRihiYTO+KPP0nIYiHxvIJpQSPgV9wPGYn7u6BhQOJQ3sFAZ5ONoXqyxsEaVSMCuObZ6DMq7
IEZx2uKKLwmrynn4+jNOCA7UczT1zlfcsuq74c9RoAY9zx6ehUFLg0TAlKePOgAIUZk0tCnrgscx
uOq5fjaA2m46CdW7FhKJQnJtYaE2JoGq4v8LOCrc8/+pwEk97xVeB/K2f1ef9V4/+Fzgy6fqWSPp
bjEMGjoxz2G8N/8d74Y8wt+Y1FFGVgadXw6cCabQxIWqC/BBOV6sBvoFKkOdU/opC+gByDL4bWCK
CBQq2j8840vjUkkOFeReRUAfY6H5XBmJCYhSEe0lRXXp8lU1Cvek926LIQuZ0E/R4g2uOzEozzGN
vK1NByppue6/szVXKpSIPS+Op9d7FAJMhaa4EwZQWU1mjOpBegg2aJNxHpI6p5PzlhjxnYftHoXC
am79GYN/s3ujvg92dr82HqsNUsE+FtFK7Ln8ILFFenmM5wxcqeGd3XqSUrqgbVXib9QRMWrHsCSX
r9g8HvqyJxYOSl9b8+HNIFLPOf86+oZYryAzbhE6KOXDLOgwqtv3dueX9a1tmPxyVGgzFxUkl/gb
9CWzqo5YCNy/Iha09yi8J0Kv+zrM4EIWBJ+26isaK+5XfeZKCypx6WQSt0gCaph8pKngrNjQ3x0+
5yjRg9yvxUzBiWnbuS9fi2Nf434tpY/jevyYpXb/OelsKWqrkX/qbxKk5dWAiqXvaRzuRkwWD9uv
LSpVOSweIYTKvicd4KpxhVAuZR/HAe89rZSm/KXqANJqP+8nCnKjUoiqfJtkFAbVMnzpb3cVuQVz
CPUbESAeNK8y63AfCCwZxERwENMyeOkXKbTQcm/j/2lSBnxSGMasx9BreMpwgdTVEzc1Hc/AFqfV
TGlqQDi0vLBzbObv6B/IQdfs5F/WCd56fxxwnKkaxwGmlEMpvoe0jEWO7fbJinETy9HBGAROtoWP
eYnsebH9SaYOe7gCPchocPzQZr15QYeBgQDiZTKJYtNTq6/D5mDs7PBd52iLZe3BpWZjqBVW6nx7
jQQkO48BMMy1vHZLWzGM7jxN7a3HRJgy2/VpfVTfrI/N/LMVghdDkgo/3Jb87qwRf6P4ozjDZ57M
q1wTFz9EeEaU6b7hf8OISN+ampnTO0Fp6quGViMDaZUGC+wTNhQT0Iv0FB2LCxEFuOhKpyWwtRP5
eqRADkCqFwRUpmS0OBQO5kVPeY5wQw/5oWlvl9lERoWy0ws9i4q+SFgxxi9OHFZfcphuMwUQA7dX
VqZk8Y8YiOPmq4ox73ESJ98uIE03Nz50quEpZKCC6/f01cK/0xozpNejdwUeJVJapMC1pavSw+L/
NePUixpg5pwJBp+xcKWGUKSSX/nw96c9H9dai1wMYEvECUnik00Kk00yQY9TnXgcdd9UFNirxpdx
6y1pc1AQh7DuFbiCnRDWcKXF0+Ecum4dIrbxkJ5Ebq1v+cP6obj+gV24Nwe9DclZB6hgm4c9MXgg
A9LrgMrkdvKxVQOoMErTXdwh0prdoPh+adf10saPClMCveuHjlwPlZbIbztyR/M4Fp4Tk2cYDq4x
/1Stvm9ln763c2wTy3WUeZqE/zLc7LWWZ2m1FyL6E4QGpfhULBoYIC9ZeNaC0CPcQojOq0oNpqR+
Id5fz20rHoHlh5AS6+vH3OM/kg7pSc/XayDa8AfYbTF9F8UwyVyt9IyzV5UICN/nfhLQD+oU4SpL
loaNdEazSYRYoz3hszGy+mnm2YcNk0Y5xpFGMdGrPxGhspCmy+hAFPUu8Ygrsm0gsjzhmYiLLc4i
V4KIrm5layTebhUWPwuzrtkKo+UsrNQeA1tyGv9xuLedCcucgwf8GNFvE1RWLpsZYsUUGd1Lczuy
2vn6gc0TBWCrnbqLvjGsX+dsaFrtv+61O0HblLeEdxdgu92IYpIHn1tOByKuV8QM4SbmBYEL9Jez
74WAuuN0WtWjm3Rp5VDO+xGV+u6MsjePj7NgrO4CU31XRdomubuR8HjoVfjT0QNQowuB7AZOw1UM
nx3CFGnqHOtPJv4mGDfacVM7ezZG/ghdIRP3N3IkhhuQ921CPDQ6oTo62OcOYCknSCIbOutFzF3H
+ieF3waBIPhLyeXxzy9J3KLaXoa3eDNUXk1KlIFccBHAyMNRTtpA17933ynX1tHvBOOkU9ICawjl
Nnvm6zB2hkNynoqWp3B2MLXp03mOXzJi05MxFYJInlqRwzgPqf3gC59HVE9++I1BhjwAyG1DB+0U
lt+JXVO8dM4t6Bnx42es7uwSXRYgCqnLnZ6oqVhWskWemOjcFxX++MVCyjt9682f5VekXGuL5Ca4
+TAKpXGG3af/XBrPZwNrfvWbjuGh1sI5b6OcQ6+HS5URqMki4A/aVo/+YelZl8RoJpP+yhRkNPVc
1LX//3P2aEBqngH4yq5934eBOvHBgzcltc2uxXjy1uL/oCtdN4wfv2fC7fFThHaq0h0yqRipjzQb
5bGebKzN8pUhSxU0HOP5oLnRJLxGo7O0FTnyH/Vqi+C8tNvgC72q0Zwmmf87CXxBauPpVe4pK288
OvwHhM9zgjJ6J++Y3Z2mWXRQjmq3vED+bZCd1Vn70EI7PHRrsAjx4O7uea3ldY17E8ben2kr5LNp
YbKI/71wxno5HTmI/YqzsjRvmAVE+lzypfOyu3ES+q7+h7qbU04k/mlQR0feyE50dS5ATIiQd0rl
fLgh/miuaL6onZPT6RkG/TuLuC/o4YhxZveC5y8X5atF09QM9S1VCY2MH7Tu9KyVvwdzsgP9rJpX
jCxnQ9axc1a8eP02oVz3UuZu1fhJw5/UDzu7H3GCv8ybZ2TWprcW4WtzgDvAehUsn0n29p4STHWp
wVafyhQ8Pk9w/2oKzeMcML8tantPFi9CX4A0h2xj27pRrTuo+/SHkeG04TwXrw+pQx/D0mbKfv2M
SPo/L4mG4E5bJpymfhWy1tZtp/bNpUDzniHpYp+nyOrl2WuM18Cacau3jfdlUg5NHva5VksjjXU0
Fq7hiOCPSgH1K4bLX7Uk3avib00Imw1pFejM9xMfDtxJ5uYpcaORqN5FBqlC759mc7z4bWfOyf7d
ZomlbqkObgXuND4PUmsodQi5vKiQVbts5FxfyZb+usmEFsn9wOSsrQ/yJxnN/mzVjYH+MEJMpYKT
u9Z2qsKmrqvs2vUEbp6K82bb8LWNeSmkHgVZjzQ0LnsTj6YAL3UXvRtF5d47A/UQ9erWMRUlEVoi
j/dJVtwsCJr5l/sIoh8ZqFkLFMQHSCHoC5U/w+1kBxgZQn9x87a5Es94D1PS6Left7md44Mc7JG7
dvQK9aUMJZd33QpdIw5Zdsnt36qRy6r2Xuf9KUBUv04SFIZhnsvJk+5qXVQXTjQjeTASFvgxTewg
d3rNRFxOLQfEPFQa+h0/8doaa6VVITGtbI4Pfr/YMDg+4xWx+WZ2df2qOQFUO6JuakKH2NoRF1FH
3Y49Gci7Jf0ZeS01E5FdCDIm0BvfU6JdQ1ZPFdJVfiHjL6sE3egf/MRuEPG9I9/j86Eegb+oDJMF
nUWJQsguH6AGmK0Sg5Iuov3ru6gNiiSRorhE4zVGhQUw7KLJRgXyrRZ7B5xAAgAkIj5DCFyKEHGN
YqhSca47xGkP1zV7sqgQ96KOkBKU++7XeDb769+pUEnfaTk8faWfsVl+C4EUz0wohEXBldT+Mr73
hfkzIRb/daKoz3kFJE8gkAS0RZag8ysHQSTteHeKCOWrhXcYJ3Gz5bysirhjHhOZnJYgC6S0B9Az
pSZ6A6s7TUdrj6Dths5Tli9iLgZTxOteWD63Yr17M4RKx0pxn8E0ul9x5IhPX+MroI52RlSwlVaq
/OaXhH2PZws8lDY3SkZI5EgUn6zin70LdBQYYK8mVibTVBD2VgasDC33nioDr74xN+9vTyMaJMj7
NsdTYh97OZz8rrFeKO7RjZlcFzw5YPtGo353/v26a8nnzcrZL/wj9k/6bsKEtd4nFUoMKTMPC1VA
YmSPtVdn6o7QN8w1U7BLlYtwQ/qMIT9/9foSiBcK9yG54TvqGUgtoj9+bZWasH6c52ykP/USg66R
OJOA3oo/rksJjLFr5kf8bQ55Gfza7SRBLU6nY9ggWjGbqIaPheU0ZCfvEjbfcnJXf6qeMWZEY8Gc
Xwtg53Zi4orRqELJDlekfKA8ZhLRa+7eyXc+v6ygOkrLGgdsLOKvX2ebBXRVdI94hQZCIX8sLdul
ok1UI0nYB0nLmw2+EKPD/EY2voo8hLfuiGs01gH0L/rkB9oMF28fqqv5KKcQPEzJHq2weOWC88Mh
uCJaaVe9MJg8i5QIUpu4ejvJNVdpkAFAnsOc8akMrNqCAMbjDD95f4E/dDEihVRX9RhsiEB/ch9/
tETJJRu5/tTsYTuYvASRhRanRYf4ynZ1/VU1BrlLe+8ge9pyF7XDz+pVB6raC915ahlT1NigH+o5
vvOJub6pFqgVrSUmqCcAsX1L5aL4R/ka2XEuRrc3e8AyUCfwLzwUyDtIGVIY/IxzhZ8BxOuTZ1nE
c3DQGwySO/KZqs6N7IF9psTY1bip8j4HTxF287JKaSpi4BOfK0G2BnnL9bHlEp+z6h1KJBRQ5bcB
kDU7qYOFxYrgRStvFz5WTwp2VIA6mGkIOqtduN3o3Ox4eDkKpywn3/E49u3EHmuFLpue5g3cpsd7
mos8PXBytumRaSTOy3iWfN0IPRHCmm+Ad8WG8lQrOb6Hds+1npiCiW7PMffQthcvnBNvmSN2+mou
gS5ICYZxlWk33+Fb1UlCShFoGdqCHip18CveihaY6Mkr5MLolJ//22zYGICWaTj9WmmTwkBsIL1R
Rap01PrmfBRhaIT9hcQIDR8cXvygVQQCSUk/iWIEZXqxpdp9t3ngi5nERx4heVmMiFyEGt84J6PA
sEibNXiCgaQMKUx5mEcyBB0CNIN4JMLvbrxQZBM0TFMUmeIe3wRjxwb7pDDWLwztE6XPMwm0ANz7
mb2A6+ej2cFGpVXCV2gkmw0SGfvts+Mz9MFUVUXSvs9z0HDdE1U5p4SRD0ozhPXTp46e+nDm5bPh
sRFT3rNpR8lxOgwUvuDvZiNbAUuioGvbLl1Pe5X3TYOfZTaHkTN3IOvsG8eiE0UeudJ1CgI/ogEV
+5lsMzCJtyhbQeEnuo0LZCdPMfRIH0wW30wGzLWnprn9xlOxNYzb6VRiyEGea+4WxNhv1s7o4g/I
AV+dzHDzEwnjHsZ3aS+szuaq05XRJqiUkppL80pH6Ra3YvgYngCtFq+lKdJPzGFqkFE3EauJ7PWS
czA794LZbItV+gXgbo9Qeo4TuGFC+ieRrDKxZ4pCkgCgRXjlbH9Y0N5ogdYRT6b7AX3OJ2rKVYyW
CiTCYhskk0Ckwy2Xy7ZILgZb+CUoCC0ac9oRbh0kSE1oKuh2jOgMi9o/Fa4MlHVF7yz6rtHVe3Tw
LgGXVefrsHb1b+wlQOyGcERA6JN3xadsfg9NfXBNACHt+zBbWl4a4bKlC9bzZZElNwaUV1i1vzYP
18pymCfkKXeeRY4EGGIS97b81skfPc3KOQu1jfV/3FpqlZrjRVM3mIN3PDOoPD8KPH8p3ppTZhhM
dmskDixZVhF4/7f30dGED/NUAwid32qVZlHnqIzYLaTgW7UD4mIBuh1apDIcLZDNA/FMvcirn3/u
sHTTdfoDo52E4e48an3MQjb+Gf88OQznO5jY6rC5tJyJx18+PEyAI7/tb3jEj7QchiRMTFKJNLgB
LWOKxLB5G81BSuCWcwKv0LJPtQduSurmp6M/o37N4S5xz10th4zHcHGxsjxgGJGYpgjkIp0/3pWy
ktiuF9RDwlAA6xnJZ/jZTTuicXuCTirNBkK9o8ar76wN8BsYWMDVqZkfox4vRgpO8n7axw4A8gxH
7PUq1vQOmlTykWbuk8TKQR8UBBImXRmMzS7qWc8+2OVpnAQ6pmr2SfgC2JE7khU1T2+uAeTDYb4x
Fn9PNbXBOKU3+ShUiei6tIrPrSWQW5JSfIsH1I2upHMNuFn3iTIgOjjknD7ljjmkrWxM11U9sZEj
Wuk+7T6GrhoS9QRYMrhwAiek1B0sFTbBFRyr2GMum+aaNdmvUamw0LAT3752olwDnrm1b1FpzkTZ
JFtIk4my41UtlfHXjTw4Z0/f318E767oEL3IuyMPDiPf171RRJ3rkbMEeVYXsuLNh8SZ9kqBY3MK
rcfviywhSZB7FHKN8scGsqX1mZACf+Hr76gmkH+QoSuPNZfsaCrGG5euf4AJKONMNEh4zlzZbxjz
1aHA932wKIPCB+hkfuVm0FTv5heo/0dbZmaxScpLiF5CVDiJD86Tken6DDTjGCfNyR7Sl6GF0Cbz
eCnIb6f7QhHKK4IBRJWBNo6gzZVTIAt1DKVd3k39g0QLDIC7GFhRF9ViD7D5KNMgByXVBr9p30bP
5QW7b3SjxLGdoNtIOSenAdqPaLcQHCRScJAGiyn2XXCuwzZMIsQB5+T4GKghcKdii2x52sI1MLIE
KnIqFkmt9xHEQYSDDR95UODa4HeSjVZYTk1RMqoTX1TqnHhdB9NaR/xg94g1aXhacYw0Jmq5WnEk
RpO7ozMW/cPsU3mMtYRARvkW8m2vtU8qx5WJ1KHN9DaOtKBDpAvQaF3yenhWv02ybeuLA9YMgRY6
qwmtCpWVizVk9zGtT4jx8uyTthhrcxDAP/hMn2pabP6eNkjKcR/cAuH6teiU2NwlzNSwv0EPuu43
ODBtzjcuQuPYQiYpQPU4hzgIntycg4CtQo68/6Jqwmsv4X5P+mlE+gzN81sigAiD40Bk8fIxzjsS
i9iUj2rsGA82erJW1yKZLDHeep1gcT1Cu28VbR9/86DH8W3G2tZ9TbkImEa+ZAGzbeFpUOYBtrI7
yfWrDW6zR6+IwFBnvTugaximQFveiUE/QxnwVyH9lp/4KS2Cw2KTyr6+4kEKF//9xF/RFsWynHrc
EaFVtzgFraXB634KLf7m/Hzly0BBZlhJRa44SyaasGFgnmhPHpLJd0J0REY05OGDCnr1nj3ySeaO
oDxwrAgi7WjH2CmNYurn3V7XUgUZFEqsOFqv+NyvVShZ5Z3vCkRdMbAkkuwxKNvTXYq+VBNvxYIU
n2/M9mDWKtgMCQFo+TA0cD+s3rbODiisAP5Y8ukE2ipPjaTq5A4qBcHfr/0GhUcYQmpzyWGVE+Ok
zPIGwYH0Y5kVr/Y6HoUPmKG0QH7BS+Hx02PpHcQI6UZ/HyoYcYU1HwgOBPrF/vILZHqT/oo0E39A
sm04jYwTsjOMdw+MDzHyCtlSDwP63iMiMtn+OsY+D/ism7HTKcMFcRL+q2nYvS22zn3fvMG0dhxE
LHWUJ91YIpyu/telHDwzBgq2T4cRAk1ybXKWyV/+cslkgEnexRklO8AvI7sQ7IzlHFJasIguaaD6
VmGNDcgAARwPwWNc8uaJaj2km5Xl87ZYhu3Lvcf/C/jz9rAkUCzO+vDIG2DeQWkBIIEURYcxVcVH
65dN89BOoUW41NvLUeO7rgETLfLWDScEK0QbGMtP3oA3cqvbtEktoYLDFN46pDLzR1JPwE7TVyBF
ImUXopjonATrPotcolgLiQA4HKS3Z3wHaOB7s5Zl2BUKW4vdHUjdp3fM+5SyCEYY1LCbNiP3aETh
WuAR+kWqudWQVUMejghuRgOF0zz50N6XGsQ6D9ciAfnoZQ9ybqUU7eD4WdF6e5RhdKzz/o7reT8S
rI3RzAPokGNNoKdOkaCB7pD6FSEEE3kI77hnoyVTuYP/TfVNREfIcBaavh1wEr3FOBeS3ZtBBfHJ
7Siw4GVi7mi0IQfpIYgHGVIJhpjgcrbtoDaa3RaedJgf+ZYnHE7qc2xMYQc36wk24hOouFd4PqLN
AnuLQtZHLuI8m58OhEBKre1ClU2FSreXQUGpGrMpENycmSwXLANX4fQ0D+AdaBNvqL07/tsi89MI
cBVWaiDkYw33WLup9OGMIZ86u7hJ3FZdgH3ZQMB/jMzIdrvG+I618AZfiVENVGRZa2rYsMMupmUY
ygIguNK5SvP2Tp69zqLuGsQjM4/vq6WV2Eq9jL8BnQYTbRFviWousokfT7qPZdJ72dN6vljNoAjM
TP0zPMbuiHclyFipy5pIXLkWg7hGZUQsSsTt4XBH/QVIEzTQHYKAVxvP0NjZ7BqrApn7+/k7+LPE
Dco3rgTjamZjRT5Ko35Vp9owoDZqVacIZ3XNXlK7kuQJAl3+qtSOC+ujCmuqPK1N2dUqn+ci6Fw9
PlfWL9x+xIbql4oG8N8HFCTufpFodi0bc52SW5KiHgEUZdkdXsudMNZUkTmBnRppXTNJhYVimbxc
Elk+5c1jxNqEwRyTUKHD4hSYV4Ejp0E7pwY9ZsDDL2RhabdE0N7PjsDsii3vd+oFa3E/W7BsxUUp
cqDbEv/9QFrLbZhT1XD9K6x8fynY0vb9aQGJnjWNst9GsAnbiDJUA/ApzLlZFmnl7hLjNlHuL4bV
zxMMvBQ7pcbJ2e88WbXH8NDYdQlczSSCq8zzvFwSPsdpCEq57zN+aGPvr7stX3fUXsJKg0FqK5gt
+7A5Y1Iz4P6yKfjbvsxcCYD5D65rgPfD4DAJGkBDjQcxDiAkUt6kMsVMn5H+VEWPp5yW77KqQxXP
sDdsaISjsoK2VGA1sNcf5YB2ExqnRYnA3ke4+AJveUxeAY0iCz5cZSnSvvaOyBVadhTUd2PW4AqZ
8PJlsFIkDUtUUbdw+9060bwpoIvBRpofisyiwMo8UOYObI9ZsDL85plfqeAzROQblZksIop9eyGT
lTzIdWvXD8gaoI/7yMGvHVywjudkeJCZuDO3peGwJfO5DW2roxxm0vpSnka1WjuTC3JcXeJNb19j
ClcMxSi37fXPnX1A6eTWuP8zFWr3ZRI5UXxa0sXssQ3XWefzppvfgA8SfJFZhwDh+wFWdTc3HOc2
KRzJLNUo8j1TmL4WYd2eUQU4ghxPlvrU0kMF32KsrcsojcMLDZS9wrXj3nz6wWpCezGvG3tCXsCm
RM5mkgAEJPn07scCcdWN/c3Gn4SKncB7ieg7zQhsahNXdpmOjnYPhPBVwuhP7o6bv8jfzzhiCFa5
P8LgtTGSl8/Vt0dW3bYATuHfIYBKKp1LinXmQVFOjiy99/M56awVCGR9KoPZFKpSZ3A2NrzK/UwW
r30DgUCASlgkr8Hp8F9KpUly1K5BxmvovbHR2yQDS5eWEso5M7qRvtvsFmhRy1Igl8JuwVbltMmZ
rC8XwxVNbIglQfBrNV3npniAo79qku2jS6HHz1JfoPRpVFElA8e3ftsXTI40O1SZqCLtf0Ex+4Th
GVNgcnIrz1ejr2wZ2A1Ckq8zoBgqwpSGie2PQaT+T7XOXoyio3AvS+AH3+mKbw4fDHavtnDToPji
PzSuR+SNBj9cv/eaGuLAq5JaX9hqHtEzw4uH1p8xq0nBsdLIDpfbCaLYa7ouHMazOP2jnkOZKDw8
aVWyp1hUoxlzbW1VGUqUhtsItwspVX8GyeEpFAEq3SHpbeFfpONul+uBB9GNTzTN/Cu3vWdCCE23
NganQ+9UyYjV627MuwP9ixEMhszESOQnNjtlS+jJoQDcvPug+zlGE2f0RNiGPO1UUODNtywj4t9R
FtlKPcdWKUmpXdecOu3ez6Cyss1GY47U5B3W43Gnu55aYU/23jd3xa+hTbseCyYlMd1LGq23Ax6y
vn8E6EBjoAzavDA6lEu6ceTSwg7POYOwwQAKN3mJdi4cAULOL+dZot67jyugKsnxTj7U2jqAGpTj
QqYWaB5M0E6GSRoh8mT0LXPuc8Vpk+QRWNNjRSAZxCKTKniWqURlWQQOFTbWM5FNrIlEvDYvgDuA
YLmVFuZYGZROx7ZYyQ/M11BrgTdDvO6cr9gOO9yT1OhpP4sHo6IVWqiWTcCQ9aQmnS2TGGKsbC2w
OG5hoTzn36BRnB84dsVPiEkBV8hlxU2l8W0Ku1+/UwWIW6vE+G+9e2t+ZN0VBBMo/q6ajMu3qqof
dcg4IK5BF+W1gstgNmSAJ/mCzV1jlgySPpVtZm0MI4hZb7tffIfpXXIxYcMHMw0S1whzIwqMzdQK
xvveW+I8pTvoVnCYT37wUivKDtjfoiESF9B3qCA9l95Z3vyw/A75hLayC4gfeo/slAQuVsPbv+C5
hSaBYJPV6fwwX02CVqTZJLfaosHOr1UxdXmmoFQnCl6A/gA7YJCNQW+R8tbHY7YisGBAmH7HZ+yf
lWZYw+yhE5CZNQi5X5feDIgQS6XEsugDFjLJV4aOMSFN6HUZPyO4BUaCi6IWmCnaOXe7YQSSsCKk
3pYZV+8XY0XoF6nR0m4br0YcJ1BbCX+6bAGDnqH/pEaM9RjJbWl9klx0j28/8NDqlaoo5wKaO3fW
S2nJgzA8zr2OpcJQu7348GrfdeUprhgPqekXOzgyWmPShb1kPuzq4QI41XigHCtYMquvgP/WPrX2
CldUsnHoqsOZ6lP46pV2deqo5qk0Y++ZZCAMxun1MHpE5CLlijcwzep0Fz4une1VEhGEgxobtdLM
WnJ8Vnq7lvoWG7YT4vy1SkVy2uzNtwZ4GMk25bD1cWF0KRQnqLCVZYYiivpJjls6wJ2aBai3954v
vTvRyAri1wUIoJcGc53C7fgLVr2w8y3WPY8pgH4ZYzN8VA68BNriQ5IHDUhW+smo5FeDwqVj8S4O
vSeDEL7mYD1X+5wYM8SDLiiyqsD7Gj0IKlkjOFup5DzFVWSxwk4o/sKY7j65RYUJ3BZliELiY1fk
y5fxwMPU356ghwiARa7zUrN1xTJoi/SJl9BU0FExzBmUGFCOCvkTzVU40dWDxGJ6mrjGbufTrBHP
PGdcLO4sGMrUEquq6sKHNjlA8oaHuvpwJ9bFeZw4ZygY+KCW3/ng36KqM2/6q++ZT18fVDn99jiC
7mNnrqPHvA1SAWEpLs51LRYTaeWZDy/z3BQWya4NNAkGGIQxHFU2i8nVgpF/+DV5OR2q7GCKTSek
8yNM/PDdJC5L4m7ie1wLbWOGLMW0P7ICZs1weF+pjGlyJX7Em7CsEc7J4ko5VefLzJ6MWIpsPG4/
LKXk9C44BpCwMmcVFHlseAHPScyJXgoHATfddjHu+RD1djO9pZ/+PPdR/gxAnCiJEoA/FPVdWA4F
BbUEakhaD/Xx8W1Fv6F4lMaxKcWfrn29nIYjjsOMyCfGS4AVRQeTargmurSfi4+6RABulkbKgGC/
bTZ/xBtth/RImtQnLCpvYHtmauXpCarrHiz11fDdFLDURaYeFGISKn+DcwM5WKGzVZkwufLsMU3H
WMWrwxxKlgH9IetVaY8HCteBQA5NpnKZVdJaJJ8U4Eb+S3f8UcKqlseoTvSwYE6/gu2/3sznAh48
SmOXhg/48TK4GM/n+G6mhZUQa8rgMxgeBCCnn8zSuZTXiEem0x4xhHrNJ9zeqrYhIRFLSieZpEdN
m3E07MSzmJxKlHh4wEg2m6BapIGGnT6gDwOUOvZ+KBJp+5MDhm1twKZq5H42F2FVe1J1NbBaat0B
J80R/s2ogLZnNJ0C/bowY+aYmvokAskKSHWNeXaYtZACDnwyID8qrQZWQsDVeBvPIr7qOXA9nPhh
eLEVRhu7PvLjoswyraMV7B/QWkaaU4lqRaY5K6HROORXt6TSwONg6Zp8Tgy/b/Q/4o6/TJKD2p/L
3VG99iVidGuBCm5Va7K4buQN7WHrjbwVPQf1X1Y+/K2vnwWkriYMQ07alyLhKgnT0Cztq5ZzimrY
9RsFRj4RCopUALSFxcqXE38zFnB9lwAcrTol5xrTtj5QXCPIVzEZRUlkmcm/XEev72tLQvpaLV0G
WGnnUisTO8ibPz3Bh4ziX02CoJVojAjEFcMUZqD+sEcjh23XDoQRP+fHNoITc+SUoPdDV3Uwt8wo
E1wHy5Lu0GCbxff3gWC1hOuTv99KTnUARJ8cAthfkYxxIrztqzqQ8D9YabCGdveMs+fYYMqasCQJ
ToJiOK9KLh4Z+dxujaBevEycOczEyoymP77t0eK9xNlb6u/QYPsmn47R+OC5ptrY6yGm5xRj9tLu
Mr7RlN0T9qWD6/Vo3ZGT0r9RLCvTOknytnA9xTwAuZbnCoUQqgqidjEvjVPNAZd4NnIEPdGOrVFj
Nlnbwn88rCmka9z/rqF7Vp4OIv9yzmUidSZsugiVzKrOIeR84YR/uf8QA+wuhlt8t6phrisAwBFh
aH3E9aTzW3wx5GYnWc4N6L78EQ56q4VWcuPsX7AXNarIBKoqmrF8sRCs2/DPxsKTWmLCUsJEu7iq
dKkX4WThyBMWPeYA4v4foh0X++KEbYnVrJuLIjdqQdfuXgCAJu9AN/+UcWH8wqMmL/jXAjdBrYXU
SflZg0cXPhmg0zh1YZbmAB/RK48m/2dXIbrWwsbPyTpTNoIuIFhNPDEABGXBhWCbuNcVIMAm9aAM
yRuKDKUyH5qaloygjw+wHpMlV2rTLaL5Kz+WiphLyCAnYB/pm6c87Pt07a8MwGW5OSVPsW0YxemC
lnjqeXYUxo11pH4uoco54Se15LT8w7omebyunzK7TpDMcDtobBlggUMI4wIXo/VFhoEUXDgjdONb
ZNo/nInEOienWndJiunqRRL6mymfpXuRtlR2V3YWLYxwjUSsrsMlh3evXISVzNcnncCSHv7SX/+M
j60TNR35pAigT0Q09Ws7PPHN/CX3QxVCsfEsW6oZT02DbMTcYTlbzi/4eu51mVmSVsv2eQiQ3M/2
e60tLmbcOEKp0daoOd9Q+01es2zoVzMnV4cVJGuoBthA0C2V9kGlHGfc84YC833fPeM/JF8Y9Y+y
cfA6oQf7GWFNmh3venx7VF8ezAbWGsOjtWpVQSLRZUOktl+cjd1eJEcvxh9cUTATafHmsGOVDNrC
OhHL8VeC+c12iyMkawbWZ77OGuWtt+YlzS/CAGAXXrKDKqbgaUnO5goNa0tkFzvgym9jphjZ3e8h
QLmaQwWEpciAEPCpb9/yB8NQff/0NGLwCN9DllWl/KNh6LulmZezNUx32AAtJHAHuX3uR10g7hrV
Xp3XM1/h1N64Bq3HyH4a2IOcgDQLAdmkqKm4QaxAEXopCz8MK9tsfR/fvS6VaD+iL8R0SyPubDd7
FidjaITzz94EHEJrDZnssCH7e8Kpa+hGb2yvorOfaJxUnmGnkto+cLVnFdOPmOt++8bOCN1CFcSG
HTvHJJuSqxbFessHa+NY4HeD2KaSggf9y3DPAes5U8zXj4UoZUxiBM/NLwtqf9vIkm3Q6/1eId6W
Xv6J9k9x4GkG5dQOd6neyfnOnTMDXJNrDq9ufp5og2+69IkHxlWsUv2XuHhfDJFtGu0r6BivWDlY
xtk1+ox0Ky8XAzHf69i/7MAnYwQ5Pu0z6yv/sBs9/HJn5j28RFMLQ50Wa0w5QwxF/EgbyfcSSk0S
LGwUj2haXIjKOowtbg22IZJz3CYm8cAOhkjZuYBnbtP0XbCH1cDkqPJreRDe1C2MhBULU/omLznk
kDQy2h2wBCwrcfBMUfDN7OzEFMGePnksQgotgziXJ1/rDLL5RXPZG0QIvt/MCTaaGOu7B3UNjL3J
AgmlFi8lLTYKzWUiexVk6h0EEFk88EI6SZDI4VZNtH2TzH+oKfeMJxw1Gz1ObIDfBUSber0NRWcC
P2vx4nQirgWtuyKxE2cVnvH4iFayEQB7Zp6dMzkcoHwi0lopWvUXh9talTvWVyMN0yrJSKEAj92F
f/BW7+YV3/RXMg8vDEYnsuJt85VZDJSyaJc6i283NZogqViNl1TlIMGJvRJoQsJHOIApBZlYD3Uh
Aj5caZN7UaHIK9TJQj0zRDtpJihR6aoq9MY75RKVwzGlzLIWNbrj41k/vuVnSdsBSbOpN62051sf
53VcQgJC19PYuly7hLCwZn84Pd8Y5MTAfE6B7W+YgmXlymkFq04Tc/L52GVqmuMh0mPw1vvGoRqH
6KdGDvBfWJYCuGY6CT6GDBlOwSlMhMVeyrfEoSLEGPjTWIMM3eW9yBWb6CHptYv7IqXTBHDyN5rE
ZftnLABKFdiNrilVtQEdHaYh0QLJDVLkQb2nESCjAvTspAmTtbdKTMQEdIRazff/BffYAciHwd4C
wJOpe+XTNb9F1xGmNhKQno/r6QTKUfN+/5Ouc4ttiyJjeM94yOpvDCyrIaYpqQsBOh6Y8iMktlkt
7AOxubhdgx0mG9yM645rprzSuMMhQ3Gut/Q0weD8SVnhmVq/zBLyd/cJrGzY20G5CykLwfLH/RWU
e9lMh03Jp4aXxPrYr5m0QMqUrja74ysXfy1Jg3OX/VmRadSim6df/lzYuAppIpbYLbX7YDI2bJkK
vJbSFNB7jyZC2F98FfqtSgGXr7dg3JwVIDdmXQzIf/P7NciO8fwukgu+d2MdxsZCUlatMZQnxcEU
iv0narMmJmb7Q0t6q+dJueTXRWYp34ngE2L9UMOY1fbw/LlGtvL9qAh4Xlq7P5OB4R6Jx96fNzcZ
22b914xu0ofomF4SP4WDTSwJlchNw3673odSiLuq8bm7mNKevxsD3mBRIZIMI2wNDCbB5koB7jk3
ZrfLuRQKEnEimF9IKMmAUSLXLo4k1qnqWc+d9Kzft987vrOLuQbAeM7ZedFXrxm6SRNcqLwVKhi7
UKbywpwAVUSZZYhRDHR8ojm3cF3pTXq414LJCw8+Q59kf/e9UvL5ci6tQKHfiFBPEQftmcHj03O7
FamwfWOffa9gEh3PEadyp83dpScOY6s0sIMQpcntC8PulKQxcAiWVYt8eKW6yX/XS7kgi9MOzhUn
XaJ6lpLxHbUo2VVqKuyhyBmxApl9ypv4imVhgdWF484H42sZ1uBt51aQRSteOtpRE42BO3/MIybH
/uslzoNPNfISRV2zx8BAe+tNB3sq7uT4rpbMaXz5zSSWSJzahAluLq/LmYvwoCcsUmkh6GJ9/Faj
JYoM+wCR00i5KsGwjfIKs17nftBrhPfPNvkXzcV6Hygj1VPVBHMJG881s/CFfa10ne31AxBThw2W
6SyzGVfnOPX5UBYdTjB7btpLq0Owgz08p+qd/ToPPEsct85T17aQs8OEonmk9B2qq6s22xLr+yM0
2dNuDV1C9RBZ/7i3VTXquUOHcq3/ullbnwHmgOQaBMQIikvycDNf1+slvcqfvPO1W6Z+As8PfHkD
7Z4kmxFqHnJa0tIlmvwWjLVRcvoIcCd6Uahd5V4WZlQ15tA8551oOTeLc8HUC0Hxux0/I5uPOcfM
WZd38NWo26uBZu0fgId1/eOy8EY5VG81+ttXtpUzEXQMFcj8MigBkJ5qoRxPQNqcnv73Yd4hhDM3
N1ElUZmBCsGoRiqSYP0pIGFSf7CdAwpEWduqWsezIaLwwVNWYkG6BHCvYOUT16ZEdzSKj+qY+jYI
4wDy0YDSv/0p6jRkjAyD5nhmR49bg+RitAu5/AL8tKIHtheyg1V1C2ALmblawsISQKnnhm5/C6Np
5ZGTBgNKhHE+MmInkd3DHA/I1vyhl5oY9cOFLOChBZ9/a9rCbqng3xUp17RypOmHBalovYL91AXJ
SBdmilM5dtMvEteeZ4Qe3Q9jOXsJW9/vKW/qwQO1dZsfeirnDQJ+dCiFT5YWBfLSB0tYl5AUmtUG
/MFTWNZ4whwKy5sf10yNcoGulkXZBWdFD1UZoS+CBcApLCIBEbE2k8OPiegTk8YqBsy5QShKz07X
QOTEKIJj0L8FyhTrGZITvTIgcYq/im5KVKouMHNvF+j+H4p2TY4IdaybDQDYYdYcXIHz8TrcDDCV
gJR9PCcEGL/Q3949xREaFegUodZlmD+l6Bcl6pNrax/Fe8NDjGZcnGP21HtNDEd4VyC0QNUyCwoB
3HPKfTer9RT2HQRxAp/iEzqVgDAmFKUQA5eMR6lZF/rJS8+jQDDh8605MDFt8QVWI408dogvy5PH
Z6gc4Da8dUkPSl7T0ZMd1qt8Y6z9XxiCgtNvlZrgcmMgAb1re6t1EJ7VEr5acAH7O9NeHERUT69o
AZ8A0P7lYX0nT5Q8xAIBtNDgs7+Z3/Nr0UsapBx+gnA7aN+F9gaKqplXcS9y0KL5a2VFe3P2K4Az
f9f48RPep0lcET1YwT6Q3WFzd0pl/0OSKLCH+v0GrmW/43nZ1E9zITNMcCk6T2FZzTFX8v2mtekr
KTfYkePjyQNyFD4vt9AXwm6dpyOqfe6+GTwz+cLm20QyroOEIAE+lYo/n+0T4bT4zukBNuLAxPSk
BI5KKrYq0gkVOOkNQPZ0b0Dyw/7PB8TaCJos3nvy/YxiDgx/VRcModNt32Jh2IqsDGfb6QfIvdIq
cuFwQW94E5QG2575no3pgjMs0OaMRcNhoKgU4oA8jpb0OAI3N3acTS3dAygxTXUhg0FtMIGBP/Vw
IrcONaj4e1EpZC8ltaMfvgruXlupCJfgM7kHqnD4HvEpN4bJeZ/hk20tISgYKLOeZLEpJkn0ZzSk
18apPaVIgjEe9GtLbFzsDcWG8jZsrjQHBundVHz+4Int2dDrSk1tPZOfey6H2f3iro+GUPoi9RAp
7lI1/IeZW0Fle4k+xOtadV3iKZmlCYRLVMxkQjKMLiwpZd/TfKDlU0TlS0P+kkh24X6a0gcPMWSP
UV94MXJYob2rQeLgZNAbEqTefxmmA/VmDI73/yJMOpkHuBeQBa2yg9n/vw+zNEJrs873aJI3DoQk
Aizd41b7Mcv19fUXUbon4hZJZD347B3ee4PPVlMxVm74yKL4BRrdayCZezJ842+LiNH9IGpmR0y6
9OsXdpP7BOLzkFKdo2kx0XZaGsV0LfDl0HZZq+K0BShm7L4nbP6OVADTncASjeUaUMfdDOLF4yQG
F8avjQNvTK/mB+4/6tcAielwPxCxfxxhsXEW7CExiIZKD4crMk1VE0EEh/Dty6WNr+h4uH+SDlrv
TTk64TZd+rb+7UKmgTKSv3+TKFUqCz2TO2/yJNaLi0raecDH4hQayNvqOTZd3Wa1mykVL690RIlB
usr9/YbpYGfdPY29GPpD30iIHliXaalN7ALd8/Qz5SgC6sAcvBUYFmIB0QkucOfb1fNqjbSffAGf
J1/nmRTdk+2zmp3CkBCQoPAFsk5+5qx5NsJfaK+TjTWSme17yjXKyunkiPxeS0TEwRS99PURoKoL
IGa7WcyJJM2lDC5ofoEBLW46NT3xzl3vYHc5Im0p3XkJwU2DAbBMKxGBSoWXfWf/KXd+dOoS2URM
vKA8GZ8KJibNmy5qXUmQCXKcZJns5/RqV8skHvng6alhNhBAN+VSWACosBsxmXlLsGXfDJBxDHJU
02OWPnGA7DysicwiWxR9IFpn8JjS02psKX+lG5QT+IgMwBED3gb0Ut8qVWdWOZHFOI1wOaE/Kq23
sin8Az1cM3ATkix0u+VglDO2WnsChuNcN4rZ4FVEOpY4gQNSbJbLHq91zIwk82Ffbiz5mLAmXQqv
1ZP53eqZ21NGhWeau9viRfX4biCN8Rvkxkahv/vBiI8rhqfdzUvvDkv4ou66CZsW6omqwqRuAd0z
s8odvCsfFFDnBxW9oJHbqhPBmGqsnYKKk976IPLluLWI7RyyHRS5XeXUpVPlPVVziru/uqRRoYgD
1ZxEyTXQmH6l+pQ8nc1Azer2UmtVA3hVuYgR7HdEgesl4mBRn/TYwBVK7EwoB64XfSgKOUrHCQHe
jgxyOe24aQna2YpP4um06v4sHFsvMPon/SDGrQpaLPR5mhekOvHsmsrN0DNt6CP2kciuf1TU5kap
lP0MeB7UTJvgnUvULvL1OHo5XvZqhVkswMH8BHUjbLqC9Oi1tsdm+QiotNDyE+0KJIk3ErNQhCvv
7n/ETVeI8gks4ZVxTa1HNgKFEjRZDkzJslMiIBHYA8xG9sJNaFt7wVOxn5VWUZb9sF8x80K7s8ms
bkzrPoeo8Eq2qfAiYHHOg5Np48lBwkXxMBu2rSB4gHxCG6sk0R51hMtVH6xF/HIR00bXSxGqtNH7
h6eF7vOzQ3PeijnnakhFxIA26kYfI5OEOuMofbWEJuw4rS2dt8ppxBMajb8ahUTTRyKph5CxVr89
dVaLJCkNdKUB2Z4Nrv98i/vnIKku/x/SrONGaNsMtZ2obiSV2HNQZa4bHZu7xG5LRoscth1bpyJC
TWeeCV0+F1RidHRCwdb2EvrYNfQN+tBbmvMACBnchTJYY1q63EsKzk+Nfij3sgutigh+1DrSN13n
GCGCVKcn6GOCcCYJbYeivdQPfWXeQjvANChxAXRUkKbawO94hT059akcp83Q+FTHMyFrro71LQYb
mVJBpJhmLbbL4Z0YlZgCLInT7MSPePzfp1EPzOtW5Ad4yLloTC0TMAv2nCiNr2UaRcQAK9kJ/oUL
8b2JPjbk0xRsZe8s75vnM4xVjGXNC1BMEngY6EW4A+/S3rtf+GpdaFOHC8XhF96jSDBFRPgS7e6r
8sGwdhdoiKx+iZ33kXW567T2fGxZ//prLyhfPlPMqnj2dqfvqbmGprcaJcnonpGOK+ldq1/D5GwL
5+9LrjwqArfnyWrkR3to4akxv4pSMFJ+uZjKBc/aop9dvMxhKBDFDoUtK74wvD8mgO7pDAv4RzwG
ktf57hRrRv4IYi1kfrNA1sjE8gP8KJKccjq6G0KfboxZg1uxwSVkSD1UtFSynLDvamwk/R+G4B9K
epgc21WjF0hzKTlJDEMl1glLX44l9tciMEKDtsTCXJFLLesA4Q15tADMVqI+qAEBYXzpfTlT67nR
LPUDFHO5Hz4TvZ9j0j80rq30YO8jA8QOS9QJJyJB6ccO1jm2ABFUiJu3wz2xkrn+8cw4dJqJZpNv
wJlzygTBGWjIHItYdtuKrIzQjlC9waO8JXp+0ZV075fmOaBb0/XnT5a7fbg7tyIczEaPjH0RTmKl
EISHLinqLIeu80MecCu8+ZNk4Dm6ZGUIf3qRSdvzd+aYkJpo9O4AhMrvYPbP/1s+rcJdAiO4R89v
2T6Eb0aVLBFZiP1DwMW1h6sudj+b6CKhNB5ETRZWXjiDRu+OTmOECmMDvdALiMQeGxUmGXwm2Mkd
KfsNJLJkZQY2F/+fqoRQLEfDFtCPusNJNHFfcW7efHwXWVA9O9YrIEHNGkwEbVEmeAaeZrN46t5Z
HD+KZk9nrgDma4pO8ch1gyKUh6BE5ucqFgoYAZehTH2Y+raaPstcnM1F+NsU4EepOWA5wXELj7mx
WMjn9GVgC4M2vhXl7XxTGH3Fi+VNB2EXRWbtn9/vNtA4oVPpyulVqEEpWvOmJlMGWHbq4liKCNFI
5ToMmzU2s6sFe/vEKRhHlOrUdiLbn0yOsHKcPPdR+EX0Xqr9D3wZib4QfUaAbEPMhYUAoB3N7yyo
liwhefdh2SII0cBnawhoPv7bSl2GFQMglUkObPeCifAYLIoO3mW1wDdAVAGWMyAhuTuSCCtOSa8x
c6vBrDDl3P2gM/KZKpG9kkFvpecrfd7lW0QuWYRtF/Cb7B6zb8XMp0jFdSrsRdghfhNRiqaUWxJK
B9kkNJ4JYUYeUz0HMy7pmJk2SxrGzapiqwceqlFD8QZ0bntwqLnqofCpSucDGS5z+xCG5cEBnExw
6SgFUP3jHQ4dDQHy2OWzVEdzHherhNi6YQ++kAt7+HAOq3wuUPu/HpHpx1xTiGST2Ki03me5OyAr
TaNR+1OD42a0x9miiWH2N/r5RR8dB4x8JevalKv6mFNNT0jrvRzUhjfIYZvwMBeFQc16gE8fG3qe
UnjZvfw3akbSDryJt8VWpVHGQP1RooyZOLMWHlrwWzlH5TSENFAb1gPGYFqFMkXy7bX+Oc8jSTMw
xwtD+8VxV4JVrlfyhbEA7k9ntdz7J4mRCh04JqxiXhSwks0iFPkUAw+crva/miqcwiiVnqSE6Rie
yha1ZXLtNjSy5/6dVDmohNZDCFM3ubv0O3aITD1WP1yjcRUq6bL7t2VtKiEsU/cM5f2cHvMp9IWI
FeWEnpA/19oaEJBWBjmd4kGbp+y2+yx+ZHYT/stEJz5LLIyWF3wdbc3Xl92NZ3+WopkoYhxrpSSF
txvS1tq2330A/0+ykVFJwCbPUMJfMLNU4Df5SC11dVIew0HVjK0Cb64gm1JZRWtqkKLzJD+YHFl+
bEO247EEpYr3ARF3raKItIJGoo/KcgeSBR3vZnXQOobDTbTkIlYLAu4iMApxdd1O5v/cgQnsYjNf
qTwYTCg+3HF5LMi0y05dMG+s7QdNTzEqqe8JSRozJDco36DE5WnvDhrD70FdN0T0hZxEmLmTOYxn
/R9eSAX1rX3I6BH5YMgRlmxk0/xdZkCgvkH5r7BTw42ZD0DeOam2ch1p9ZoBUcCEGAp6qaSvNyWp
0lYCjpTjDaL0G/V7W52oRKl27kUJemdF0luvlaUsoiXIWtOfPgCuevWJvUjip0Ts8zAM42aJfWKV
W/PlNwQZuam6GoE1LTNwNPrax4BAhJNx+0qiEWWEfoO/P8XMUwW3XkryCdV+3e23bjGdSS1GHjqz
xbFMRWbncrRByzebu7JKzdmenm0CUcPTjsYAQrbi67yEMdJQ54P+RwBpIIEzGVnJvaXgVSzeUseN
a0bUk1N0P/EkeQDu0deco7L0XlaHwDl+qllQwYQidx1z0oEWJC6ktRN/aSYfgQYxYdnDdkPxTQrV
0WBTxn7Lhbm7iBge1vbs1uh6amjZkH1DyVf6L7W3AaNoquoDvfBD29OB5oNG2gca0DB1EwNuHGz6
0w4jXrm8NTK1Jk7kG5arv2VS82GN02tlNhbbHwxDmLWRa1Hl0wqujiJVZP1X1arDo89aY8m2M3AH
xZT2qaRSnRM2KUKzF4hN1mgKOfpzFy4CCVmhHBec1nNkkaU2h0P35qkl32j9MoAw9Iipbgd9XeSi
NjiQMnTQG7l4ga9lEDU8jz4XPk9hm5HV+WtG/6AfPtZRMwh/iIRwtBL6Bs9xmgAV76h+WWbNaclW
mouZHrHLMHIDexUzHrGRqU1pSnGIwJf0ApyogF2V5UVzuSJkOlduCzKg9NtFqrp3lJ4VfZgxfJqu
qwv7O0T1FTNJCqjdq1wG5rZWn6xEWMJjIeqsH9R5LPutRRREy1dFwvFu2ZRPbUEGJ5kujztrgYU7
TAPYNR6eXl8rF6OMkc73FMgBp+7ZXEnSrdO2NMkcOURT1+ZfJ01XR8x/ZSh5gHWHHslMCHC7oYL4
b00RuoKJUiOrZyTa1GIB9Gx387G3miCgDuJHEM43WzbtULq13DoZYiGlIod08PR7ZuSkbkQXiKOm
QmcqX5NoMP7Peh9C/fGdv+Oan/dhcDThvLrOutUbAAe6TKjJwnTp7zQsbwv93vk1++EQ4+2jLB+K
D+K62+VKNM8uvvUSFmLXcI1LlDFaZ6r17pvFTsvDBU+tVM4D6ERv2KPWdNcJgXMYkjvea0SL8MgA
idGumkPDIxiOhsBDNDCesnGIezFKMDX2GvpwmU0EoK5FVmcgWwM+D0QdIvpws0HO+DoElAX4IZCc
PHdwxqPHi2ou9MYk6uOQxAfLe1nkE2fmZgrBCz1L66YqCahPFZlHdYuHpNfpxyUPjAhgoJk4nkaM
TPn6Oy2d5dFW6N7LeR+tEqyyJqfOITRQQ54HqBA/xWA+ozPlYx4txHUxShy/afftGQH0XQBQsWlP
VKMm+K8mhCur1ITF0j/8ndCB541OZP7G8Uyr3+tg0+8/SnLLUsO5LxnI/4R1GSPg9Ghhf31/bYcK
a8tAn++5SrEMBanUYjf+9nRG/2r5+DcaiECER9WUOEWy0atVktZOMYdIDUqEtxf42hArzTHakVUR
jFwL/CtwW3lkatuPRQ4ADO2/Z7Kg0w/KhTBfewfssCiqytBDD7uaJfmGj7qgvbB9coA+cXMUaHHP
A4X+PjV2ElcfwTFNF0Y/u9d+TCgVqGIpuhqQhYCombBenHdcd8t7x9O6c2qRkfrqyx3iBU+bhvFN
iAEsii4/4KeLoIdJFhFPigLC2LAGqIPsCRTVETyCHR0NFdIYnuqoYfOxObcjvySEHzWxYSdWvydN
l4XfG0XmydjOMT7Ymom3H8gVJ6jGkKKuCTZrN2JtMSdNaWyMJbWRkOQRUnFxA13x4XCsM56ateYZ
TqCYV8zXcsUfFEUL1Z0i0/jYABi4n4bXcBrhroyFP8SaYROdv6dcTS20h+ebuv9zaLQza8CG4TdL
BlFewZdORKNVQLssPLq/5UG6nysT793ez/94JUNBOMtQIe47Hwkt0YxRjVACsPPul/VDG79xODvz
kRvHKLTo9LVMG0oxYd16MsW1FNLeKIX9gbs7KosIEUmDDJdHJKyvAT7H5xhkQq7kxi8UVUuV0xGi
nhfd++j4hbQN0BJGKqZ1w99KVK8sYwilkZ1gaYHs1kw5JNYrDCVQt0ofYLWXvS7WcV/DQjbkKkz1
qC2xRPWF3ybLJDFjHYmWdmrlNKuBVN6LfyexGZ17aCLvbGegiZOVUoIs0t86lk9Mrp+pRyFYE6V8
WA11XLAyFc9+WG5rjov82YW315loyZ2CQ6ReQp+qqlWaXQcraezsbwbr+cBlOswTaFZx/7NvLojH
5RccIbkQMN+twW2ijG4JiEIXbIdDJCZKJk4Nhb+3eT7Wq7/Fpik+TqMYEie1owkmjJ/ZUXJY5Ymn
97BS7R8PCG7X8i9QqEklQP09hx0BPjmJ0WeFS9F6v3iI3bYnjMKzC31sEHoJ/kxqOo1bF5F22yS2
dJJ1l+Ke7BcVRECqHbhkcBiA6TAP7pUfvR4+x+pQNDU172QKKw04wsqrwCGuCr0vYdFsJj9FFY7u
mx8fedVXgGY4HqNsnxEHWyDS3Ke/wzlEbMOlgigOLjIV8ccwEp3I0ltvMs5a2V8RwOIgb/V76+rC
2J6r1hyPwqwA1kjj9LEnGIn1ZqXC+PBFffb+qaMpOqnQiyE41v/A1YbeniiP5aLYzigmPUQKGc42
CKNwcj/9zqWuvZuPNVWQDdM2UeD6M47bi1TWIi2XspmvykRzg3B3iXhM+TG607J1bWwxuYs8i/3W
TlA/Od4aN8gO2rHxeuF80ZVzUmwAb26dsAZYx9YeD3sJSafUF56y9bRMzgBvmNXWtSpAmEbXAtLu
DhAiyhxh0Vm3o8297VaOnw8f3qCQJ33gn1ckuGxp0EhkgjiAIU+Smsmv7+Mys46I8vvGlnuBfeXC
trhKyAnt2K+UgLMvFnEOyg5QzDPDFPwPwynURe42jxZwD1b9c3pDUIz+1PocMTFBejZbR+rbp/7C
t5UaPeR7QJ2QvwcUdGHhaE9gCrrvzKqnW0k/hEhyMAA+VPsF+OTpLyc78tXGB0iZTV4XwwweeLde
G/p1kO0De8p9Hcho4uIE8hxsKNy7wiHv8ls5M/3WMU8YXmhWUd1skbbi1Xy3HMf8ZC2nhIds21ry
Wd4gs2fsdevAyJUzC/YKcyxevZ5s7YNGXkTYZOtNYnq5daD6V7T9cyZseE8p/Yq0OOOQIm9hkpa2
byCO8iOCKfZB3NXh+ayFrbO9Zf6xC4KICXhguTbprljbYz2kQnw6iGmpU3JGjDuMFAUu/Db4/GoU
tqDaMDLpP/LX3M6FGmyZ1/WUXdDE4/Ya2AJfrHOAiwTUe2oTWopTmsvysmfJwsLfShoTOV8nFr3l
NCnJdW4ESVvBarQt2JzQQQl5sEgi6FlPKtZV+MqKFzvkMNOLfJxXXGyqRrXnIJ/kCsDfZWzj31nc
FGZSxB6cEt0CFOvBw6S1hfYMIItNFTO3v+Ru4KWlJwDTZi9FuovH8mBxEQzDr8/umeuTxuMK1B1g
IVrIZ55Dg/jPeqOk+fl4SaW/4aAteeIufuH9m3uLib44HBm7xoE+83m9y8bKnw3Tj6HkRuT1h3Tn
QULankZJGwUAYwAy36e7Tk2Mb9o+KbMxhxlhTLqcPejkYfbp6u74ir28CZYGFD0SvmtpclW/6DsK
wL2zZ4myQEMnVV8E400ReYd3MWvAkfiyBOkf0091kQnDqc71Wf2PNd4qlwx1pMBgA8JqttENB0XD
ewok+Wi1XJ6k9V6+n3vyqIavRz3er7ksERCs1VWmLN0h+v9PjpckjiVydzs0qOJhJtdilmHO7iUE
mvhqOk46jFCz67SMevbb69u3/cEfTj+21MPBnO3Ea+sjFQK/eTiJvggXuFV/8Fr9cA2YZWX4RSWL
7r67BRqIU3QE8/lUFZjMK1/m0NvGKQY/w1FwZC/PPksEPC7icyF2mWriNC/tOSTFZhPZc0SeXKtb
TjokxnIA6ale7gncUSOGCLfooHb4NsXLXvVyaywsW7gSnaslb1CWR21xGyCV5Y7aFDare1pR/khT
+SCxe4DSKJWcsNs4OqY99n7n7lQbxafR6mGMgT7PDaoYwUEZTHrA2xHUvbgNCWz2UdiWJmMxJM6+
mSjOoyogzWCWLsEUq9N1mgj6DC+R+gTU6fIGBf+vLFwAZ6hdZyNbDn3A6uqYgdYido5HnCTZ4NW+
cLYBEDfyC+aGnxnACNrjleZiT2aktWltHkHK1oqxs88njI3RyP1fGl/3svCGjmTfwwVfFJzGTGct
vWbHhGbWOodUJG/4bonNzlJci7z6eVUoeBGah1GzJGFCsydOqI+kBHipUEA3wVtFFbjsOqTL/wE7
gBpIUHjzBOiJomo1HOwIzvZfu0E+x95qCnnpk5cFlETCzE6vZr++dRipw97A9JTdo56B4z9Zft5T
k4+PgJmJN6U1TlMAFIGYRjAvpWMOyqYA4AntCfqZY7WY2aOjqiRX8C2MrpDAZoB7EJ7a9MMPL2SQ
XTPlnEMI80JNWLEr/W+4D8rRhgNeV2ju3NnrQqJCqplT45/kYh5rl+MnzN4VxmEr3hYA5S/x9WV8
8y5szOw+dwLceB02+AF4UiB8WhRwU/UPISQUATSgI6/5DmD8tWfZjUMva03zWFiu+WTgEbcQ74Yc
jdlSeyhB5iCtfgE34VPLyY8YQYG5KhHyn35jLQVGoLOkO9nW9V5ASP3V6WVtMLThKZ7AbaMICKv+
EQHEuiU9PyXGrm/dfvaT98JCi3as/BJNZFD9U1ch51ST/p2L8isrLnJohgCaEfQz+6RGbikEf93v
nWhKzFuJELPjuAHJKAohUa5Af8uL+QmlWD7rCyu/ojqESzMkoCtL5Ka/XV5JVMOxsrN7/+S0ApsY
sBQong6Aev8gdahPYTAQF8WNimKMcruN2wnHQcEgUrVHRZzC5yM5fbtPWDNo1d8GWoPyNqnbL6m9
PpNxy+q8lelnWGYCvN+rs3tXYvulLAMeVXcNKDkcjW1UcS7xua7i78VqIDscxx9q0UMPy0YW/aDo
I5ym7i4VMYTXeBGUlgZBEatwjVH2rzYB0YhY0imJ5zPYrYDpkz//F5zLru471m15OWpIkw7iF/vv
g/mte2XkuhdZsKqvET9b+jxnKGlUfv63bMX8/3dm8yClTvO7QieWuubY/78wXciEoQ8d6AHyj1jx
ZiKoxsrOmqjl7sGzyeTHylakHIS3o7M8ddd2fJ+bHqVYK18RlzqBiU7B5xQQ9P8MOMYqLqvC6ZXl
qWJY49jUYyCfvCka+QpuIRQzXZ3RTnTxhC19/f/15gpxmJstOrAay+72+9e1x3EeLU2BvDVNxadY
QknJAGkCG1EyD8JCmfINxX9BnDo7RHs5Pf3hqh2rV6X8cAYIFvk3BpNHjjzo77I6kPp8nXvo0pQs
Hvhku4cb4/vX406drO5Pp2uHfiOmdv8k7DQ2EAlW9UehtH/A+Pz2Oh3CxpEwp68hn4TnZHhJueoy
xQ6EBA3I+hu1ZoSF/kcViuyRztCercXMea6CunTDQMcd2lYkqlknMuMcsnvWmN/Z/jlYbX29NcuG
OEadWJrS0hmsZYSWUICzJxpTzL+tmhgUNqRRF9Dp55znog2NoTZWXSQmmp3Auw45y0yhwdXqyJSU
jZuzoz7DGhxlaSVqiSUFRUHENQCwZJq4tnuTb1vm1KfKWjsfALc010lv5y9XKqBpX2AlgQXb9uST
Gzowv7xyS8oxvzP0Y8JtaxSJKgSU+eyJztjeg9WSLdrzZsu+/iZQ9oixPtmY8vYZqTPznodIdf22
hn1g1wQOWOmbozde/Qhsxn6tv2uzm/ZBlI4aXvMOBzrv8wEa3ZivG1ZuCsbbd7LncawxAUTSvgfa
GHIt8c7wkGDjA5sOhEdqyN58ExB6VwxPLsxgHTzP7NZropv4BrtmDfJ4nC7QMwr1jHEuf6dabK80
S+KuH0m+lwxIY5pAsLZrmuf3pFxnBuvU3CxvwHuBamkhVpCQy82OlP0cCHQMTQMj4FlzwL17V2CT
Ma9PkZlbPgQVGZI/8aRyPBuO4x/OcngPnmLWeOxEii4lKvDWunz1uPRSU/gxE666Iu1VlymJc87l
NnZVhNz5D3DbJXnh2IcXVls8SxzMQqYt3J/tIjWW6LHNJzeYXiQhqjwfsND9+JT8BQlXAPkiXfo3
VL0ZhXjV4D5VcbS4SGzSFjuNZ6Xd6tv2ETAK4uTeDZkg2rB92fLNh965ku+wlaaK8EVwIzGx1FTX
LELnnQKw5kAASAfHGaTM9mkqBpTH4WevxM0T1OdCHHGXzB9+3pomer95r1vdESTw2dFzYClrnNpW
2OgVGCqaQde1dKqByKX767Cw4tL3U947Y+Ifr8pkVRfZp67v3TYwXBkZdmaViwFGSmUkpDp2crRP
OiKW0asZFiQiSkhoynD7umiXChOzPShVLOKvtiw5myzRBFOqZg9C49wSna11Y1JLbBbhXvYaxSCC
hjgLp239/PS0TQbsczfKa07IHPeQLt7GLpKoRaqnWtg3z90lt1JeeU1RLoMVoD8UDu54hcUP7B7M
HDoPni/54GThH0Q3G+0gXreCW9UyFnEz/h7EPzIBC/+um+u42aYc7dqybsq46sc9qjfoVuAP/e/a
WDP2Mn5vUjJlDm0FbXjsOfGPpDqp7xiPjkcxtI5EcuDdSmyWl77pCxRkIafdKiT3fTcKwYSSFyzW
pFq6c8UFnf1uS6EqSeoOUKBXBCCtEwengQ/2YUMUpmarwYsqHbohjdTqIR7cECj05oBAF3XjgNs1
U//sXatlzpdH3Emd/9vnMthLYwbWInWeow7AcrPANMxjMBrtZkPhZkb8PZIlmmy8/R5quLTEFOR6
LU0pDp+K4snabsICrmZg5h/OQMJyzNFoLEMd5+XOf3HgPOJtLgtoDQXLC4JaNdKM+eYqxmsQp2ED
/SyI16IHWV5x3e99bkgu7Y9S0fYyu/b4miB158lnMbpD/GBOiEFH/cUY/xwjjrBi9jp5z4oTYN7n
ySuE9LNAByFtXVmS8SEUUUR+DWJI9r6d/vGDb4rzP+F2MKAVy+VQ+u+TfUM0eLfYhBi+fYspT9O7
Xr1ZkfR7Swq/XxYYsyDo9PrH+jcuFUDMs6Kasj+oPjNrSGeNpWxFwxW8AUf6szda81zNOQP/iTRR
Sh+jDnIn15f3HLFZAJ3Uxy1qApylNMWaLTP/XjtzKDj90A/ypqkDZZKMtL8Fwjw31JKCuO3gMdvM
W0vH2g5JSe7acOrMoD7MFIanoD4A3g9sP1LJfKXkbIkyMz7IeJK5+vFFDsKPdupRkidLgIZ8wavt
3QYpyqZpxSAie0WhohZnuyAAqNsZ9gSKmIigE7ahtFs83eYHA1HpQXou3CR5YVZEKZJtvk3QqB0T
MNjHJ2LG/bB+mNGwm/IHGav9tkXXvRXyR/NlVQBJsqQc7C/iu/riU1upA1vaT/GBRopkXAoltwfh
PzmfExYxtOHpILYyHzmNfNRPn2BSTg37bsUy3FNldm2Y8DwCQVYaegJ/YfR62QQJABZ0VeDjWJ8i
vIXEErGlk5/jxvAlygVy11jbMQqFuUVq2za4yFcJMgUqBbuWSyfagZ9LSr5jNj6s0i8RMZ/2mw10
HlWbnByxBjFyOUPhtw8orid5M+j51DJq5NnIQQZIbQHIGEHyQSfsvaaraFWqmM9XyLCS6JqiGSf7
1N1y7vy8MxO27ZMNhdJdqyglUJzejnuAU3N+hNpXogg1RdWKqlDojvXrfM/+PfG0g7zyLOTJRZPx
xHxtFXLi4NCCDdpcjeo2dCrIaCCpdnHP0micah50KdcI9NRP0iL4BVi5tTiTCH5SjcuGGNnZPGOz
0qQ56HWotxkM11rkTWhmI2aaKJhlJQCEf9+SNUJBZi/Xohw52JIJE43ZAnjDbJp7zCEtWFt7NQY/
w7La3y6dKdnXF5MXfL/Hvb9AX+5QYhRW+Xi6kOYQkv3vSDFXRMIAGKokba89ptrHLf/rO82UvnV9
kTnsD608OlTjbcljl5p87GwWvElgbSfOayavXQJlpfhFOisn6ki+RzT6K/tF6Ekc2C7KX415bMjp
VXpa+DRYG9iZpPLABQhUt/dATZWPcgw+RKCpfM2l/OWClyrHaC/O9LrvbKfg+x3T3o/+DUvBJa5W
5n283L2tAw+xwKDK/7PzzJO7qvkkCWz/u6nWr2jQrhO8dv8XNgtuEvIeF8bj9FovZEJb6vGGU6jF
+zFuSVlIueGC5G5aSpIIVxptqY3mrRgPancZ4UqX9jgkjZWzOYV2df+N+6GowlDlB5HXuPYCjp1+
6IwK0Fkd9bc3ZlfTzTxqkeoPozmJxq1uHolmnWwLY+6ELJ3cDg8nOInJ8VZJMaFnXvvjLbmj182p
7dagg4i3L8t3k+VGSizIjKX6QboB6mbmYjfeS4FqDLkJ9oeWvD85ehmvdBFmVzvBHh07cVaxIlsb
BJUV4BCePZjiLQp1NGzoXxe8DGaSRejoLz3XuJHOkQec8pkHT5es1WNOA1Be4fYUJmzlUo36LqwV
opDltGaGtHOvSy9CYf7e5h2kBqzy2r2Llb4F92SAlnOhwm4xNrXxrboo6of3J4HK1Mr8G4FF6GrI
T4JOTcHtx49+h74ZDf8ElDJ8GHuMr3tiYY0o0HySfZ/y+DrO5A5igYEpOZC6X/ivhhcaAKak9ECJ
5W9u67+cXT1HWWvjqI5yetDeCuY+nXcjJIwsUgomOWwEG+hLmTdVOAQXY4gzrdjWbZx5+C97Laes
8ArQ+OMxmhBWLZ/mBHJ2qpjK0U8GH52zV/OYBqirDiJqclwv88Xt6YkRMVcbehS3Dy+ph3WAk9j6
PPSbKe2HvLQXxodofeh1SpUQuwt4Q8oQhg0n6L7wLQ8Zhyoou5HsnTBOYDntIM34heXxFecjyHvw
MV3R1BpbNrUM2jY0o02C/dYMJ3aKiYsfspl9QMYnQXXmQSa8juS9jiiFggG3/m23PI8jaoHJusG/
vB1jwg4vLav2lmOs0EvCV7fO55BnHuYBsicisN4f8k71ZcW9LJkce8KFI5p/9hux7hbVtTd/CDp6
R9kEsYxNUENowpo6+TVd2OpiqmivybawTBVYip9vKqRg4iSEHlNqmmOZvZzEQSk37Aq08CW/Eabt
hVvAvpFHkUMiCpMPX3WaElop86KXlsgVuGRH9sFo6bEHqRnSaqS6J/LahZ8eN1+P+PRS5uuoJdzW
DibRB/bMEJDx6JtzFuRQgX/1GPXFqvMldDEmyEkxYFmfltI1Joau1KhxhEKum1hiivoaBjuzAwEC
hbUl7SUI5xb9mYGor29gQxHDaSxpfJB4RHkQdyTXZKwu53AO0BZHxb3CQZkuug0NWU0c/rl4r7vf
Km3I4sVFEq7de5GaRLNT00qqYXoIdzFVzZ0IFbxWnTyMdG7EOk/fEF8NgR9zCU9GV1/d6yBOvmGf
dlGpUKiQWrJt69QL/k6xPR0zDmviznxxFNZZc7PgJrk9UqfvugYXgmwSsZMmuFgXEoVHqxqp5bf9
NS31eZWSTgHG6OZqhwEcQXWbgwCntzq6CnnEe76VzeznwRZAdtb9qJGlQcuFbSHzTd57hXj09orx
b5cZmtQBqzColxSXkSVdkgMKGITgyaXoSJZBxmwAleD9AXKbAR9VpwOIrXI/doxJyDc6JBbcG1Hi
Z4L6S9nf/I+Xa4p2abYmyPguBZ0yS8QoRis9s/U2D5S5GCTUpQ1NdisW2wZScu8qb/PrlvWYuNJI
ak89fjVeBT+v/3hXTjiy+Amo/fwYZD/kkfP4cpLYicJEia1sV5BKQ9Tg2dffH55djh3MF1zJ49ya
DgpoFaFueo5eAZNn+fsTbMMdH/8Cksk1vKxCsmrWzTlMkriCP4mO3FnsoTko+lbYuR03GpTS52dD
5MzjeVj+fV+iEH8ntUlzPVCHOZsEM2NIqeblMc8+p/M2OccKiM/3aVU4klFWf0ZdWBrZkejaFkUJ
/a/1Ql60FMnaggUTwwvfnqD4VO8l4D1E/c0KK4Ofh/A1cYHRpy39c8ZWnzqev2OOTqB2AKd6CbLV
14L1Kx9fsyCj5Pk4kV7BZIvO/v+2peobaW/4MtLi1coTRMP++TcSlTEo0TjWkFJfFz8JUk4QjqOy
hceBFAjO1mgHluA4On6Fx1NlTz1uJpZ/q9B2PBNZpCE4mcslwDEkN1Z3PV9mjZsN9XKDJDypT0Qa
HiwVsV0RSFQCD81nAh/LTHae03mJ1qg4RBOgrew9yRd1608dr89WwvcNiA2Z4osbUdg/6p4n7Gd+
3aPIn5bvFcFcvAl2fbHMRnNi9ZaqYXk2omM5dEdCBzP1SeSPga0U3VyQDoZqwVmNbkHydubNDD1l
FKj6E0ffClmx53zj/gA4QP7vna+6XQu4Tpvl4lVMbcofgumYHIe4ELANrE9XzTHCjTgf/d/2J89E
BZv65b4mmu5eXWlnbG1UyCHELQswVEhLEx7QwpsWGFjYaRXHZssEOqe+3WOVGGQmqU9i+VEgzm3G
sIn7QWxph1DmZ2aVZH+Vz7HvXJ9USbckgYhy01htXu7MucKeWC2J2QWXYbVtcqOEah43yD7hYN2G
vTVDReIG6dgfY/5q6+8GZqBISUyFIAUjFm5eN7mlUfs59XTztMZbJ8SQ8iTEGj47ysjHbyJRdNJF
nOVQbtw4W0K+l5+O8gI475kUlyaDzZ/OQKFKgZH5RasNlUqMFXo+AaDGsaImDirSLMhALhRjt/UD
r7QQZQKfdn7x/oGl0pRksqVUUWDoWUiN2TQQA9N3Yz9MHlB0N2l51nZtpciq5ifllJf1OXOZYs6T
SNQlyW+H/WED8pZn5uN6lKlZVRfSpJu61uKqtCabI3KUhBRhx3sTjQ+LhlOxfzIFd0RODWyGdmHl
rNo6W09+1lv1Wsr1kMAnfD+cXtyVr/RfBVDiSoKsmFqBqvb3K24A1V7+nAIVJY4nA8Zx7rww7XRO
Xs1YSoPvX9HRHlwQd7jutCG2FNeIUr0kp1TiuOYGmQgPruDDZLJO7wDA0nZbmOYxEIiaLb/Z2fiO
0RT1Wrgm8jY6/E+3umZeVnLugPtnpoSnWm10yp6GO/1KIWJU7LuR1YHtbaqg1jGl0iWJNlXbCNua
pZSMrksIzu7pPPhiGFzPnFPFUVK6OoOiKzmPa0JasM30W+hbfhxij8LVJjApIcw9IuaVkiJPC4TK
sxOs5YWdvGU3KMlHxPfNEL8I75mJ/nmdn1PZcCdTQiUMQ5qLgP0+bAzo6fRjglUFua//EgEtOrYv
EwRjWJQUCSquSJ8UHUOdTSFgMf1eiJDDG9/iLz2Kr2Go5phnxrIhVvhy+i0fmlkw/flvz1wbMnZz
AnUSV5jFRDKCeGs47gOqcD1D1Y5BKDbd0GOKAP85CJ85SPLZlSMvdlc9/V/3SfIsa7DNkNpZBT+l
ZsBpdcKxFnr1cF5GRB42wZXoJDIuRi4obJE6qcBpf4Fmxv3fdPexFKv7gZujlrXlQEK9xDi0CL9D
nAmUwqrVJfth2vbH8PvVeHPO0NkMsfbF3jpEUbGxGjNtoCYluMz0hDBSS+qnHDynBb/+uf0DF7Su
B8bk5ud5JtXLvh/dY3+S91Imov+7rnc7coLp+inGk8qlfZhkI13FNBxOlFWHuyXiUsLXmKVNaomI
5zQaECmLJnJFnfLghqzOHEWxbLkom/cTp81LkWl0bQQyuNHyipzAzWbOu6uMXbpfbpfTdsrekr8V
D1xHVNmWcdFzVvDAC7tFQOg8HquixHPM31obAYJ9HqN7Gpq4GzU+H1//OtDatmvtKN7sjv4XZAgy
19FxtxDuv3iSnVOdPe6HfDtu6SRKs7ksqoO9VETqtmFyu0oif1wDVvrQ6D/kcq+xQStrbTJ0fAe4
6LtzFXsla0XYa1aXj7Qnls8i/oJahX2lKH1huGnnVSmZpxd2SvXkF1ZCXF28ylFiVrHnP/a6Nmna
jop+M+dJctsImRJEX+YV9v1ItjsRv+4+BGNnAQ/nkuXZcsF7z8TMVq67e2AaTL3ggFCb3AmaSynT
dxncvLVtVISmb2BT6rrKHxGshAomFhVIyOPZXFtU7GaNhM6RjnsK+Dpf0eNpY+H5mCoLHPp9p8ni
p4vUwGMUWhGvPU7ZWMurtZKAKykzV/X7O8ljxkhOqt6T1AqoKPnrvEHKL7YjsiVbHpdtvT0OVPT5
w9XJQo48mydnVzV1cBThL/hES65O/xfTuY/jv1k5m1ykyQ0cJAw7qo3fAi4wDCFy1kguMc9M/UDm
DyeOKB3Cqi20UZ/uPanv+n93D85x+yZIRaYU3CrA8KFHafP6wy4NSNXzJjVw0f/ZzFuZ88fbO9vB
yUNGUJWmSWG/dYF7SxU1bzdbPNBxjN5ERjbrbVHnGMk88aipvkRsRsqHSx9k11idYLZsgSCHI9Oh
f5iBs5wIpgviUtniLniDFtgMdevn5dSb0zn/M2nvNM+3AgSbcnNgbtTXztuZFuGsu4sG1osNn6QJ
OM/a8C+w1j0hE2OqHAEys6jOwlwbSIDBg1RIcIY1k7lUkaHOdWyjzkAtGQPKjZeUtenLhIC8eKq4
MaPaUI0ZfHLv+QcYXmS4kDskEd+mJPfXG/eNKOt3rvETK/iMZuG/tQxD6pNC9++tO3WHHzdWuGf/
i6SW2JpHu/Q8EVJK/FKq7JB1kdhtlWYfkw13IhysanO9totFfEKNLi4/cyKhWmAugNgA/gbrVxSB
y9rLYhg2diJYveDT0cD3wvhEgkdA2CeNi2Pu6+lXdaIaXbKYw61FVG7ZffPpXI6lg+/iwtDzAAd3
HwYS1p81MeuCtTAYeSq53I4yNoQe17gQW3KFBxXi62E4RSdOe2XJmComFQXx8tvrX7RXOLgnBY50
mXIizmyGLpdiD5mRCGbgq76jJZBKom++qmzkiNLSQ4dmMiDDQc3VQEq28uVMc7/2f1JrsVhSLlmi
kRWQJnZrGKFq1a0Ymvu8NNTGGulx/G97L6GbOcOgm53Jod+Rum0LWLoPgcaXqFq9hGYmL52FCcWH
IMYs4AsVs8vVxtNsg9iSaKIsTIEj6iF72zh04kuyQ3lP3o6nstbQDePumkRDRJtdlilAaRwBBlb+
Cmdr10d/BWvy+B4qEhD7XB8IsCm5hbBfZUOKWA5+Qovzd42vFOTDBmSNy0GAddR/nDLhBvmlGNx8
DTEPjEzaFg+0h14JS/XOSYwPyltmjCVkC9hBtxUBuWIq/y8zLS0yPWJWcvRSx6p1VDJd5wrbyGD+
DI74UpNeFZkFiit2jlaW7rDRLr7PT3CaV5pUSDlq//NsVKFrIatUf85mrf0P5e5KhojC6M2d0Xic
vJYiUmD3zBcqEW2RRS8ndHyRPRz6FFOvSxcCYLSIWpNXfGQgEs59P8tWSvQUfiAc00xG4zHzwJ7P
DmVufqjqGxSr6+MFR1f4GepRCBpqMFPNrlCzzE0UH+wk1qOGUWSxH1hz2rUBeCNuKI3J8r9Wp8x+
9E6T1Y5nYLKnkS9iRPIEudwkLQUmxpLkoznzSLhAw7XJCjUaNJvnSw6zzVd7Tqt5U5k4SprNNMOX
Eq7tNhaEYwxH676HSsaLiCIy18FEtHjmsB9C9bxfCTepQwUldavq3rNAuNteM/ylKBdbufQC4jsP
Hc1CI2pGC9eh73sbitlMh6iyqdxOq3iJ/7WKw3XhUO1mCF+0c2vLqm2ZZH9L/fb+uTmRk0nnu23N
fuq4cbVH6cIO2lrieJFKUP0CTamIRmv+aKON2sXM5qYJ/tNsfxxEztq9Qmu67GlBZ1Y9qdi+iZSj
GulfB5vPXed2voxG2Jym8PkIt1V0Efkn+UcASmwpdD+6GhnXYkEeNBbS3SkI8ULJj2XcBh+QfC+w
qjmREjaxDN3Gm3E51r3Li1GcwWHQnLjzJTe++aKSUipXNOFkEYUyMn3hzoJIk0180aTCVDcr480C
vdxIbrnNSuzCaCiepgiHbMTJpvd0GyRLIY1myKL1ZAeLKnB8a6BnBpRFyxNgOKNh+tONDhWhUr2q
iNC+xC01C9d7zL7EwiTgOtEBIH7CwLqf7xi7UjBlc/+bnYoghx4Uo6jh2ZXwkBwoxyRBbGYKe32z
CbUghUW1uJpJSmfTNvySEfvCdyyVYGpScKtpi0MrrelJiTXr/9ZO8VYZJDz4DA3D7XP3+9D/q/20
6bAtBqIxfNCxL9xtjFQ99/BaEyxAqzQUSPYNH4m3jA7AkVWYnjlXe7JlSWxP02KLSJUEzJe9Xpie
jTcFUzwgj940Th3aErh9mGH+IxHE+qnZJtF4YIoK6qLxGazl38aeEBJgSet7KWm1AH7JhQG/8lKD
qorJlcB89SUMSLZdXUI9OjHHX1Ve1TgzWwbIe5gIVy2AynF8KGQeNgCI77rFMmZ3ZYIDaFfb5qro
sH4iWiiJxUT1Q3YqsV4Ql0/tl0m4neDQvrgw6t7Y5+Jw1uVdoaL6gzc7f6OJiBZ09xYDIOKz7zdf
MIUZWhAbi+s01Qr7iOYBhDmitbjuxp6FGqzuSgjrkAczjdvEho04jm4i6L2m1U+5zIviKAnwTadc
cdBazR+02Fpjf+fiYmHFc8ZDTWTMvxQpYtPoBf6s1iRm3goJW8VDDfFq6FmMyujJNzmxAn9jOQiB
AZLr5esVI8NLuifdevMwZaTCxGdZ9hGtHK1vCVifW/bzyCjHmb1ioO2OTaylT+Thy2hsMRG3aSLa
fyVPnI3ffMODstKN5ZQ/K5saCCxyUD6/1cexa687qIdnkjGmmZjxNe5D5ygjwuktYgYaEKLjz3ID
wpIW+IGxTKVxKOsIXD09nXWInw/t9uyUdJkTIXOfu9fJF6P7nLclkcAjKmUQl7aElLq+iP6boKGh
of7eTWYuZjjlaph6QafQcLdueSktbicRJTYnzJEeeCKhEzNv+pDmr5xUvsR8kUtZ0LW1hGFhX6FG
q+fzWPpLoQgdZeazLJOBPJyaWZcC5xYB/HHvsRYI+mgQbFuflOZP6oiH3TadjUkcgKXolZcVmTIw
lU5Uo7RahRC2G2VUcNCWHTV83N69N8QpgUgbKEiLn8M5zLc4mkmTxS1L6twg8XzTqPPHtDQuXqx4
QfLHQN/jZFcIdFtKCphc9jeXqY1pgpnTp+0NREYn6VmbBUGChQodeffD+yZEE/ALjgrkf1+VejBk
SXrFRqf991Xyr30OacUDHabJOP5VOcaL/Q51vU+9xiJt03eDgDZXxUAsF8xn/+FVpKJqP9lW/W6w
i8wWc+mPxghqkpAS05E+E6EUKOEC+44ug1tuRaGz/D4qfm1nMczf+9FfKn1EsMq9CneaZ0q1jdbI
Ijho3HXMabit8K1jcO+T6kOahMuL78bGKO4B0xxrvQHrDFyvDhxy6JjTN1+X3RZ2yqK7ay4CEHNk
gtjLxKolks8JUvTn/FY9G3h5QhNDSc2WSeL43d8qcIzLVbyb4EHuMSsLzd41BUcrmhgakSyyCrnZ
hTdUrZbacIsB4fTCcHD1t1h811j3LgpC5ctFdFCLbdVzJQFjLWtNmBcXVhBrsK/CnsfYmL3UTjg8
JgU9PMbz7Vc82rLEeqHmC5nQQcSTS8gbAFl0Vm1eFqZSH4rvolw7YsAgcPYgyTTOV6J16CoNBou9
SXIS8QtTQM6092iSERikqLyASFqeCZnbWKXzcINtxhwsrHi2/w7EKqYRR+NnFvlMee7wPxWwv0yt
xGfA1BrvwUD124jyzgIOJY4WoocOJTzzrhSS2AvtN6YZMoalXS7Ury4HI6APO2vpWNi4fY7ZOdDr
AN4QFLw6pUFzf8DqfjUpFwmvXwaSvrQQZjEzuhKKKst6Qde5N8Ce7pYKKWYGVcTfn5W08rVCMHaI
n4QMRLG/KP3hJvVuZhrL2Fj3DP6WSil7ZRQCYlSSRa0O4y4n/Ldl2ieW40klIE5XsX5itatxH8aI
FkdsibvwmxESliih0V3TikkhiEJmNJeaMwy54HE5CsJSAxR71YdWOVfuHvjgSzoJ0GMebk9iFiKL
qSpGkwqTXIyQPwWt4M99WAuihebwoqQSvC0AE3v61RMmpMvgafF29j3Wc5BaaIFv9u7nb6Q+PE8i
bsv0rFIzfsJnhqo3Iujtus2LC4YBktcsiosdevEctmbC/3rWtApV2FNLB1dj2Q5tbuj3UUFJO1Tm
64GGnzTAU6lBTlPYLLWrFri5XiTq/BinbnAKWQB1DvFAXlWQW+zhe5dPgF/tj5dNEH1F183M7pYZ
DIfyODlQzM8SbNl9BhtDzYnUe81YOBp+6QEgyejz410RimDBacjAmOfL2OPnghMlWPe6JqYsYLdN
c2gQ2U/G0t6+VDM3/h6EHYHhUo+q582TusOun4PFWeDXcdUtn30xSg9LE7csuoyqI8DQQTBcU9l9
PD0oKm6XiEThueAYYAv+5webkbeOE/KXt33L34be0zn+9BqCMcXT8w7B1Yiz8LOWmAX3xaBDFClV
Kw++riZm3flEePX8nw2OhuKpOP6XTBmwU3BJAeRSAg69M1iQaoaK6p6PyDTXlgndsfY2ofe/klKY
/8YN+PprIcWN8Xha4Eab2W5SdAcmh3zgw3AAs2B0vskV09a5XK23Q28iHW/Dh69Mz5x3/6F93eh7
olDpeaASGbufvr1CqSYtQGZ7g474E1I8qw8c/zZjtnNxE+9wUi7257JCJoNWfym/rDkQWHXt/sKT
IpZN7SfRkFdNrmBlBRgXF+M2Q1o41FOdLF3lbnXBfrOI7ylEtmtSFsqPAjdcygJBiuh9j7fdTQ0d
m43FOsyVZRO9NoptovQga6rU13SUL4iunltxehk7qHeSXgNawtgM8YH/68xJLcLNngaebmPOxDeJ
RcIDtOow5RQGnidABLa3BkgpsyaTeK2ja1/McLnhNKHAMsRpBiF6aV8t8VFGrqnpG7jdRO1/f11t
38Fgo2iPJ7xoGIlX4/cnOcTSTqPCbzLzgE2rjqd6ZQSZzg8d6YjOfmcjqOsj/eFDcAFS3RgCo6iO
BUytpCoZqZtXlVzFj/2toNv1iRUrc0esh/gXLFc3PfXwByApedoY8Scz4jkapTyPJ7wJoaIf9goP
9/tOAe2QqyBlceZq54XyAD/keYgbfe9njPj36ge4GYcVFd38sGzLjjn6lb/vwKVOwl9KioW2beiL
xj70L80W00kb76c/EO5wbBPBs4rbOh+dh4xKh8aqGXlrw3kNXEG6Q01U2/wXULgMCqOtzw/mw7ED
g5t9oS039elERH/q63EC6EffJaIoSTsvMY86qArBjjlWnqTy/68vdGRbsAtmanZWQhlmuvNl79Ra
Yko0sjjLT9KNS2Z7/HxPGikx0SZ2mtUIUtw0ZWd/iqb4aUrsTiMjo0FeRpUI4dUrYI8c7opU1jJn
PmJBiyfp4pSKVEfpkGF5QxCs7JLDw1y53HZTXZX65CXiXKAjbwNg61HFuGWghPEAkShMAeoTt+Xc
qCccr0Dqnghit4tPesnGNT6GFpE02Nw3ACo5XaxP9IRg+8jhAQRO0PNalRkV7EgzsV77AKPSJumZ
xbyUl2d4wpGcnQadahlM9wMEvkoQcyO1lGRYjWPE0dHIJAYQL2t7rlRs8UMRybnV5S5NDZ+epOMQ
y4hkIpRtCQkE9K6f86w4vpSVxkt+3yZdoXQa0QC5THJ1lZWoGXoHpRqsqOHyzivyGjUZ5zgYJAcA
54B/YMlMma0jP51UL+/fTaXHkv5Egd2Judp5KyemIpRyoGprduI76mAmIriLOqMvpeGBSBvzjLpX
tsPPA3P9TZU6ti5OeqlPV6KQP3hOvIOQk8B6OyB37vrIOqgaW7hnTv/2hYAm4rJ0YZaaaG9kkMVF
5Vna6+QGEchTZOVUQZcu4DRC/XWNG88UrcK+sGb5af1Ypm2ESLa+HdxCasqz7njH42n7kjpD/kYK
ehM3LO9oXcnSCJg+q5oP0L6f91J5l7MQ4AtXiUq6PsWJHl5pnhlZluK/3bjXs9lNbhNWxcZUiRzS
6Bl83hCes96LIJMjJY0LoVA+JhaX9Q7sTwhj5DhCNWI+9TviOKeyekNoe4AQW6Ikw7NwAIHVZasn
gxDnm8/xbivydz/e2Dci5YwClb4l5ejMrobY+heh+3fqDMVg6hKbcqRr2mMGgJiPeo930gIkHW4E
yVIHnL5lOIOI1U72/SmFx3QZQQ+kATMd/q6d9QlcYTfNHx/kaCESgvxjndVKqS9GSRFeb9lpzUc2
1HKaHRoOX6yoAKNC8RfvU4LkwtsNF9fYYTHx99YuzqcwENJa37XX4Xq12arRzTXBFI0kJzIlAMr3
OtXrrzF+Vtow4HVjAfs7FEpAjhTZ0HcWHtKfls3EIHFQybZZ/U1I4aHPPrH3VvPlZhRw3M03ZE2y
7OCNO9Uh0clpYveNBDTbmsn32Vx00IYDg0CdCj0nik+z9x0uUb/h46kkQP2GEblhzdmveicZk3AQ
yVLKKXtan4hWF8m1AaT1Nds1IPWSUgby9hwO58dwByD8tYJAOUHV2tlknPwq+OmmSYIFnJH9sjH5
8ESFEjqGwIE76mcPFSz4dhkYzLzH+LEZHLNnVcOqduvdEwu14S7dorSei9xKbDjb2RhlV2/eqs05
lAasHP2ZxscPi6XrRmpLRlNsXUjznEWUDYuyUFoGiPRMRUZHW/I34b5T/EaVUmGPs7EsqiweCldw
PPiw5WJNnvf9ogoyrgJg+PQmYgV6OYR0WPIfHmHnMC8XE5GaVO6yq/Zit7FA44a5Q7oad+jXbyVt
hkz7GwZHxh1gRa5NX3L87DB2Er9+l++SNCnnsyitAx3fzvzR/TVpAiBdGy54yXa7Qqh4kzIYfHoN
0CWAHlGhwqa5dmMPHQnSNUmJDaLUw/XDqSaFvzqbYQ6NyuUwydDNmBO3AKG5XCirhrA9B6Z+WV/p
Gr8+NcRlYsrUXJVOXc6zFj0/mbhOkQ1SnWp0prIclL+M6uigLAooEBZjQw9xrYiGdpBxENNo2gu0
aIr5vMajxEcGHloLYHMesTTJNMK0yp1AQFkNqczGhCEgNgO+3mFdBcREKR6DJLTxTCwp2fHcz825
fHpsS6ujgze/ING05lFQc2pJjelePkz3bqBhJYLDQAaWuDqR50lfzQanS+cFSmlOiMn7POZiYDKo
xlO6g0PX1LLaA8TQpNLOABi/jvAesJgCrEu5kj8j8sL6lzOYyGZb8s6y0uzmWBhHwLd0hJZiZD0V
+2twHiNyl6y1fub+gg3Q15kkrBOelxUwUvOrPN2AgFAvhScJKCajWWGiOokO7B7fBJ8yFWqb+AkF
9AmUkMzQVhN/Xo6DExmTrW0vBvRc22k6VbE3VrULwvJdk4QCSf5lt8KJvciExDEkRiX565wuoe3a
meHNDFqhwXKxFswZ3wFbcBImWFdPj4uOivzgAZTH5R09JUR37TUJoLcnflhSyFmuMjC7afxx3ftu
vhma6rMj8sZIg41ZmnVrUlgkvNtR/CGq553/1RcdI4eLMWFeoGAlbTUxPguErcyVUGLjTVESJecG
gQdUndUEFqUrvQuO4fNxP8RDt8dYWIHJ6GAsufoBv7eP72+PXnMnjYkhZCHKsoQucWYE+bp4T3cQ
Nkwp9AQBi/i0dyC51Q3pBPfpgsFXd8COf6ngXp1a70GUx4aJ/YoJIwq6ivFPH4TmmobCANlvevHD
5oC2q9vx9eRYFydeCsirycLKpvKJSLlcuJWBUgTBndeJ8WRlgfiCXjkzOLL35sRfy0mAySaUMtWT
vXPUqMDdD7Lutwg0mxMDj6okkxr+qWvdYmpS23eX78I7kVoTiUYDpfFRY9WqFGZpohHx4oUAU72C
UAuyu2rGIjAN6tWnCVKs0Emq+oZZkHC2VKw4Og9CoTrzjZnqpYPBqsTS++Q7eMl0ACa6X12lTcYU
Cf1cfFjlnW2tOyGV3dT49FDiND1q8TladdzGWadEKc2dDklpirvJzMul2srX0Q7mC/dnUXjf3Mtw
mDezNurg5FGx86vtf1goqzIY02vBDH7CjAYA4ItGUPeschiiwTKMIQOhQ9bgYxi76PzSA9uLBdHf
5NITZhhuBLOdSfqWSp23BGmhDLKMsGv/MsfVHo3FBu3kGbAXQuvEdch7IBYf+u+OpCRq1AfhF0V4
GhsZ3HnroUrOGegx+YscT2LZ7PJtpmPGfOTgBkLSrUN4k9Ka759KmJTKhKtXrv/cJ3Z6LWuxoe/3
dqjjfG5mykvFZUHbqHLto9RizipRMI+A+oG1mFNJR+/0g2xHMawcfVBaF98GSvb9d0VTjsfF+gq7
kqXUjtKud2523C2angiJEbuJrgG1xI7xu1Q7MpB44HgmYOzwf/sn3AJj+/WHxWRohA/BrcZ7n3sv
My9kZj867n2N6sH0XTMoypQBpxbzl4AOIrycL72oa4ef8dqTrFf5BFRj4glt94Muy9V1RLMSlqQw
n/eG/YvFkQEglVY7lzWxcZgBQId0E/3zhPUsNob3QSBBdaR51+scgjkOlUgxxXhdlhpTq2UKTKUW
e9sP1BRkpLnGX6/Cx2k0mjFg9Tq7ABvgQ0KU5JlmijhfULXjbY2YIj0NazzVDmpALBCHsBaar2UR
85ztNHjJJBzIB6Zflf18W4utlN3jJne4LwLiYwxlpGAfJZi7a8mREq0HjaOOsEV4jqPVAX3/yU9P
dt974LzAX4gLuHuY9Rylx7AMtSvg3QowwEPfpxDkL7LuW+YCRPvRXaMcB0r0Rb6a+bceQhCq8jw/
iNs38XQlwzcO7SGsTNcP3OgjqqYR/QUYdsyK6OBxbToSB5jzMilv8TOciJXecpJCnBvZQQ6/5s4Y
cC6GZgryq+bnLK5fWkpbY4Kpfn7ntrubg/aSENTQMxf3SEUDzXBookzbTu4Fyfi0T2A8abwreD6q
4D8Pr5JwZWRPHSYySGV9WvMyOPLGpynBGwmDl40+G4gwr36Z/1SaDXWPYv42215L61I4Wamayfxf
+WvBucQF706hXq9K/BpcrJi7nG8NHKcfdVSirLsVabx82wy634kOBsuMdJxyNPkgvYK/RE7p4uur
OQX0E86JOJogMSWgIPrrIKd/QoRPp9aePcdU0WNwZWvfjFG1M2mTATPge4cv5QBw7r0UmJ6lAm1b
qk8DpyHY9jmrenp8cHk8eE6DJiqBE5aKrtVZxAxUSF6L06XXAKvtwV+tFiAiQAA2uEDhHlWC+3Ke
hY2+4ZxO5KJdGY0zHPX44gdocQ8YCDWlEDUuRNYJPg9onAWO+Gr/+RWy6cN6X9U/YFv2SyKsgIBs
B/nLa1/B2EfGc49R+1mHn18cIosLhCWRT+YNGQ5BKLC2iIjMF1Ii5LxMdk4jGOnnZg35EyAOD613
s6yMzYrCW5CRyAQLbxs3pmE7SMgY1kofFShOMHUtfsi+I4XwN9ufhVZBZG1E1NIuxT1UFiVrPF19
NuiaU//miAkHU6yPeyKPZuqu3+vBClOpEyLRJsMfiXQwSvbKOK+j4vi8qdc6Sec9oEbx/+V9jX70
qxFVxdK1RxWJyD3tJp9lQCAM7ZJ1xfAL4uI8lRLjOUjPEOvfl1vH12PSRKyzJFUBquh1j6JnbQ+W
g2i3xXaihIPpHIRF9PYAk3Kx+ijuYZ+yWHXkpw1FRnliqnbIOWWSCeLoTpGYOJB1fzsDTrqSLNju
MUgNmbnlQGfHOuzL+Htzv3tJim274KiK7KodLeV3GWYapxcqYL5UnCpXITJ4d45d9a5y86PXKCwv
23WvZxyGsQlQ3jSACOzkAJti/53NGmhRWfiYDmcxHlU1Of0/O2dQtmp+E1Lf0WeKJ4SpykSzTbQT
pyOSp6VcagD+V35LS9VnGB0LdsIczloyHNGKCiZgSrNXCQ0gXHKj324kv2GQAFKh1CGyRY0BAw5a
U2emfDCRiYaAEPVriN5krl0e9gxUSWrAWPvFffROY2QJnyikJo8yg6H7b39A+ypPV+UvixwBFXk7
3urvZyKaMSZftnJx5C/rqWf5VBvZkwz/2Ub8+R/fag6WEgWyfLsnDd3u4oCUWc5OoofevFdWuyqC
SFsX8wbLTJm359niuzC1DuNwiMR1gFT2DxLxFhln7WnVSvGyPEgFbibahVLxz/0DnSgIv299Izh3
/lVCos7kn6sKjOazCHJMgfpMBSIXqlzRchFTGCFuUR4iaPcFRz4UG32AigkWoabVgi1TjftNl3dE
I6Ku9AU2v/a6b/XSmh66Y6HH5juhLxnv/Xm9wq2E8+WtalBLlkrNBxNoO4vt+cuMxiwq7IWxxqOx
t2zjmDOwtsIcqcbsNGRKIHt4tqGgBuUfnFhhTXhMHIAKvgDf/0tqOX7MXpX+Nf1KJCKRWdRTdmhr
BdP3OILZOls0uHLuPtEor5SJDVUjh9+NKUui5pOfvHeph5a0q3t9zyYLab7Hihpbifrte9V5R6gV
mlRP2MwGialrVzLWZpQ4sQ1uC/fqlmNj6nvWJz3oJyxDdkSwnYU7CL4VRl0rCWydOwOPXsmb08G9
C9VsAIqh4EWz4Pp5scj7WlIOLLEskZB29lu8BzwXCc+ZEI1F2o+DBV/2wwFsn8rx4shc3XqFIync
7bgKsljwnXAaFTWdRoq7v7I1A2izonC7+Lg+3wTG7yVfArcxnjO2EKjItHFs5vohCR8C3oRQ6crT
YHK0LokfSwXDqX2w/uCJPzMt4QzAKg2QWYm7WmaUdb+6imXxL00E8o81DjL/Lbv9Ut99zZyhc/RO
Uih2DXSui4K3slleF424HLX6l4/ldn7LXsk347PH4Sx1+Ds4PX6GvtaGWdVFdQUmM3qowdLZJOL6
wSYRz5qvW/3qBCwpcbThR+UA1Vw6e46XCgx4oMeKBZ2hEphu350LsI7sUboJnIC9boYqX2zKWqIb
rScf9yZSGriHbPbB/K4GC80i0XEpOv3rC9EVMRQ+bwY7GQeWNy4FsygogLxGkezaUgU6BA/Tc8kx
GHll4O4xDilj2lBNBZzL/jiVxaIVMRCZUBDAH38Wx85Mv2I9raoi9Uq16I8PBLVX5Igr8HZ1hlkz
c2V9UBJsWPNu7tey4U28uNEf24sjiklCrEtWYSbdUpDFDy4MKpC3BF/Ak9g5J7erBtKwnBFA28iN
PtfPMy/olvjia7Cy+SSIRCvTJw3iLAk25opCXJ6L/ENrdHkNBQFwtvYO2D+xd31FULfTrL6hLMrK
Ros/Lcee/AcYsQ76bcCiWEUqqMp0dYMy88Ik1sHG54r5XRWT2jqTK3zDgDobf4VXGla2JXrJf4Sy
7l7DVhvVopZViyX6d2fuNOFohmTp/cYgZAMe+geU1IWjfIKgD7y6C9Ww5PDpeTqLikKKUeaVGM7Y
X79nspo4dwboOVHHQ4M51z6OZKUOzWsTbCwGFhh8us3cKGGmoICGTnfhza7FsaZh0/XGAHROPw+K
TMgv6cv00xc8rvUbOr8tkMOldmlasr8Z54DZuAxYmaa98DquJZWOfCWeWmEb0xzGAiH+C/KLRA2R
tvBEXy5R+ExGzpRx1wOq5Un1/y+QJadvDLax4gMdlcBfCZT6RQk55PPRwcEynLiFMJ7qlCKzirDA
/2ckPTrmEKOJzNFyxUK81pGMkxZAALGvo2mm2ij4RxrkHRrfgA1TjZcUA0/isQRsHR6yMRr1FWr9
KfbIKgrM5ztqdtQjG4pu5Vg+hhaSftevDsI5Z6vC0O6wjMUBALfIoiqGdu8zh0uuntHmkAFq+Y41
moylzbGIt2s27jYZ8CWKaLvBN9KGiSN2i1GPtA0ugmc11S0BleMt5jS9LX2i1afcxH6dfHOYJevt
5cEgjQmUCVk2LFi+JRiT1MNmQamGRWuBZpAVUENyjIxjhlLXoL/zLvhFy/gPb/F4J1ycOP38IgFw
0S6JrJsq1AtNCVh3K+GGpH2yaHYx9jF6FntPRL6ePNccaXMyi1LbhuEXbFwdybh77zVa2jGrUkT6
MDXb+lYoUYl0rn3Q9ohqb5HVMlJ0H5bGdymb2u1vafvChD9na1rFfuHaEnDViiV5aF3ijl4xgn1e
rYtdIRV6uCtfQsxKQ29gX7yZ0I6bsLtMWaVQ3aRhyXaC/tWgzernlhbD+kXs/gPSY9gTPqDi7DJX
VehMNq8CwQbyRceLI5TITI9ZOTsnluL9mMR7ZAeas8tMGNm6Xg4R8XDqTlvY89t0WNS4CswKVNbg
0amTsx+1hVE+vTBbys33VGooSALZcmUQQsyEbLfkKaN/wmzZ1biAOZt8vWDHYurQcSChVr4L6e1d
sgE7VcxzouT6fSE2Y//XmGDmby5+6RB1SihFCEbO4qDDRQQf2784qridOxs+HpWr5qWYzKjh4OWr
EoiZRl8tQGXYC/mIo6texyjseMa3ZT8tBNQWUqXtglNujAz93wTeZ66RVe/1dgtebY7nzTHAuYsM
tg0BwItVdfK+vL24amVOKvWSgSBQvaCTypDt7/kSZrrUHULJWNm87SoXyfZ9bf+Fx+zfuMrPqT/o
XViSSvmYQ8XYlIr+7VT7pCsD9E6sMA3iKXmNI1NK1biXcFoPFw1LE5mVEoxwJHnEMe8vcp5Hyw7D
53s4P103eqbj/nj4dHRvWBs9W9AL2xuJaA3Vsc7ESIXgK9H5XPGi1woTjHAfpdrAGR0vO7gJB2um
1VuUo73UPVBI6aXAhYFJJtfX2+FCxrzcEs+wTi2/4gQw9CqnvQz43jxiIIBLQXp9+JT9JFxUqQP4
ikj8DSiSYxJ6+QSVV5ZRUa/Yvllr2NL2tjHvUAteqgCByaPDxXwg6Gm6yEvgjXxCzP4Kv5XRjYr8
PIexFEbL277gzWroEFJiz3FY/ek+oidZQsVmDf6OZZMHprC5X0htnF+yufTIbfV+RrNZLVUujaDH
VkAlGtZASWOy4lZy80ipWh79pV/ONXlPq+bpwUhh1s3fX8rtR5gr/lOHuBMjNll2WLTnUNX/2Cqp
uhYzI/VVrP2nNEYE5emXjfwWdg+jbJpzeErTrFnma28rOuzovHS6vFrPexoTJtZR8M5433iV+cNw
wZF6MQzGSo3jRd8E8vCkqvCwqR1UqfHPgwwFn8Yw0q/0pBgSFukRzlDG4e5cbtA/vSS1rCN1nQca
tmDdOimxsfIyiQDPza2sIe0WqAY3rb1ifnWR7uDssQkeScpcVLNL8OI97D07wY4vWq2Cbji3rUha
MQYg8C6hbdIII4GlPsZT3lao/HCz+foLj2aHXDG6dGeMenlAPUIwQySa/5W+RqHzN/O+NIcnt7Mf
RlYRViWGxbOT04WGwNI4VGg4gv6c0nVi8CPV2955ZdFsboHf7dna/Lb5auI7SAOQreNwtNpj5ZyJ
NsekBMUGXQrVbm68SK/lK7uLTn3ZvgD0Jn2kCcsC41wM9Fq+lJjwvOKZi7GIMiUpR6TCfAMpVUBR
Upm2hDhqsLIUuj6MyfWloCC8Co1yQFptldpiVP5Bg2yE1aj908L/7YnVg7shqTfgXtWjAE1L+luY
YCmUmu8gRxacHPe4UdtpRaieu8FMCCuey/L0ACmTKygOd/ommipqkF/YHmzdwLPUfTaqi5Gn1ot3
L60SJBUQX0ncoc5YTx0rRIMN/w0fHrYBBh1DsUoGJmjvLqf2K1WjPvAkJzzPkqA7aAEoA1D3nKSk
XGpy2AfdkNtxo4mE+W6pKGsCmSRBdCww/URTzSifMQRbJ/VVJvNHz7+Tn5exW1AKioM+ev5dhBhE
9kvbYTBwK8J2hM3oz1/lxIGAeOOzRgJBtDrg7nNGe5/E40Gr27Qay9fBclyColzWzanY9iwJkff8
tjyuhS0uPwT6NB3V/wiP3aaQXCbWRwllx53aOZrDVQZC//vlIMgMVROagkkQigPqg0D1kcmZCgDi
3vHeiERDBQV2m133EmJo8fEuGcFT1cNhc1GUcHKW1RKx1nLSjZMIWnLQudm4ORSdgjvUDrakmFeo
4JOzosLuB84PH5km5f9g3zEvM22YXQxpbEDkuIcUrn7aCNXW/zjTNTrW0DMcPOvYHsxuaedqbFPR
/gcDKYh+byEeOnCSq2Zy11dj3kbfpMe1AbynrTFrEIN9/LNW3QbOGXHKJQCN+6vhrj0gKFSEfEYE
r+ynCCbE1bxQQ2bI5d12ywwcFqxUkcuaiMdlC0Avfd6XWJVpu3CvzgqXQTX+DQAwPOPFgzdhNcS3
SY7wcXmLkodt8yHJ9AoGRT85JPdLnlxMiZ0iLj6dUrRXTtYCUPKVVH7Lmu3NKxa9TKy1ilPklm1R
Z3JlU0VRfJ0feNj4AwEJ+KIAlj1AQ+nO0z9+44/k3sPVsJSNQ3j6tBBpvkNBqnQPq+hMvaNUEuv7
VPtAO/cR2kr1frtQTDVRpJrAWr3Qgy0J3R2R0ZqYPVUvs7Y/bMYf3b74QZ7rUZrf15THa+1mPbU0
yNixH/IkeuANj1KbJJ5+ptbYKTShgJ3JlbxJlNH5J4jmdmyFhPXsBNkWLPyxfsv4IHV1lYCaLhIo
CMr+FUOw6dGV4gq8GgVxktUALO1X1/ZSj8443aYl1V0Io3Imf4eDBWibYbi4CzpZvyyNxR+fYXXS
Dxkvje3UX+javOZfvrXSy4oEmkRH/f5RIDFFoGuICzZilNpeKBDgovUkbz21LB17mNgndEcKxpfp
ERUfv9E1ZFEXvWW/gJmiN61HKN7kZtqKHDH7pjSxWonHQY3Q50xyAvbWyfTCkD8JvqMyv5VHzg0V
PCdG04XLeumEn63TvYrRXz6IA0TiAOg4e/WRir5QKEFlG6Q5kq7OSaOuRgi8mGG3BL41VsgJO+Rf
0MLO/rz7EYa5Dl4qA5waLINrQHixrDOeU2nx36VFgxDIi0xnI7blx07gKwW0fyoNQESYS4+9OPNB
XlMVF2Nv5s0PmHFF/LnIukyZvZKfMCiHdOrdvRv8xCT+nZaM3IUA4tirvJehG33ot4gDvc5Iw+TI
OmT+ifRm2XVaIVQuRIHq9XkE+s7kMdgX0f10R393+SlB/+Ed5n4OEuIGd/flMLNQJBU3OCWWizfL
YTuZogifFJnlQ9AGpgXgrG60ldJfjt52ZAiMuTJZdcPnObcYTV423vp9+Og5OWhlmV9MnfYLuTJX
ofLtw3EIDgQ8nek9i+51jGi4HsRwufsT2FEWJtWoAjpIkcxHjOeIbRh71UuYXTbk6O+bU8EZoyb9
uwKzJdeOEpw8c4ZiUzxULmFwezcdezzGQrv/zZ4vD2uU0gDdbeEG/YiaKKNeaf9VsN0+pLUJAWUE
wespPMo0d3VGJUgCWmtf8jUmXUanKq2WUFLf7kzKfJjrsr8YyIjComL9ymSUIjWquxmKO6pnGceY
zBd6yTHdlUjlfuSZ5a+nECraiFmHxiYA98PJ5X3uilavuXheMpPduCtzan4eZaLsLEVTR62lEwCM
T63fTLQaMx3w7mYMk1bcRPfoqoT9jXBWPHwKpW0cljsSm5o8V9H6hiy+CbgD4zeHL6L9iGtqWMDA
vd4M0KAvFipaoJwIcv8F3OAIZbiN0zVZjKmAf9nAwOtWv/snYde+/gSKQY1dWMzHxsC0DcbpoUHg
uw2EsROWMwyDgKh2l7jPOn8b8A8G1+qJAm4D+WjDL5ZwEdUzDpH+U7H81Wgh+aZG6JVnkgbc/gtD
rJ64HYKioz4F90NZRbEzYGTFVkG1ge7qrkX827QfvzzWdn8WpTbF4lWyuMUMyLIC/QrdpVBLnwD2
d0t+iRv1mmAWZtB49OWUCpkHahzMssrQJlWwTK4PTNrGz+fQ4r608kG1dCuPCrWqvv2m6f+/q+V9
fzSiRRdgxZSmRhQQ5U9R7HTpbNPRplDRhS8bck1GpQA1WBlW5CwZtMp1HzgqxRAVoLfXhGTC92dq
fgKjvT3n2dXoQJghRvxTbNQejvb662Up/zdC11dkyVysWw6Pjpzu0Lo6adcyb3irCvlw2LQSU9F3
0Hpk/Ue7s1PORA1ezhfKDNGgs1GEp9lJVmfDW7nB21S+F08bVWahrZOMN13EIyF5665UeGrgJlpA
XnB8e6UItEc1FIA35Mi9z1UCIDsbFVS+2lfGTY6lhfNkjpacz4nDW4Pj/CRBTsojHgcH9oTool23
0lEzAoL0aQm+hRg1UZhl0Jn+97Suq1YbjIsICDR3cR1TKkZ8JYRIzmQa7WvB28c1luEKbIo5ofIx
pLWVeZz9azBcz08wvpRgZjcYdasDdVNoTR2S0NVZfAaiF1o7T+W1aaEnUcWbQUpwOqKTopAPolcB
PAHRQJDcZFU2h2rGEJtNytu25aAXbsUx8v2uUSzuGLmZMexWw3WZVX1V6dQXsseTYWR7Uz92uzC2
WsNNK2PDXi+Ch01vGQk0gTUqgGSjrcYBobMmvAs3w7rlR+zkWwjooCSC14XorXRUPw48cQD3oUDw
iC98eSo3UvkcAVx7SRIvQ52myF/Hv4wNtWzG2PCXOKo0AZjjAPk4L5CKG8ibo+1kRNy0BeEgRlWj
+H7s8X6W773fia2cuwrTbJ4Idnvq/2kZ9izel3VfoU18stfhy6eGa5KIzEb4mHJurbPsGQLOzg7M
Nb9lJK2eQMjXxKHbiwftM0/3KUQp0m4gOJev9bzfYb/vyJh84lDoH913farGBFvt6y4HGUOrbyyQ
xeUBOXvJauywoxqcRkd5Pt+LfoJ+fDSUmQsW10rPgoFBmNKzLi3Lv7Y/UUN0LhvFqjjVDiiUjKTM
DJMMBU9Ou0IaunKmgEJHbnRqLTXTIWquAwRqqZD8qdMMhoyLLcZ8Z2tsiJUV1zhhVpwKHK3cnqx5
Jbhy0FfziwJL+S6mkLIrKMth37JYaQIkmCC5lDv4UJw0oRifXuW2FFlae4Mz2P3B2fLfWScXOchr
T7L55tmQ/2f+HvFZYS1hb5vSZ+L9dxVlFs6VM9nEXkK14o3hUc9L8YupO6I/Eskicbhafdj1/Nu2
gxRmkJCngFHYzwBHn8n99oT9JAoj0AB0YnN66YZS6tOdBoxa7ueQdwBOfr2TwuKsDMg+X65Vfl6M
BI1mtO3nc6IICDAvoQeA8FQPqeBs1MomqZfZnNFtr3aHck+gqvwdQo90BHDzqseD7bPkXb4dDGGb
4IMI3b6K5qM4PBJFQTibEtHK2d9r5zTIm9RK6QfyTBWxpBpkrSj88wymVun9r9iT6hkN3WyaOxzV
dwrCIRuM9FN87ZX0pJYp5FbWuMV3ZDrkqzU0PJl3tbvsUqXltFisCZrxJvu+sOvgvabzlzh0iEBl
MZz7fvziYXPtCOGajgI3aaLISFLq2RUxPO3N0+Egqk/ZMDoQTIpq9EXxAF/39rrREKqjhRctVOzJ
Ggb6AO0iNQpwnUn2Hd7tcyVZmW3QRVd4xPWlr/RnGcwrlFsrLB9VuW7VvzAOQUGJ+lv8c8cx3BMH
XI+DXhyZXjxvW/fCec7hfc7+XjCSCxMh5bUTfypkCrDVCfoSchRAw0+Q/zGkxrcJVeS9SHdUBdIH
BeRIeI8pnvpasIk2tkW6VKicK+pi+XwkH6opSW4dKg0/es8pq/nFK9xT147wqY7FgDTAWLDvd9Ad
2nxeVYVuT4WjOSYwjO7mYAD49ueqq7QYv5QvmTO3w+PifLk2QcBLznlMfE3Gzj0y0S1dqoeZ8eT6
xCBZTVB46ZeIJ0TYh/vW4ZHzSMf6Axi7ABJTC6kj8KBRZomU+0vGRbWlqUdi2k+9ClrJo/8kfYge
8b7vZDQaTrF5sux7etWvKG7bI61vfJ/puyklwxDwAdh2t5ypOcm5Si3iV9/KHX73chR8CJHdWJBU
IrW1bYOArEvme5ZlKscvpWtprK2ONbbp77fAQFx2JMguNDtzupRg18I/GGYLTGLmZK4DfALBfM4C
3s545jssvnAh6OZD9ohGyuQkAiirLDZOJAHLoR2Trpjf7f/GUS+bH9sWC/eFCyG9R0JDN3aAoTBs
dHZtsrIUtGFSTzMJLv6T+mmU0yL7MToCI6mQq7+uu9oidUdUF/WKsvssKNrhGqyut3W6FzR/Lqa0
nC0pHdRDN1+VopDpSAF2Rp9BNqIUWqrVKnQzsvKZk1ezIPcSkM4IFUIcxBZWHctITVvkJL3W4sTl
ICkOddHNMq+FgzRODGV3yi3CntrFGqgLz+9uUuGU9HOhfZb7TWyknCYkA09MauQ4tpfkTTCQI4D6
mI3y1JPI5kXl7xmJIx/Upzl3os87rlwjOGmqakKpKSiYhobHJkAZwN2qTJqLahQRF190tLjWq6op
ldxgkliMzP6NaoVELGspxM8G3/imDwEj7ejarAm0Mu2VtJv8iZUyKEbjyoDxD10BotrKwmjYhQ3f
8Zljh6//DCtNYbs3MabcuyL/IQ32sNOGZ3ackOWkJXFkr6AcIS0UDDL0vejtrUgQjjnA+V+OhEN1
Hcb2Vhhvbn6h6qWwC4CCq+ZgI0Vg3wzY2ayTa9F4stpdLXolO0xHNyoI1JMWYNROQ/Z1PVt9ngNN
2ZAwftPyh0Z2U92pKT1ys2upXt2OmyW0s8H/QQRn3feujkiuVZpkIszybjMgnPzwjSRaFTC6reMT
CxzKyGIa9mO71lriW4ifZGxGG71I8VedFiOElUEWHpbl/GDVJLilpKpkl48gQtCeL2SHrhbImk9F
Ro3lNbC5uR9kG/X/LnSeRyxVdasvwvtOi7tl/d75uvnQmQVOG2VQqohLFC38a1uyk8Z4Ohyc5CfY
JUv7M4ZKiGKgPz/hoENp6z8nJrRKMRHTd6yuHwmMCOaSS1FgyiDHOwPqiAHbbo9htcIUQV6o0wd7
ugHuRUCg7hIXN4ZNdKqETYWo8dP9tcVhirbQrVEhQPc3OHC1xdiSoQEEaS1XtytLvz3ix9LzVcrd
c68lsufCYqAT3rZSFhgYL7IClmI0G2RckUFJXW4uDSnMS7l504ydGa87bw8+uRP5C9nVPvU2//w9
utcFoDajZQf2PML+R8ANzAmkL2yHR6rrx4Goy0xH4ywQVrGXmzERON8f2gqifccjv/pvIiXVzQyH
/eVloC5GYB9rMB0VIWHpVDmw8lb2t+syGoxaS21FPD0MSae1r9Vs1aN3I3hbCCmag8Z7sRmt2Sr4
ENQgCnuQprwJfirsh07hFqm2RqT0icxxDTQdsIen2Jw0xcDbOR5x8oNQdlqGIyd8AS/BLiaXoBuD
xLVzT3vOjLCQEtCcVdx8Ww5eusqm6/nqbhhbOgyjVd1Pd4rbh1ZywghyoV7KxL+JkKIkjekDobBb
uEitO+SDsMvaWtk+wXxQNPHnxWbf8ykzaytq49wrb/92XfIwLcHWfMT4aQ4emGDfLJgAP7mh99ax
OZRMd9DoxAmlgOqC+dReXpqD+MWnbNHFopVOWZAzZp8ZZzcj8ED0XlGj2968zTALOQa+FSEjir8b
PnjCW43u2PZ7P5jKMYFvG+WgKA89r1NKNKblSsilpPyLnweKBuUsH2u8XGeunmKCCWDLhgsbStXk
WUlZrqlliN7tqhriHt+sns/mbeN98EHAZJJh3CIERmP/i7b2Q0Rp1T0fc3ON8ngmu23gVT5O7s0d
eIS9fARIlsasRnsEcpAy+I0dwk2M8VlXsxwqw4pIhC9DIKG5Q9UgHLjRAQskbeQ18Y5o20Q7bt1l
UxR+j7yuYLHtiMy6HqNaPuejusfW2RzEHu4CtLXF+9hkeywzGSKq2FjSnIZ4Hv17Vk+Dg4SqG4X5
bY8FAGJ00b/maLT+oIgDBBpikETDKeTT6c6wTqH6mGvYaVRHBsBFwxsxjg89jsV/TbZi8CFWgtH+
ig5C4U1HCUm/KPcyxi0eBNf5TNUj3L8V3XIdgD8MupopWw0B0w6LGPqP545mhal24QfzzpdWg6vC
kIvRnuVhrncI3/Z5stXYU7rH7CE7xPQLKj9h3E9oGY1AARQ7I8Emdg2tcM0Ra2FKn3M481VQvNTy
ZtaLWu3nG2aC/yAswrRupwA16ngeiPLL59gbUdr2B++6BdX9buAKKWaOwU6fktNXk2fRufNmmAC5
CPc8wBSAubhmxoU4pz5143/PCPH9TAkqLBuC4FxnyGV/aJXhjaQn6i2cpaMrZd5F7zA4DjVM5ZxA
/+03h8zvxyu8agpTfLER/AYkr5vt9+UOHt1zXFpr6N3aKQW2eruNwZ7IBgpqj/dbsqDCY6yAYPqo
XvOXgNg8tE+sE2YlA4/f6XoFYS3/o/ZoflZksY825OrOFbmFAk7vIy0ZBZQJVx3tALGlQ56pRV4n
1ZA2tc1h8tKZmQSrH1m+hQRVAuEfXZQiw1k0pcYrYedCiMMkDu22830izqkX8qXoz44sczNNov9D
gz85gh6DIcmhATE/L/TApLc3xTAO0UYpGsSMaZFmD8CHIUJs1IlEVNp7ShBDOqWptO0CESvfNB4L
AIe484kxXU7jeObrdGbSxpINE/tz9XqWdX1RAxsCbGHkcf7TKAu6No4lD2Kuqqqa2LUkU8ZvzIjJ
xAnVmOPKVw6BO8KSul19T/BrLiwHzcBGLul3GSdXTq08gw5E94Mq01aZ2a1atOBqELJdTizZ8Wut
5L/YvvpLpeg61Qgx4s64QIUXDLFlYoh4mjQqIbxqj3FieVSP8uE69zU0MhHKmGBCzIOJ0nuufft2
2a6azG1q8SD/fmSCog4hGmsa8Zze+IB39XLbQx4k79zVLwDgmrvfl6nFDqAugieiYnmmh9KxGhnK
/Ig25LpFCXYupIN2kD273i1nvcE35j2HjKydmTGk07Qk5CF6+1pLEL5miOsXd2qWN0myFFHQV8cJ
u1AJfzTC04gbytGmLybzOLAEHugnevnTWBn1fv4GsuyjjqxR1SEHn6wRngEywK2MLsn46B3W5vld
5OYHvgx9HXlozGMgHoUExKxbjCOnLz03IzvzqlKKOqbljTyCydQR4VlxoK+sZCGVYRgFm3X3vUGZ
v04oSWpP/ZeeC3gYY4kazvvvxjk+Oczas5N2RnE5SDN4JoiFAX7nssNMPyQEbUoR5r93vM2SM8Bh
0omcNKW3cIdvhlxpmlmStJcR7zCN69g5stLiqVqPtZk2Fu/GjUrjbahGs+QHnqyvt1ILQretodIU
WM/EeqVLsyti4483NH2pe+hKYSPBRzbAlW3nFSgalu7XuT0psxSvC62sCjc8/qcv2jF6PaaJsnZy
SHbTdXAXiTaKrO9hxIsV5sMUemMb7E6BBBx89W8EaEOtHC62Mp0GyE8E61rIfFMpHneaL2Jj5kB7
24GJoDmWyJH6HQFc40JFQAwuB1nixJUw9CA7xG7p1pMqS0ot6SLHotoI78qEvRT4o+oIZpgiUuGN
XflAVcJis+cz1iODyQ34ZRfjcX2iTnAh/HBSSuCKU8/Ebtm5d4kIdBVZMtE5tFhLO4a/dcV0fFay
7ElayaWomKT4yWzhumMXWDPx7Dd/XWxuUeHiXrNTg/XSPv2YBsgEbpE0K2f5TqPEUGDfYii/iK2O
IVXf6iGw4kmadBFUrn45GeUB6S10T4fKFUZKaqX4c7C1I9FjetX0EwUT1+km4b8rYjFitLNgsN2l
yeXOY5MWrQpxAiDkQvmb98pXSKmKp6myujU6ymoMTGGzDJao37x90Jjt88cnPo/X6sjhWCwcUPZm
cPNrbwWwjJrSKMT6YJeDIzlJjyAXr3hN4sWyXWoByE9bl5jkH9YhRBJDS+SFR9vvcXJpXqqwqoT1
uEus4QtmM2PljwFSueFVknsvVTmrkDypiIolIppEkcY7WxIJOxeAftWqZd91M7IEa18F6ZwruTfY
8AWb4/IWmVXlz6Tz4GQfjgcJxki4YIXklSa8Z5rTit2K1J/NqVxkM0QaxlkER/ogrVdMzGcBIqIC
EObwvmvZCGNrcdRBs4H9UAa85uPSN28iOY3fpEjoQIP6pCHrDye82SZVQXx4IUiTHV8/9Q40mXsy
JAMXv7NYHk73+AJaYe+Ybr/WCZmb06WlRh8rgpU2dl433PacTsvF9pwLZZGuvUswkaSlnPygLYqr
/vYmjQLW7juxhJRlje5wMGvTTnwGz54O2tWCNJjaxOUZoXZeKwQVkbpv5xEQFL1gjmj+HCQ+s3FY
aOSAnozyYmy7zH43L/2JKMqRyQ6y4+uQvAhgtZrSnQfpKUnz2k9Gl8K3D1tpGWNeFDjJKJHBA600
FvJDLWj3m7groHnyzBgNGCtHQJUFi8UHWbSQ380kEOxWdfnzRYWb06TaX50L7sFwL2/2p80zWvX5
TdFIvm7sfbFQaGn6Rgg5duLRd67YBXnw8wVF/jmCr7jvP6XoXqHkp0tnCtAY0GnaxZOUNGW0iCW3
Zc4QiITxoa19glN2aWx/x4OngnMJKn5j7+8nScTq3BbLTVFnmeU4+OaW0+Mb3IEH+PxTgSUzuhwf
K+4FDq6LW2/Fzv21EqJZBd99o0weY3PCfOVAqC5yhvDJ0FMWFXJVMZKS8zfjdCN7/9f8jSSv0enx
h0cfN9MMSK6QMx/YRnqAVV/ZEhZc2hpPDEa9xNcDFJRwyxPg5+LLUOWb6Taf8o3h+NJiDINKU7pi
+wMtbUx1a6vvUk9GkBcNIjKjklwa+WVAzPlL4btAiFHWfOLnrRDLd5JkZmYHTq0k6Zn5yiPEqmyK
UTbJ31OGkAB7SPsWObMvDyw6mmBab7ORpeWjZ5KYYT3XADBa96epBbaOrT+QQGMerfFTYFBw8+8L
J1Dt+tvx7DOBCFpzLzYjWu10TldKSAeBEQBTFCHVboamIR49RdzDnjFbINpTsk1Vf5PSV/++rPBN
mLU3sbxIAzmwWQEeK2wk9Nx6mVvfZbKWlzr0knC5QFU1YVaE3cIchA6MAPSdMBzplOIdhlMGBvo/
DrIFBQs+Egkqvy50OI/aMNZbhcrLLpCMzKx6T96oqdHo2qlpZKzKpUL3hhAwDeOOjkWZSLsJHVpE
xnMWDzPzKHjK1VaTI9ftfQHVg3wX5Ekn64Cmo4QlhzzMFLC/aO7BB6qOjgnmOpvtSX5+r/6hJ7Fc
YVKuut3iigvadJe3K75huZTgKQfjbjJqWSq2EPTY/soW6e+eQTBIYCjNrHtYVbqWMPezHh7SJox0
XmzQnP9ST8c+stAAtqKN5JIEub1UvZrYbHZADwOd9ukuyZZzuQtZt9xr+XAWaxtzpAQukAopNaJU
AyhKYsRv5tLQR67OojxljYbH708mZqfycQ+ya9g0RicVRqGl1W5x15akdhi8mRKZoeFXusI6RbV0
b12FyRiXGtq1CT7TOuGwJz5Y9gZoDs61RyhvrpyvXwy/hzP9xbE+k7AEoLe4BmT5sLivBcPTzmb8
lzCLNP7eYX5ybF8vLSz18n3gnyRJN8WfozmOMoz+7G5UnX3EtidmIflDE5/07gRlIUU1bcgLIgaQ
1A3TUB39SftQmmTZb0orUj7JNT3oIIgpXRSr9zva8mcXcZJejLZggOWkZGwwc3Nv+TM4rXeVHZ5C
WiwUNx1b0PMbKafq9JvWatbkGBuBp9qlgXjBZcYeFDGkWiz/MhtdgKc3+e7Pltj/szFzmWdTSI71
oKi/C/X5MdHwn2Gqycg1/EbvBQ7ovUW0JR54CbPWszS3cSWR8I2x1tXmp2/uAjcDgUqOCTiFS3Vy
wrdm2dgECngDyDJrQPOg4PsLls4NLWowcVwZLIKnPd1Kq8O8wupRgD3Zd7uvr2CCcXyVnaIZn01W
lkBisoTOdnZnL8aK03xrMj2CEY1OZrcgg9VDuXTJvIr5ye1onarpFC8nhvcG3TTjAeIcVQ/VOwTq
A2876V1/OayZlmL2z3iGf7ockTt9LNZm4nFc4EXS8IOloz0LlpTy67aZtsNkSr8G/JdQGWtNIGdp
fDYR/SemsNDPLqXDGh2QSFZ3QAqn0s37NK/ivtd7KuygqX1bi/GzfG58w6pdUOHJBmZlXNWC1VUl
zMS/gd8Zw7RmC2xNO3uQfEV4r3u9oSPbxFV041mvi/rZFP5RY2IsTkoAp4ZF6+psXZvkX3xIsBUz
M/knzbLvMevFQdVRIDpgLgRPLGAaJEBQxfko1UhwXPqdqQU9sntc4yfVjRenApNJAmqYt9evp+3z
uIr0a/yZtjFW/JF37xBiNp9M5L6r/bKoYa2HBg9ttrWNWcMGddcRp7ATljI0TXiGrdRDF/UOgQfw
nm5b15KoWLcO+ZJSYdNyigiB5nUAje2sijh1vL+qou7mZkkIJLfXwevAwHWemsKLy6Sx9b5chAk5
f59K1KluvTjQuLsur8SSltchM+Qigu5IhuhUlP3boZ3/RnzARGU0gL0jml1YmbnQT2vr8p4tOxDp
qECB1q7yn1NtIrlETJ5Gd0tY5+6c/3M24mZBq9HXIsPF+fVDtYvfNZBalHajNJmQzIaaAwDR0CFN
h7GpdSF+PJB5Z2ya/Q6z5M8iKCb0I5m1TaZ11KSVUAC7UkGdqrpN55wZUVWQq7qDWjwrWtGu91GU
oCFCRn8U/AH4bMWH7rvvayj9whW3yyqwi7eFWKDBtiFy0COhreZmL7uB0VHgn3qNVHo5uC+v1eex
yTY9HvIJz/Pihw1RJ2c/zQSEwqSkx9p0qQgzAE6RqjLSQx4LtykJXv+EC8+HsnFkVjYVprrms/al
ezN4rkiWd6s12+woMcdtVnPh72Z/hAPHW5mNDp9MCzkA6WKzLgOGdOuAG5Hu7juF9IjKXA8pg00/
WBg9BYrlbeH0WxYlISrRUJW16nLEC/9cKZKw4JLkLteiM3/AsAFroh0nqp12pbNls4CBq1Pat4ba
sEQ+BsumgV9442WNXiWEHnNjwyfMjBFNV1ylB8S6JnaJBlDa05eJ382C/8agymtB/dDe7Ztw/SJc
dgvv/Em5KRBfTHNi/w0Wn1o5GLVNmdEQ7X8EwPeBKUTBpU/TOA5bow+iFO4vM4ZEfdFfS6OiLnTh
KvKxnA1n1rJ98USP/n7i+VhIa+2/MJBPLLcFV6QUCZMKt7aItry462bTIK4FFAwXI9MkqlisJSDq
coaOLUNOltik0+/uEXSzJIHef1ssLq/e/m+RCFLl+ZBd5pXcgxB+aoC+IMzY85+vS16AmBdMHeIv
PIBAocvwK2KrB0qvcKMmXVkm5YsOwVhFyzSihr/2529CI0QYTA0J1Qq3Q9M/NUm6Ann03yOGejVH
WwgGqnKiqdubY3JCr823VidZI4secCEhHYbg9qkgeBkxp7DpYZ49rf3qKRgOYRXFTYJFUyb3gJCn
lYESLGRMHs71zUpGdLLD9JogT7H/2FDCaGb1fnZKHo0/mVsXv1NqE5cH0OxVrxosoNmat48M5vJC
IBHkSbhkWAP06aW7PkYHFaIUZWqUKc3A7f7KJv7GJ+tLRLjY449lL2igkWzDhZCTOGs1On5SEU7g
L3OyhRXRrXZmbzsF3ttbI22Vo2mUqg5QfqldOIlxkSBxZuOQkLxEP1GJBCB63e3zKQ0iUNlR+yj5
SHWA4lD5YvL5OzNy/bF3bNQjOTQmtZO21UiCGqwChkbLY1XarPbZYRR+zGisJ3lG5ibPFR0o58Mr
OzRqaJlbe9BrWiRtgLd7u/UF2eXi725TsT9Cak7oJ0dISeFzBE7pAKJDuniPrmzxVex+xf3VhCuE
Vs11Y024aO06EOCV9CPnXPpNw//3IxVi7F7P3x8khWYIMnQlWzoQJICOnc8KmgHgK642KO/p3COw
tUIP5jV0chntx/MGpkTF0DcPVWPdF+1GQn718TBoWJ+sbGSj4iLBMPl3x3DDh+5MjHURHiV2Gccw
cxwg1/TNjyJlfiag3VkbvM2hluFIZr7ijtzM6QP1dpP4BPSdzMMkvvd54iEJ/Ig81gm8/vsemZMT
MkaJggfwa47ipCxuUjvBOFZUpOi6N99dCCRYDxKO0nUEdrT+M7rqERGLemlpEQcz0ohGFsnkV1Pf
03svk/7wyNiyGJ5ZkAMKSXapYvmomnR6GUyP1lCe2ArCw7ORVgN4TWio5HRkPUnC1/RlEqIQPcoQ
YLZrSoj0LItk2abKTnOzX50rANbZZ8cbmGVUsDTtuya/bowpoSAInzi4HBMho4SS3YIn+hYfQoMo
v3sztcX+4VTCDVq74HmUKXmUvoLVe7Su/WUtbYjsOC9boXBjeoKrcL+FtS3Uf5WtUocsIeFOXPtP
SsNlaL7xFO+bQJfIyB1I2i1/OShYcDmp1zBeJSciUmHgSDv9JkzHZxfVri5St5OCTlb6K4aocI7b
/IcldBlxcgFHnVTZ15adkcrbMlxY6m4I99X/wLKRG8bZC+QNq5tzQrtQfYQx0TNOxqkf1X77SNIg
eY8mONyJv/sdOiLBrr1jEiX1XOfuDpZ9c2dvOdrj07g3D2dOjBF+e0ColOyt2UL8qKCAMb25vnGs
Wu43wSmRSClgE2l8pU8ab4Lc8m7mPuuT3Qto2buxDC3WmdkZjHPtCGE6a/h7T2X5sHq5zk2wbqnb
lwD9tZGOYuVk1HReLGLXUaZTgfhdqofNx6OnaC9GGvjpdxEbHUZ2JPxR+4aezQzji9qJpyBaO8OY
9vKkWJYjKUMRI0M/yeVONxHAP6LKHW11EQp3gcDJE8Y+6tGmWr9rJedXtYUI1MwzbMgSxLrRdnKx
gZWlKzaTe2ee9whuOESUzggK6997StLgkFwSpuHaSedRE8io/HkdSTDG+SCzMrGstNZclNsto5h2
h4VvXr2CvIFKoPDuCcWABMgZgbzyypExu5McLpjAPZ8zxNY/DBPcYviYzKkluAFIiJT/eRs+92mj
w6QvZLcS/gYfBZE2B8G8yFR1kPcFlUl7YCQJWr2GGb/oPpbwcI6OOjeYKWZXE+WIcCvbF5pNvej+
jUOdLhZsRKgr5IMnWcvkGU6Vvco5mV3l+MLI4m57OarpsLpBwz3pRDqjm3vxA6CqFt9tKHAjP9oT
WeEM3pJ3/bphvvJY6IGmiAKegs/Ji6cnTlgEuCjGYKssov+FusupSozqVM8O/9QoBxC0/emen+PN
K9i1oj69dYA/ua7bUb86CbFhRS/RFQyqyFdWoPL2Eo0e6M3mEVw1Qes3tmlyBPUastQj1pBjN7rk
lemsnqUD4ndzkNeixw5UkMAQ9Tn3VaAulod8UaL5PqJaIzcY9BZ3XDcYKKZv59zKDe3tPGIJXs44
iNXNR6eS3jOdzqRgcu2wrIFygmlr9bKRLc+HDw0yeookTiaRipQfB5Fve4q8Ol4KS4LEhY4Lpk7a
9wZPgtmrJvKK23gQB9pLNO5/N9I4PE+pxS8SV/f1xr84APFXfJ/ugdtJSoyVTlVqv8iMhhA2R99v
juXdAerJxTHW7Og25BYAeNF3KHIA8cEVUXWjfsQ2spwJylTCwJjpjQbbCoXVSyyM8ffWicLwDsnU
FrWnUn1O1TdYn2HA4exHJpHFl+FkGT/m9HSwJ7QPybHuGdQeDqhrQa77rm/ax7t6T2urQ0dAzNQ2
jUEIEwFcwphpGEXxaleXmErcQP2KtC3y+hHAIkDYHboR/FIkjA8433bLkaryA9oIyYYzSaL4LhKR
pS5miaJLo/i5QotnxEhOTh1Ts5FjzvjNk2QUSkDygcl1RWv6nDCi6p+6YB7xaKalJPLy+u/kL981
9adCEaJckv+KZgvcSRGmmjhl4FyvyMnuMZXAOCQvZwxE/hhgwRlP5ANJKxxcMsN7taM+3M8Pb4YN
9ikBX7NXP4uPenOHg5DaD4NzwI5jf68NvRe6czIYEqpYCGgGX5zK86rom3o15fTLf+MHdNzSk/Ws
lHSsEsRMlZM1ko8lpmL6jd5HhSSCjRKGmnHZcpiyGnu1T08qHw8w8fPO6qRa6jXN0tq2iVOp7T7p
yTwn9EKzvGmu+NRm3EwMGkBkMjCvIxbYn5/HDHQxwATI0oflvNp7scdcfv9DA19+pb3G9KgS0+cm
wXyenlSJmxHmGM1SPZMjsZITXQ4Xgo8xyRvtMqxQtgtWq5UxKS9c2yxwfpT1+qqX/m4IAKLBg1Uy
1O1q9GyYN4CIKuNzkW9rgPUPvMwp0eWh7ITk+e8GflqwaioKnBS1RNOyS1H6RBYJULJ74pHIOUBy
JHFrdftB0cZH8lac35zgVq/Ci4VKq887Jmtzm2dco/Z12Sn0WHAPXXXczfm5L6nitgyKXrByXZEj
xpNLqNsnYzogF3m9mq5G1oxqSL1cD4xngwCMUPd4KI/nWsNDDr1Am5qAMf1W6oGJ3flx0F4r4xlR
JG+hB2XEOD8gTuTRS5EHSUcryG5HjSdW4GeMKR7ZSQd8JT6H9liwC49ZTaLasOZNoVfNR6EVyaV9
d+tA2hmUCUf1mznjWphMIbfez1eWZZr7A/0ybZE+1+3qHT19OIUwFv6l6J9ZA03BIxrkuwX1dCYh
Kgdm28RtJ2ajWYihvmES9Rl0qfqFnxCjVkFx+U8q/wH0MwiU0fq4zTGzJZIfH27giCEOqyO7Tj82
MVt7QqDHNTtnMHi5A7mwB9TDRo7PaAwSu/L0qK+sisvYjh0b/QzO2vO4wO7WuydKXxzEU+ylABwY
OdGhtglYFVERz/p8JF3467hl3OKxgwfMyDI/h/Sc+Bg3uWawvKKLuY83SdCneH3ubHPj9WJ5SZop
bSQH9pyjOPFV1qPC00b/vjSkTpnClkZ8yrKq5nUth89KqqiRQwnn6qxYgOEif46PF+HEwnHTUbQU
28eaSTVz21zwGFhIWmILQN9kU3M1/Vr+hukhNHHUZI8FhR6C/H19ObG2yeOjkfGblJoSUxMFsCVR
xsJK5kjd/DdeOHPDv8HaHn50R0Fq4pDgwONVOBDSysHOX4NtDJ6wDdqMcf61J0eXR35O9EhNQLNn
mCJqdOc697avlEae2dXH6fzXr1CbRIiMHQMgM9/eptwCj5X0323leSqu6XeWfKhLaZUfw8Q9kzEv
/EYxPiDCSbn8K9taDylM3cLKiy6O7Jsk9JedyBqYAubrO9lRd8gmJF7orTguOgUlQi+WmMi+LLaJ
y5OG4xAwWgrEIpK9N+CCQYd+0kDqiSG1wgYp3SJeHzig5POjWY6tZE76UTfw10KU2gu6EDebtsDR
Yt6q9cLi0Ks7q4Tl+gtUkm5zDVthIU7vzA5ipI4m+rzkDeILpUiacer1bD6ypKuIjSmSedP/Ygqg
2jNqNaPySK+KsrYIpoaLUE4/IhmF/GnQ493LFTa3KMtzj4Bgwk4l5XeCh2pUyttqPkXmYmV79dhm
W2wlOJs6vQW7xfT7GbVpAtshKhvlDut5oBpF/FSvYQqbOb59UXZEsKiK9M5XnqvdJDoTtoLKrU8k
WKDLr/nTUaLDCGpbLoM1+jn2FDERzOatLx032JWmEHbepAeTIsAbDzmFC7XmPy4NVC7dOnJa8LUG
xlqc6QYwbVm+ahW9AOe75Wejq3RTjMh2N22CyMX+DOU1byo9L0/i0PpDglZimhXJLu4tnAJJSRw6
WpMVUmw7hPnG9FzZr0vECdtB0pneZQI9iJu4W6PyVptel4wC2wiu6mKllK7S9sAlVMgsC5P0Ro0b
2ihz2p98EGA8F5lORO8Q57V6SzaEzlyNzfq2oEoHCq6L/LT1vBu4HYuNCuXCTloM7LiWJ7kN2wbU
wNxRj59CtR6Lw4Lox+H0VEtqnrS7/YXE9xqaWwUwnDTVOs2oypVGHf1LD/56tzydSmKnS0VLtmYI
HAPZN3cbsC4m/CXJuWhoqbkmxyNPqmROdd311G1WBAxC8G6t/Q2W9u8eT2xOSjiAqBkNTU7h9UeU
thpVDu5XBXjAP31kPAkztvbpdl6ZugRk4GVIVH8gwI7zQtyqdieFJHNlVbxOcxFIxhLKjDbAle+G
9x31P35grh5p3AVDMUEwwiBIJ9LRP156R9Q7pUy5q5g12ngvm/qwTQ0EVsjegt+lGmKhYXBHLlPV
LBe9J2FZD98XEPdYGQaHL3Tuy1AQ3vahIkYRItDSRVc1i2cSbwwZWx8J6RG4kvdWpayNNrNoooxK
xJ+a4ZoVmn9wgJgzb5jdQN9njoeAmSvA2DX6pSCcSPPTknHcCz/sfvHesQAe9oToEFnRgcS6nIcT
Bo84GEiIkv8lkyTXFW7LVkSPp+ZIRC8OiLJL7Yad0FNnOE9WNNZgADsz6NATUUzRSGTYaVuLbtnZ
IyKUBOfK33s0Pamo2esMUV1PqPkoB6O9pRaE997EEpqMCR3FOyeJPaTrUw+6P+ivoYj60QiTVK4F
ZTY6wE9yvqoL94uMYgVHrQhY0ur1KSTfLQ6mtf9W3rfBwx7TE3rA/Bbh64+LAbx63xqoDLmuNYef
R2wDMimV50Kk0PcI0Afp3ygNtgc+Ex3w6VO1R8rsG/LOmGSHLYZDspWFnAmR6En2Ou1OjdO90f32
O04jaaQvBmPzWAeAHRMEMBwlLXvoDhdMwAkrvbYCamVs9dSo1fi4XzQ5VuwVJFRz7WhTy/A9p7hN
cGtkO8xZtAKC5cd0ZdoY1r6P3E5R5+LcVI3oOd7xiikCyFbV+U/dj9VBPlmM7zovlSJ7sfeEkuj5
haKxw5Sy5mdWWLllRY5bRes3BO8dakPJlMDyxC+aYWddYq2MVKwDjVgOnNXbMqlW13iClhm5nIMT
GKwGAzoJbL8mKwujCtUg0CF5qCpggzVEtTwaNTvq283xjlrvbyYtX25rIS1JfmXJCzyaOuo1pqa/
1hei0E/84llHc3QiQ6UVFUEr2NBfc3oJSXP33OSyLKy/4nZ22TEWh+rou/nydjCh0ccoVgfYhXYI
Dk00xk3249xpD4wg/fy29DI2ey+pa50cgigGXoiApSiGqObdLkS7mUPFwy/LgFdf5oxCNau2/ij/
0l+XYhPRjqTDZpc9egOw01wegXxBZBez5d9uHFB6EmzfQMzi5oU/ypbewc0xpYGpsVNQeKbgypPu
SHPRcgrCmn0DZvFQ2fYAympOE+VNTmqdj6BKBbn/kaf/Tg/Z3xeHsHNJueB4uxGnL1baW99ap4oR
QUvfUwW6+c0HxGJ8FVhdRNgnhyH/m2U1+mRVw/O0NMTTqc1knPbruD/R1uJZFOy/pgS0LzbJS62S
h+lqhHrwvTFHqidso1AUp0ZICSCYWm3mBSIv5Pa3WRGxbwEeZhoYPjR4gwvoV1+P9vyg3rxT/7r9
r2CFHon7jo8MKdo6MeaWI1ZQE/FkICJ+CT9pDwgOAhnoKIjcm9NEC+8s2urrWmO/PKY/TVyMFdnX
2wIjtNp14Odp97RVgAlEczAN0QcNSMmAWzhFdZb13tyucWj71lF3w65jXIQbZV+9XaHYHlFx7gsY
Rsq51mdLSbxqMz5LOIIXXY801maxOaR65BvI0QLcBocyCAwOVsQierhIFYYGarBOc8xErE6bclvN
aCAvxUsXTNuAmjh+ivGEqtsGfPOjYgIYhYG55PFmPujDwTS74OvmIsiOSWLsPtv7EtZj00EB2Yl+
59yC5cwHITcXgKhM7lQO/OsAiTTSLjRPYNUncMNvRIMp0A8CzAKjJ4cgajr94VhVTIixyjs01170
9CLtveXvAD12LZNVzkOh/uAf18slasOB9dRp8Xd4iY1mXaya6wyrsMpfqbqVirCMUh1hGmGufb2u
np7hEEx2AhYtVAZS2hIFAhdUfbTgiOcP+WwNUTn6scRDxOb0+fhFwE5BcKXaet+R+AKMWke/ET0B
gwK46sJzs4/Yk7I4bVNsLBAF/1hs52jlOLXQxLuw7j97dZcs8CjtHb1j3KpKpEe3QOPNFSEKDWcq
QIf4+TlSiy/U6iirY5B9+BJ5G2Fx3fC7WlBT/2yos+Ouj2tJomAKATUPmfXm0hnJLMXol9IfUXI9
dFXGrZgXWMoFsMo0I8oz3c1C4pACyOGyZjlrOxyAjeAVClWiWG/i2vxD5khDZjvKv3Y9+ZiXheOz
bUxXzZUdkLjoSPs1HmyITqEhCp/86eddpv6sKSB9ZvEQSa/3Xvc+RROiz0GwvnWOw0Kk+zsb3Zq8
NZVhIyiqvCPaJ3urLN+2s9HV/Qcjln2ltdxK5OMWyTjgN2ZbjWL+MQcvc+WMRXg36IJtiRuX3VWt
SvQNRAgAlrpoBJ+ZNV7beOaXkNnDh5HTQLGz/tDAsTi5QjZwgNHxcVmJeq+DGFmsbwyclktnP4eY
fDyK0TALkZPlAu4G3kAWJztxofgQrcYMdAgUn8qwtRBoozlMG6eQ1Q3DnjaDETpWtyrEybqQpr2y
v4LzKsU88r/2ebhwyAOQ+VhXULpJoDzj1etYX7MNnuHy0CLAl9CuvMNBzwoZADiZA82YKnQ2Iz5+
ElaLNZ4zJsuRaRbq3Rp0EMK48d1zzx5Ku7cunwkPcezP7O4lOd+0JBa7m06aOueWTgMH83P+oRku
PRxaINnmgaFla6wh6zt14rn6nVF+CDkdLA/boKE4Mh1B4/sYx82awD5kDgQwFBjIEv1TiYEi6S0P
sS2srHvg1AxfwcIs5kzuZn8kZ3tfYWhR/PAs3k3YrL8zReDqr0ioQUPvXdxGMwhNfq3C83c5PAQF
sMLs2o5jIRPrOPOSzQpAGffc1oLVbzJAgBd/ImOK46smSv39NQRQgeke9ufULiasJYUc29s2ZTc+
aYWeBS+DiW2JBH2RUIhNSsCyobxshslRfJ/6Ag7DsrDoLpsLgEY4k2EvOmY11lKpQgz7KoeC7HJW
Q/SaCIuwAxo0qRrXyWIEiWMiY7Kz1kFotMQjCcxk17ARtpeTR+qrPyoWzZ/Qx3o63Fl3i6OjHKOQ
uDIh3r2JGPIgskx0DnjTbsJaJ1syfyOUjAhgxuKyrNfguCJ+Nfw63XuJTe3KB7a0ODQriJAbEjvp
g+U7i8bI0AhLK0gy5z+6qK8xVglSCdJpcVv1TuUJ2eeDPZMl5Bc1i087zuGDHIzJpKz09xeHzLcz
7gz0jpwbDvL5Gtu8/aUI4G3KDUP6c+M0oTZjaaIIqS1Ad6c6h4z164Q6s/fkL0/b/htl+vOz3wdC
VCG+r1Ws2rcNrxl2YjC6080IVkCCcSngF/F/nRjQ6KsLSAB8lFTCkKGKJmjYrfIsHf3PbjviSSZc
4gadBU5HVhBUnILWIyeMo5QTZFnauEvSukxXeIJCTnIssYuMjx9M0VR5pf48UFpGPaaQyUPLuenK
/00t7Iw7Uqq41YNjar/WWXIOUc+x6a0Ik9yU21oF9lKjPU3u2pyPQoOffWxutnlGkI43EAr9QkDx
CMzqbOGhxhijfz7ftzRXL99OZHEMqVv/Res5i2CeHBWtJ7P4kE/NlU+hXZfL4sortdNEv2sRI51Z
zw2tYq01ttqLeDW+pLojmGy41nyy1UmbWqLNgp5LoZ5jmOOf9bsvFyaLDMBxI17tGZLkNXxUux2Q
jPOt4ZKHLhlhA1RiBmRA9yR+NsshnSfMqP7htPwhUC+fM8UD7pnw/2BCbLaqeR4XPhuEqYPGJDYi
Uukx2mSJVaCahDs+d0V65EBri2wLwELBn7bPFoMxSMf5Lv5WKf7vbWh453sQQTF98jF9uh60ih0x
5IDE8fepOyWCsv6byPK4X/yW02fRIuDy89HUmInxyzmkyqtyX+uLhQnrM4uRUu1b39kqn4th4uXZ
1SgKeOAJ/Zp2ILdp8SntL1yzTHIUCblCa20Cw9/eR621h4neu88VGQc5QHxPTuaq4gFUnf7aBwjl
RnYPirDpRJwmTTZbv9SCL4ddfFm9DcrdeS+Rg6aUoaRvtc9EUqTyFL9vg7pohOjxKlkjqrT6hxRR
xv6XuIZVU59mwlfiNt1ZlchieffL9I4mdfwtBP4ADGFd3RjSDfB8R1smCPGX16vy4Dh//utQ6Qxc
bV6kgwuKA1wc6+qsbwtEHoBBbk5mATIt1l5Xa9WzJjPGJILZ4KQhvvyilyAqO0qN+ZmEnHVtM+kd
na02JCZA6oL4nrpJ0ZUBR0hmKrLwjIm9Qe2AQLXaKlDtL5SRGGIdFyKGWAsSct9Q8uij4tzpa1o2
uTVmZDLtccHh9KXTJrnzOq7X3qBjkFb1r4VjSTM6e4sFM74u0m0wWw7o41BQdKjibd0y+7DPcRY9
4y0+Q1D4ti1YkCCUJX9EWTAbr7RdvUee8RyzqxS5Pf0JuDYJl2GrBCLQnC+uqIejzsoiXmfjVlz0
2MAnt4c0dDlNye+Ow+mcSZV+PStT4HaohG54g+erbXk6lawSRcsTPJULk2IWNDvopojlwWrRFUNL
PEGwVLyjQ2akbkcFJpvxxBgbdTQZ5MUhIMzvHQgksxIvOoOFY+1W/uvHHiTvHL/lvmkD4WaneihU
YQruLJ1C0NQ5E2ew/BlPHp0g4r79P/Y/gs+3Gpvetu9QMQ1oJNFH0zvvBqadm88vb5YXaHuyVZEq
gLPePtmi1865pcL/m6l43AqnhNx+i3vY3jq8sO3X3GK5i7roNP8VJDV8UnLNTNL0se6TWCZU4Nui
vi7VKnVDF7l4TDHmZL2MIs4+J/Whf5LHkOBzqfWocBUvICgTrwtPii8v4JjVsfZ2+ZmcKMvaYi7U
jmz4BTkgUoTdcWBRaLRLOxHGOZ2IGr5Wf1/Lbnby3UJQt5biNcoi4YkyVZlGNWR17BL/CM3RxKv2
kZY8pTpstg/+siA1h/Lefzw2IPyfYPqlXH8DMK7gpIZjVDH+XiJEYRIppdlueTZPTe/DKcXw/L9/
hDsaPTaLGuT1ljFMj5/Hr6F4I3d295LcAW+qOGeKk65MvQWa4OvNj3hI/9D3KArFvzECKad/8lls
EdAKuHA+CJ31EJrWILNptwB7IGldXs4V+ZMeAIShLxQjF3P49Z2tflKBgLotN3ahzpIlMYyujjJQ
VE32Sl6HAozpxct21B7SCLOSXka1e96fZdVvvcSL+OrUTQAcPsWivQ2cy+ZLjzxyIgwSS32VZonp
Cf9OVCWD1Z0UjD2u/7AHg5NAom7vRBdEZnJ1o7+EffoGM3GKI1LKmjyr8eQkNaUbhrp4vPwvkuJJ
eaLmDTPr4UmkpfaUcPox10Al0mPeFkKu4KyjVUy3wmjQwb9rhYCtdgr3NJzL3SESVPuMeFJ77tz8
+ByauMHLz2M0T7nt/yzqftCrtj8jdNSoIC1c4L2yfKnRtxXdPA/39VMQj0TD8RznaZAfyZYqgsIh
/0qPyOcmhLtMTF8xZL3SBp8e4eE7yVI1zeBiQC67llKvofNZSBkIBJAGVuJFti0/wfsFhaCUn4FD
pp+f83ms3abG4LwNGc+CjTz/slb6Lias3h94Zia35MyEK+DK0VB6+DnmF7A1TXHZLMa/1/PgkSFS
R3r0OwDDMdK0m77QXw8B1ftccCb/APPjzgq+iHlQPPYD0+9ByTRVmUvzHnqLLhujt4LvRDDM30JU
hpOWo4wyc7wB0U771SLm6Xs7UX9OMDsjVMT2ZPO+t3Rno7zPn8Eo0wV6ioXnL2HA1mgEoNiBcOus
NPhi2+AkyYXxMbxUPuuO85wzPrfXF5SRQmf/Xo+dsV9PskKrQyNjPJ6wVfIrqmphV3owF6SBybob
8GEBMVP1QtFChB+HPj70++kdsH8cPAB1Lx3SAGdaxb2h40q+rB249dZYiGq6RJLy2hpG7L13bzM5
PP4rvxm8AqTLfsCIqB9UimcJy46MokLSMz8B5B5xUfr5PlkSL1UcEUWQKCTOCdeU7vLTJU41lr/c
GbESQbJS+lvcykdVox2Q5fl84TaUKPqGv/T85SjJwQdHDAtT5Iv7pkKFtz6N9C1EG6b7SVU/yArL
rCQzk6LgYH5UBTRaChz69jUnNAMQ6E3yYa22aVz1L9jljTL0pF6x41v8QPuJLCh8av6+hRxR5sAW
eptus8WITDPrv2qi86dXJxxXPI8fL27dNF0oI3dJWinnve6kfvweMw6g1HM4tGxtFRcxldc8Nf9w
25SgsEzjpojChKM4H/pOVzDiN2zKXIAT2lYeDqr+DZHrkXlkFJpSHN3EdpsXNPKN7HsfwqjRq7CT
Nb46GyLf55hC6ptkFWZ5OHP0njbW3WMmwyOXMGZOvG03e27fDyQIiGBg/3HeHM+UgYuj3U4DHcZq
lkCTdBO3YYtzckgmc45Tojy0I2NNQ0nYbOq34HYUP4YzOy0BPLIY2rhhu8xlh5a6hLRqi1F/JX5b
TysN/Iln9z8ZRZ6iqMz0lrRr+uAAdgCGK8kslOBmvtMOzMNjz5dcq5FKljQoFfJf2kdmAuwU9cr3
vrQAuWdHVuTOHQcgrkc/bb1Ol5999t+lbjmB8Mpv2W1ItM5tmYGZAwydc5dByVZu7J0a6bWzJHdJ
LTEMD8yugACrrUXIHURjdusaDh24086YSFAmzFZNfmjyVctOWqp9xePekhCImk41kcrMlvl38Wuw
SqYdeVRaa9JX7jbd8C7AzgCQPQMOKv1IOfp0A/zcgJzB/ye4Is4zM9FY+zyuVRc/9DT6TfSzy6XP
ozwfMrKGEz3VIVEVE5ejvD8eQ4RpdD5P3B0BSCRP2PUldsAtRn5yGYZa8RTJ4tEGyrbgA2RJLKZm
F2OJdkMmHewDPN8hxGLzv9PWqKWAFb9MckUzUr9c0/wpqKTbKk6rrNW75lV20ycijqp4mReHpnUZ
DUq8yAEL/CUAZS25eRyn+YJmpDRMGWpUWMeCbZdL1FvsEeUnsH2TZpk84JtFn//PrQlR4TjuEEXY
56OSBDBFUisotAmx1ih13p4Sr+rswTpg8BuoNCnHFr/SzRuJPALMirGj+wS8o8cMRYdf5Fewqape
mBy7V9hXRgKLmLjBRhei338OoVjBjeOQ92qYbBI5SQAcD/S3UgxkX6sbkY4URQCiXn5MxX211u1w
Y2QtrXHDvnV2Q44cL6XV2EV0Rmfu2YUTqRxkdTHGnAS42665T4tOGEcbXFINoLXv6GTZIgY6crx7
kq6FGGMb27spXp7L6JiQBvYzwy3+ZQcirV7V36IHiNjCCyAZmoHntE0QBPznUiEu9BUewKCvwY2p
0YZNRi2b36yAJDH4Uqg6Dv9vZen/sJyDZakrqUgoGxb+Bk+LKAqHAhhW/Z7EcKG06pC2EXpXSq0B
lyT++zhEVOpEbbkQWnDD9sv73ryNfE6QCfRtgxHBH2azPDYWeYKfSTFQijVj6f6sORow+35RsHZS
NvBrFG9AUhaixULpqzWcmUT3SAytFdS/8+69k0Sjng2CyJ6ECKSKad1y2pHdVmpXqR50r0R3sG50
t/W6/Z0vFdajt7wdwlRBo7uTv4vf/RQ925l2O72xvICqCppKaMhoGNsP6h2QUJmHQvSeC1HHq6wv
tdwaAveAl7Nl2lYceMb5WQVB/Zmr1gcKtCD9qi+JGNj5zQ6DoWThpWW5uDkvmRc9jNOq+ghqzoVr
pu31/iATHqSVMT7jmVPLfnHoc7h3vrG7zctryFyG0wZNswdc6GT2gwTgSt2XLSxQs1R95+RtfuoB
T7ZNS3GxIcr/aAkMKH0Hq41sk2spbV/Molqji+nyk06ekyHPts6Rai0qpKVJbsbYrFolnaltWj7P
2MUbciEQayRKvJqXWYteqP1AvtRKXd9LnMTDFSBev93lx+uZupp0qSjsuvXtjSh5MAuQzMDf1bA1
HazAR4Izy/GufS274tV6LWofjJJpL4GNUhz/wjJaZeb/zdsM8oTgfugD7wiPoMFLvSaRQ1PTJnZ2
bcaS66dwyg8Br3YJiG7JGSHJwF49uUZX1KoulBPrDl7lYBcMQQhZqWnZjXHauxmOLYzGZJB6dlAz
wfOnsfF+l//VvV7QjVmJe5i8lBSwtpN/PuMC6fLygvjK9+oQFRtqesXhXvZh9RYj6gPfEmCVTbBi
aCINR3dtpESw+FndgDVJj3ZNthXVzm8npYGJFlbu4LZoDOCFwHVeOMnqkpjTFpSGqDMdQVUzfUZs
pNljnKamdTQiDDpNy2p9ip/Qeg8EbVnT9aMWQvhHbDBuRt+96KELIkCN3RGuoLbxW5p0wnMe7rWU
WderoDcCep1tBVcKURYg2d3kwqhe8OXAkz0GT2Axfug2re79cEvkQbX1MjxBtbAH3maCbYUIWaKN
/AbUAaZHrcoh/ZFFEF9bpC77/FJMI+8EHtqGh3ahU7MQRGixa/JdX49V8M9MaVPsPrBSKQwV8GpS
ma2oRDLSL6ccf7Qi6oJZaoY5HH5Klckhw86ZnoQJuuaIU2TSP/n69cQoY3LJBdgTw4frZsWh0L9m
xMB1s0hoN55ndeYB3FnwDlqbfiKyfNBU2mShuW9gwUQZyVhZ6OHaczBToj6TwUS3fgte4YJqaZmr
ja16pnqyNrd0M3T4rsdAvakuXUbEDRpPnMY8wjHLIVY+RkqRCQn/6seQgbTqVIYZ3As8fXfCrOjA
BIsWCa7WQ7vuzUdBlCbafIGAn6ycgDXXnaIdzdxa+GqskPXO+eyCs4kfxNt6ph5NL193vQP3cLFd
wnsF5Nv0zAXS/+2hls1rXvhUNjp2G5jdu6aT7Tf/DykxYpXsH26ReKckfsXN2n0lELSNDVmmW+hp
QseAHtYItvARECOyp1tgPNFMErhd4k3HnFO7Nd/FeyG6gWzCXP+us7Ao6ROKq+JGdjYgUYOnVlwy
dP749rwfcWMKrfaJ6QqWSun3yeGGmySS2ZASiBvcJTxrEUei4zDE8dYRRMkWNK/LPIEi9/VLTKGD
aUfQ5VKBeg4MrxTfFZdwpaedYBCDGu6TzTxJKPobBr/RyLke5V5BJnb9CqLgAuy5CALa4M0oRg8r
M5gaoNXEtZwzFlEG1lb/HuKCsyx2Fj4ZPSh9r/ibzMa9syFEXq3VNtWgwJT8uQoCcT+KFUNV2sOI
NVjmJOL9NkuuPSbQJYZAGmN3HU669Lf6rqegxSoYilrDf5NeSiA037ZMHIqkpsmLOmbnEkrvfu2w
inNIGy1Apfhgfo/4GhmsHoajyCUXRvwQVV/92+mDANPA+JqHQnc2T4A7USdUmZs1lPMeRAt6C+XL
p/ZsqK/LDHDtZRHsNPoEab9iRGTTALpUaEVML8XwjVj7ytTZ2dqYW/V/h7AY0ASOafCfYksOgokn
jhkR+LfzMYqTiczBw3W6vevc0upYfg5ys31kLbOj3pKY8LRl1QrLHA23zIsVMVvyJ+OKWRzEpL/x
oeKzX262w7OVYN+74OEJecr2uDSqF0RFbn8pd2EeiWqwaPL1ITuNyjU5u/x90XwxotcoOwEaPPK3
uehkyMIzF5Livyf+VFysHDSsCcgqPdG3gtHCM8dfFry6syDjmg65icTxrW8lt2RAXW4h0oX81OwN
HsU1MPUuESAxqOEZveAaWihnG/2wHcJNokhvsjj8dXthX6wE62L2jJaaq5tWUpTsTBeyAGFS/pPI
hMF+UpOXQ2n/vxZQdzc4YzYelAL18gqEwppKvQy0SeQs/TEH9IvpL+ikrQXQrCMD0toSuNbkYiWp
SzdcukF3OVEXqPmpyRDpZi78PkPIop8KynK3Z53C5HAHyiMGBniRgPpBqTQ9I3co8xQ+UnNp7Q9z
PXDJQ3MlKh+BJaqZTL7ShtbjXJjaQq6etU34+ZCEodrxHDsNgCmS1nHi/f+GhZU6ePF+urLHCbab
fuyluTsXMXI+4+mT8POP9ZfGdiyG2yTYzrlHPi9dqZzvxGiLbh759c2s+aRtU1M2bqGIVRbOOPEX
4OYzEFx03C6vkrUN8MhEs7oK+ufME+kTdD+k7jhu1yYe98blLwblZ5ee08qcH8/ycvxiXmxYEB8L
ojj+6jaVE28UejL5pv+nbeiIWHxjmE2so7KNlTepF395opY4F9s0mM6TiCZeevO9PJlgD6rmqAta
PEJXxMpvavvPtFCNgHzqN977PdZj38gf8T/4sj/nfZzJGttTVqOYD3gAg5pnUgD7p3rDtoiLomVO
wBpd3o5ujADBCb9o8AJwsRRfcPVN1Q5hRcg7OzqtNLimO4LWlkLkhOQ+Ffk2RH1fjP8R3aje2dYa
AxJEp0+3WLIZII83M3Zf/syZeFNjVSVbqCQgtiBNf4umh7QNe9KKSMxLfTIoe2owHQbmlLyHXZJm
FqJtHBytgNHPfcgE14YOCrjWbZZEpGDavzAefDbj/mVkocKRQqwLqp9S8VaHx2H81QLQfPsJWNxA
WOIoqWH0gjAbHB5o81vUKxfXo41VfqcVuW4PewhoPsqfzRGfCMDNI14sptd4U3uYtD/uBK/AdZUE
03g1FgDxgberize/B1+ESwwsRg6OAl8MLFglQUKNrw0VGI6o1UKpoJD7st8u04s0EixZRgZfChOz
9I7P1o1b+jnc+aFMhn60AhKkabnF2w93OPDRFrB5Ygl1nz3+QjM23B0iQ4xZ4DCTpKtUq7owbOCz
uX7eGlAe9Ts+tUt9RVoN4XQn32E6ScvVeovBxYlPTV5vSs6vXlTuo2O3Pt1JizTUng7dykHwkZhA
bo2d4EOmHSEY98jRkvAisrgP15FlnbyXqXGNUuxERRY0ZZTFEfV7oz7cQZsDD0xcnz3fJZZGFjPg
8i03/6tuNoV/Yx9kEe5eNUtOc62AVt/rtLgoXyDJboqPfkXGBihGTI9Y6OFUOh0rOq9/pi2v5tv+
sTsXm0hWaI9oOkShwBmsNPbZynCcwDgb3WGxnOCCpmeKIRd8wCty5ZCikkGYrE7BLNDM72XhTCYg
VUNZc7qZLpdf6R6i1vhBflBBHnlHMdtO3WBppHrm6FtV82pp76dNYmTGaU2p0cd4TaEzSAYIDOQe
iHnJF6hggnS4awErBqykA1LoxpVLqJO9EIU5f7N1LnthV+XQZt0Kfflx6B9S6+fAqczi94AfcHeH
sGqyF6z2ne/57+cO177aMtuLuGoOi/CjPGkc9m75rMewSMmvJlBjaQDFj65b5MLxOPLe0mBAl5YO
np/+h6R1AHv7FHC0M93QdXGm1mqxtXVSBx4nBHdziPbXQR1QxrRUf4tvEujlv80m9Tv1OgY3YoqX
iNZW2OHb4Qc7S1CoXlvf0u5z18yk2XSRSvnHGXjABKqadkz2uZu7W+kTYnQulUaXdw1UfCmC17jA
t7GHl7BmTw3G2Z7Eqd4HgSYsL8BlSLhH49my4foNI+qRRgqwXzdRYFbmgCLSSJIXz3LWiXOif5NV
NtKYZ0dTaUdLaaqubvUR+IZAVuceaNQjSVHvxTzUa3xkCE42g5zoJxaG5JYEO52RAedsroJqAiBG
IU0pC+w9E50+blJJ0waGyZi+pSTfwPrAz8OiUDdLZWi1aIRIwSvPafsC18XwFrmFhiR7V87DapCS
XknTeJTrPU6mtf3PWmDsvr9JZdYtmYiK/9rVcUVlKT9w8reVYpM0TGvbvSVAMFMWAuzWX32lAe12
OrIQjJvz3HQOLDHb7IVT1pIi37h2L8ek5EV4vaDLXKjkr4YTsNDt4UL8BJaY1LMReqygvJaqZqRn
9qEqGU2auR/Aj8+iO9a339w+9IC1fZ5dy0NjcdgpQEKCywOaFz2DkVORkXuVTAA3S9z+I9ad8P3H
A8uBLf3cf8pSAjPUMbRU/UhzWY68KaS4MuWqpes9IBbcXT3cpJLT0rakDqcJc/iiMclWvQFSp3Yc
76CLM2D3yb7i2aJXSK2DzoPRfYtbL88w9+0JFod5EbDOmbmmfjFySMEZymyM3IaGd6G+159ZvKgV
QMDz55hGgpbwCeZPm40EPUE8OhzLwGxxeEOcqY5jbimrqGVjflql5DWGMukimt0hd0JIX1/riETF
O0ms/aZVIEPd/2bivQFPPWXai1/NST1WBnlP48w7p3w73SlQL1IiAKD/KWb1HPWC0TB34MHdGxlN
m3haK+W4IkW+fofQTUC1GwM49cTA8uIGqfWZylXltGPR9u4NC3tcRbzJ6nGdGkztj/V6FjypfJuz
BnttlFuejxEEb8DHPvDxQO8uatQGczNAmeS8MZ1nPKo7L7PAxVHw3n/IJVhRiI823luBSMwxoHJ0
tBl7hvBQk83uSwTPrUJFT+UJHTcjEOhbtbBQiv1fPBBzi/26wwOqp5U0SECJb2W3/Hu4iuRbQVN/
jRZbFL2pR+5osEJclGB4kZsbxWEUzjPd7TW10Sa69SJoVYneBuAzWDc1IbOxYNDzoG4Y9GoK+Iqs
3maMxsz80F3u/+j/LiUQFA75Bg9faeQvFSfyBVLr7ACcQFMeg0Ce5Ukw+5n3+RBSBs2oLFSCSJ9Q
kpCAThsGdHeku5iTXQI1lRwvshYZoNDDXHEL3gxy6NIwMwZz7DSJiZ9b9mkfB/EE6Kaei9tTsUis
UqWiQWXpw/C3ASeLLXRbfjesSIdICX92V8flyjcOglKFGoFHQKwjaMjMH9zfx62Urty2L96I6kkl
yJ+U9cx0tAYOVeuMTC5M0vvt+TP8C76hNgKieAXxOwg6f3TJquRVZuWevRyRvTDHcHOyYEl/bvv5
/vAwZ4slpQP+f5/Esh+7jNmVAhsW1BDGv9B/C3NG5q/9p3HaaqChK/WTbiGlPour6fXkB3pbnojo
uIoil2R97TRLOz55h/CvFqmos3cin07tXisNBa2a6DdPqm7XPFJtlluQ+XhwxWQmujPaz5V7nQD8
9hdo2PWC2XZvC1XfSL3ehwKJ5HN9Hqzu2rkZaCIGIOKtLEl88cg77TnsDgMfRHFuPv17xUbwR93j
/XTp+74subto/IFhTdx7VHu0UAW33NOxkllO/TjMAaPkt6aOy6pnLz9tkEWnX7lwR2JqncrHigFw
ddSPzc+H6i+u7yaIiOvmVlD5YTCvoBLQKphaghiYggW4OvlLqpne7a7jahTw6PQsX7qQG8Qqk0ow
8AyJQlzCZq0utbfz7bn8KX0HdC5zJ0m55PTfjHBsI8ZTZHDjbTDTyteSj6UB/6YDYIaiQMC8wzcs
my09Avy6Ysy+xW01tz4yd3haWawQdbVt42Qz8QZm4u63uhUSQXcDVJCYk+MjvFi7QKtRx6YK8J/B
+y3OlZtiwuO6vdEjoB0aR4Dbg9orF92JNSHjr3q+D3O6gVMZARPA9UuqjAIczM5VC7l0DQW9TXy5
9176PgjBsjFBIJhTAN1Vu4RLOfossaWVerTxJ5V1RJGmXC5RuLKbLL0uigzRASTc6CKpAmRvfRHM
lWfCSHgrGh7AYYmUaGcqY1Lj7nXZEZ/4OotW9clco318yEJjX42nR5lGC6LVbmAgMG1BW/4ZBeDu
NAjPop0XYovjuFK4Bv0T/OI9/CJyydXycdxlsUHM+5NwzDifYtdH0esbD7lHYLxSJ4VOTuhwPAB2
eVMXk8tEIZV7MwBsi3aORlht8Kj7zo1GBTujSC+JVg7/QLjxcZ4ejBZpZ/RjqWE7PF9VNCL5WUKP
UtKpCLee+zgm509/cyugfc9Bwly2fPGQw5SoV0d5XhVR8PSFyxn5cYvzwUb/S09hzt1NUkGr8UfV
TBmDNL5MQ29dQ4KjX9NJujh82fydrvjcpYhf1NC1M2mrfkHujwK38eO6ScPzRNY0/xJiS7JoWLwW
Jj1EzJNaOxlzXss9mmmR3GS3f2Otd+alaQjyRQEFpzFfUVZ9YQrBJIHTDBtoPQ+EfQye0cRr3QBA
DJLPAKaPJWDM2weHVY4908kC5qcBNx/A/AupKyGt/6f0GElKdu4Zi/86gmy0R+EtAdt961D+wttB
bv2b40Jx/xJa3JrEReudWyp5zzsF33KoC9GIGSwpXXyJRHQsbzX4HwnNaYaWVl91YVavUnMmXe0S
QMPoUSyz2DhR5kcOs1w91GXXgMduqIFhixZpvl2+AmgBDdiUR3uHdoPn3EXD/+f7viwGhvhotSmO
mzYS7d3AJF8R5Ok3DHcKksjiU7G8fJ4HC9bXrJhPqXSFDtgOSv9QyM0PjLUOwUjmGAZ8WwS6Ge9y
ErfUZzWw3VryRet0rWqPLmkh0IhZkmeWGrJZurZR7AD/2qgPJ8n3xkx9CVgQVHZmZ5lnHEVVq1jM
Ax8sHqkCPqS40Ys0WnQsC0nNuNp/FT+WvvZyNHfWGvKivHp4fiSqmBBywK2lbc8pPUtERuz4ULaa
D9SfttvBu55nizMumXlTJs/JL7Bp5GWDCUJ4rGK6zeiSbBOGxg1hSjc6xXkAFXVXmPG8Em+BRgut
peocuWDIi5LDuFjyYLwE7C3vzWGUGbxAyyrjFcccHt3xLI/DhBXfYQw8Vjdc4xBlrjiT0FxH22yZ
LQXHGNmNHHZ2fjdrqmE31MXXPb+VduPZmokF0ZRGwj+EjubAfUxaR++Wd5pm0NzCwpH2Kerx2PYg
k2z9QiQg5X0E+ccUHSfiIhu+1tY/pEngIe01iRQOAc4AxpAXFrB6kTbH8Wp7lmdz/A/IvYJee9f4
rSjiEa1TUEDfnSsaSpSMcYBFoHx+62Komn/hx6BWoXuN1c2+MGveCk/od7WQx93uUMe+K/9xExhA
09NJenvbKJ2EdESInU8RCDGBP6t0kKaKgnRlvtki5mb0S5CRzZQvD5pLpZLitQmaedrnr2dPdh6Y
bsx1YIywrMBDfnZCIIx0jpJfTcUhq0ED9oNnxGz3VvbQOZ9qo+iHEiZbjc80pHWljo+54U9gshZ/
PB+bteO3OujOiYxK+EsRisZXjNTONBxl2FZh2xveOxwXF+0U+zfypmmDrYcJx4Zdyr3q76kMg55U
SRvJeP8391p+QN/pvxGeLOfv9LCgvGQq5Er2sNWPujFQZd9fIXQywdR50PZlw3sG2prhnyR2k4Yh
aH38WOillalc97iUohBMKXJZN4Zm+UK+3kvZCpQeqcC5rSQbSoNeL2OgrJug2jLErS02Wtrk6ZX9
9w7gkooml0igktbwfwxrC6deSZFV0jS6G1j5fgIv5e3LF0ZaAFp1GeLxXesdahqVZzZ/GUrpxrR3
9sjj19GBvBtQP69EoQGg3p42tQLBP1Oo5atvAMRPVdvoF5uJ+NsWzaLqv0xzuKuNTg7uu8owN0Iq
8uDPAEaYw4GrB8+A/qntOdC1ypb1X6TvpZoXAkrqC64ECtfmzu2Rrte6hW9QXlHOwXsjzlGtU6gZ
f7+W9eMlHNnPlIDGFDa96qKeybVCJYv6WGDqIaWEA+RLN8fBj9gixgcWCC3GAbYP9KNu+wQXvhqe
wH2kGGuTW/UJR8umc/IMw1/yJVy2gnchqNSYDNcKiQ6LsGtpxmzHZ1eAeY7xnXjrxdznbRNjeg6W
NoKjEivWojVj0y74Qgp0nTaBoSEz9A8Uhp3bB5ZxfyC9YMCRc/KoaqD7+OKy3E+0LgRwOY60ciot
wENw+cjbcHCuo7Ta2aw+9uqOXe35wKuOvxaWD+nFSTtP8y/6MS6PZXd8e5keffsrak0wi+x7Hvef
iJ/+7IG0REzvADJy4Zd5RxHjOdbgt4N+Gyduez2bzICUW/R0HyScBFDFegD4BPT3lMybCMe8M9Y+
ja19B5bzlCmTOZT8vFS1UQU9wMpJUmBKrU2KUAA/4feGEVcNpePuR7Kt4/IHs6iyhW8giw9xZ5bv
ylHAL1S/FTWGKIA6IQzhK/D1eJlz8x2guTaVQH60V3PHXf9oRZBwv5l+HTKWiCvx/wF2i2Q4b/Mn
V31Kq9peKteOljEkzUZ1jW5obZNsfTlF1rgdqR1iuZlKp4oiLB+X1WM+ENdqEDT8SDGPl0RdiDmy
QRzYeQtWvED3d3PxyxTgQbNlnLUA08Lsd+0bXguQhh7R+y09eXR1RLbA//GQgFNo5DBJfI+QU6lD
pwJRLWmzFBY4ODiD8xRI7d/yLl6BomsrFKP6eaQVH3PtKC2XIkaYls5+b8l95WZZ8VuRXKmRkMWm
CIvFWZ2FBM6aS1jutLdMiUM9nsZZVLbXA2/qtLGkvs5jwtLzGWEkxgqjbsyloK/mBbikJI3blMKu
1B4A2+NKWEiUUjsNoii0CRujPu0hbUcVasfSW5vFrmKEc6gOWb4x8SfabT0YIUzf2hr1KbsAsG3Q
bvXIGmdx6ME8XKTZ2KR24akQXrkdx93RBNrb63SaotgDMTYwk73mlQox4jxt87sYNjWE56EfiCm7
8uYSJAbA/rCxHGNSTJRxnNPdEV6z2AczKKRf5TWCMURI9Bnn9+IRfc6RHeiT0oNJ3fe5B9x25TNO
aX8Z0CRsU2T0kI9ejPFtFyq6avFR6Mc9qG7kFPWxCS+tA72glsVURARm/3+A9u4cwr4I57G48f5q
CAF00zA/WnltfbKlPfyq9Ww+yvbZ+C6DMRqP87feCyX7pW3DUgj9jyxebbbzgb+aci78RsavUrwy
oLgzI952eyx3d4WQwbWocMyTQMR5VjS6Y60JkvV4mrFimdM1fG7YD69SMOx2O68Vozow8mdhRUVv
8LZ0VVfpYzGyEqKlW/HPw8uxg3Qc1yJHFGvjKO9gS234Geoxq5BxaxbO/Y9UNZu0nXjsFHWIbJkN
734OwsEJPbXqqrPaIxLCtpyJ5mZd+Zk3aIbUuvvqkKKm85cnaXEfwH8n4n8aHaxIpsv7OVtPMroL
W03WN+zVJ5Ny5aliVmWLLbzr5TqJwYnYVxfuY0suduPsgPzuqAkLQ/K6/oSHd0yscNNjuQ2KWSDk
BrwLHd4uRD+TSI2CttXPMIDzFVsSZQfKuiNL1MusPx20UbUFcqDVLf+cxM4WwK7JUJ2DWmI3Jnn1
M3dlRJmi6E4v3M0VqDtPfjAQuXPzc1I2mWNVGM9SMd/RZ0/P5vpVZjp/ZegjinLMFnjVYa2iazPC
UzWqUVZkATevOeA2LqnP8fKf6nL1jVgcCjEz5vBXpiCkuirI6Hvp2n3aNPs4LFJQVaCOjgrrQcLQ
3jGNg+3Jczm6ibkhQVRCL+kkv/EgHbd6yDuSUksmjdqjNIMDtK346z721x4l1Z+gj56mzIq8Giy2
3/4sNXMBriGalRFpn7h7DkVJPIIpSYPNIPF9JTCutUk8a6OxkAC+alviwvapBpZ3z/SxpKwnpsEP
Gg2tMM7oxUoz8iJUbTI4sGcm2+2Q2V6pXy6d4G7BdPIh5v4DzCfdv31sPuVBh8DmjWnoQ5iuO8Vl
n7EbItckcbApAwdRDd+TpHdrTGtnUu5IwuBKtz1cDjsfc4Kjw7VW+cD9YHHop6RuFS5MnvbpJLKl
AV/u7j59jJjp9oojl7NdqyLm7wbdC9XfVdUECMwF6PW1kt+fLvnjKpDNATd7B50XlNaKB+aPI5VZ
yWaP4mVZlK8ut9EOeJeDTZuTEFZRunWskis8ReiEkzfbz/U5DKYghVtQ4l+FNSDlLkHB9f9Sy5GC
OMNooAni6MdW2IQyAzwl1RC3BOLhzTtwreokJNjFnwNy7CCwSb03JOUh2K/JKvj6pKwNkqH9d2rK
ZMRCp+VQUkWjJ/C1p1zMcOIi/g0LTe2C0k+wX6BoGWzOac1D4Pmw8EKwUS4SVRSfP70jzKk4Ngp/
3qNJdoNfMIOJH5LuYJ2AUHOLWwEKLcjnP7aVclb0L5Wc2VjQpQrXLD0+wlcuwjEk+Q980GW0bJPy
zF1vkiuZSfTEPudxb0Q9V+qagKghBL8J2H27IlqgmLP0//bMv9zdl0Q7ZQfZ9hTEQhVQWeUwFENC
LB4DWshO45O4zaeXlO8WrX+l6prh5V7jXlqROFss5oiDuIfpbjW4bvnPYpXa7M3vPTcesBtbn0qZ
cvrdP2v0d5RBvvDZFc3uz0Rb9CdVlAXgSMDZL+2ankdQc5r9qPVQL9A/OMONbAuelDtx3pZiaQXo
ohhL/S04Ejezns9bjxwoLHswxWVx5RH6PaIUMoAcltdX+LEHyMhoobrTknJ19FnJFOAZE8b89JrI
tZi4MwKJqnEJy3IfbAjC5v731lEu188iTTMtivxBpgNYJDaypfFB2+zYYVOZjojHyPVZfa26p0su
qiSF1i3rffhJT1J5Q7pUpClIJksb9oVC0Ai8YfjRYX3WD4IMdLnvoneb/wBfGTaxZGUDc0hnPOxL
5th3hjOU3avjkNRUFhHK0MomVDrin14e//z8y9EvoU0JyNlobV7qtEbml9EJ9lAHkItmc5S6AsOv
BZfj/lubQ5r9JjyRvg/Dc48GPnTM0nWLYZwiPo4ohdgkIFZc7V/uW/gS3hdARR1P5cU1JUsV11j2
m1MiG2kfznbSA0QKTrPxqXbEmfLOeP3SCSA/zAdIy5LbZicPhFP7F5HD6X9EI+VKSt2iGnsE4PXT
rFqW0Xti8E4Z7Wck6C35WOOaSGuUCF4eqZNOuNB8WJj/gzaurG+3+9nZO0UV44mTnMlvGFn8FyAs
H33NXrB3v6hfSDdtfR3NKriMomEiDEJhyjjn8Pfz9KJHsYTB6QKi7giCSm+YhuEsllyr+XC25VUx
L/TDIIq/CimVGSxeiNZJYap4KSQtjTXNMa9lmzX6Eu4+kv8wmzQ/s4/mO8BOScNTzjsV6rta8YGO
xbRgNSvNYipBYCaCuo4SGYA/OdpKlt0pgziQTDw2E7XrjvX/rG0+AU3D1a4J+phUoy/S2bEC0wYc
k9zAI9LaTj2d0QSdEgI4YUnV7Cg+jTso57ulz4zZOkIRMxy0HWu3Zn+9azOBDs9hz2BDdJ2J8Uz6
lI4qMWWxBnzA+3aJwSEfp2WH/S7wHg1GIZAwtv6Sprli+kahcvOhCY5U8+OYW9xcrN71l4qtlm68
/vQBUNZt1SojADtCtD+hwhEHoS0VLIgINqVaNUttbSgNU/5aDWmzyYKrwrAS56xSoTgdIED3xHwO
Z/hiwyjrqV4Y30WmX5n/LZEaddgvqRCykHABUZpgOwAEAgtnV3SgiXMUfHBsDRvOEheutoSvrVTj
eRNBnJhXzOfISup5q60e1S4lCAGtkCec/TFdkM/yvDIpXEHY60EOQm15Fat55RX7n2+6oFFYsyBl
x+VUz4zJNWyu8PQxSs6YAgIhBSWI1yc4YcVqgk3tlsRBrzS3067d41M0jfhLI/05RErWMbOxcxvF
6ZN1PL4FplzbEmj54U1DU2jRHGRImkUbAOp63px+i8MvRJaFVwJy309ENcEEdGg/AZJIXO3KwALa
nxH7W9GjIpMyIDp5y6xf3TiTkwn9mM0s67hCx/dYv3FCdWoIhljFkeywmtkiZq3cVXkD94EllSEo
xN1yCzcZ/YetEcIpJVZXAMNDl8Dem575iiJBCpu9jhfsHMUm4HI8UnrZq+gVgxtKKDGHxJwhoT7G
1odpk8tOTnrBYqVNHMpfIK14kQ9pK6HTYLq29QYfalanXHwpNAA6gkE152NTmsjweMYewytZkUFr
EAuoF9tGJ+UVQPNzisUKIk/7uUn0OSPYUr/azGLUxJvylrmQ9UxszeRjdtkvx9H3Aq2b0xRkXIPH
jP0r4nKo6Zi6E76iWELSQwk3kDJgYIcNxU1okGa0RUdBQEBcb1KTT/zNjI1ai6aLTVpuRcqm8Gan
AD6JPUyYfSoCAVoUVo1guzIuTyQa4gEu0MZC4YIMUmBNxjppul9V2RbHF1E1tJKhA1jKDs0DsWn3
7xiZ0nkZBrdjeCYjFRYojoFN3gfsfwkqaSbOBX6boe4QTW8i2nHa1giAe3fJZTt4wzVycixp+NUg
8/IZy/Eg3TjPDxJM9mWjShLY4ivnbtl8wjS9wlnxMAqzHPhsA3v5o9ju+6KXCvwNNiu65K6NKsAK
SIEo4o6Yt1tt6K2INXNGGMZFRBUYNRALGeCBqtBZ8rR1daqESGxuiwKgmEJB1Q5UfOddrofhbwLm
2Ow+V2M9xpxBvd1i+uK/dKeXeEl58RP4qlqHrFhVa8JmwyofCK8l7o1p9XugJ3LkQA84p5l1w57w
iBe9IkGAXkCvTlg5vb9J0GqSPG4Vwrx9uu9HWFqgekgPnePbMhCbjyznYZVLDQKXVqRC11IN1jcN
8F54s0Tqu21qokQqugfWW97WP5rIpUjdamiy7KVQwlq/VG3CD5lptLR3dXspScxWA5mX7CmvFpvk
W3uAqPdCivQB9sgoQXbjynVcdCmTfnbYXru0mY9jY8kDrlyRidkgAX6B4MLtQlVvGazUmqlWa2xD
m92TikgBkD2P+meTi6jb2kfafxvASbq9SYfjAZD3kvIVxtEXM/TStKtXHUUiFRY3cisOL9cNiIT8
Mn1ilN5K7jMDQ2zEnRuUzWNTQGrk/pYmjQpNx+b2A30WKUrF6SzDieWk52n73eAB/18cJ3bUEaoR
eaSUBLlUFxdLYcpdaEPqPm7nzpkMl3BdyPhXJqqCqz3YMOLutYzhXwFKZ9Rr/6Iph6/m/2IuoQgE
eBORedBNNiWC5KNBaYE2nb+Bf16lPVxqHphkhFrJjO/3Ua59p/PT0rmqHuvn9EeDzuv3ECRDKR8c
4fCbXDS51zrxrpZXM/kVIWSqS6G6Sp56KZO95Qb3B1Nk0D8+X26EbXv9QWdUBtKh8viknbLa+bYP
H8XJuaKlKM3LBhlMgK2nqHq6zS96NVUg3h5fFVIIth6OvnMl0vsU2uU+DTedn7WGUihV4n0C0eDr
SFlHkBLwP+ex+SWAMVtzotVnKTg1BEvcI/0RJX2LNmLR3V5/AxoLO2Knk1KPBfkj+h4+y3FEDFFs
UrZL43+/MQYE9Ai2C8OMfT18I7HhgzV6NxB/9BMmqYSnMzrw/UIKku+MOkLkm8tt81G+xpSiZA+Q
e7oAYn1EcZf4JLWjcK7GzqeAuZQhi7safnqeNTiRL3bxbSAcKTuiLPzPep+6YQBge7fLPhAr2Sj2
6AQ8JXsIUVD1zWIbRoJV++NtyT8f+UH4Ws/eoCpY3qFNYqmPUgvbfrQAMe2fNhtHE6oiL/xAoNO5
bpIk748jc+Z4qux7bGvtEnUcg3Ly9ma7W0UrTTUptJWVcdb1GTox2ZNj2UD9PcQHG4BBn7uhvvSr
v0FKGyyns8Foj4YV1pXLOiB3Ylfp0PKyp7sVglkZZ418/dnxQC4QL7tywBaL7dWucFKCPHeNrehl
ztLiJjEL4qXE6e/y0W1GSlPsqXboQYI6XlPzbE/qh6yqqYOtCHTjQFNZIwmMDPfGPhbU7mnWcIv+
/eytEeZTUdvBWLVyAXSoMSj3m2aaAPQmKGo578KbDXnj+KO4aKiwZm7aIlCsWYGlx2I37eXHKbJh
Cr+RWzsOr+cFtzVoIciB+3t5Hwha01LQ+CctDVqwSneDMHCdS523ZKJpAlI3iYTOd+bDwI4M9Xov
qmlx1zSk4q3B1kjwTl1O0J/A3FGoN/k7i6+LOeYmkpJCqvK+r0L6mJzbgf6lQBnMFpRaFsu22NZG
UjZVKSxXlhmWSlNgFqxsHEnmCfKXXGnpYiW6KmZ3fzhbpyZlCrDSe+2rjPNfamhP9IIk4RmD80DR
NGlLpQSxfcJ3AjvkBZxPEXHDY80BqamCZFkwY355GzRf8S0dVqTJHkAH44/GSSlp6Yl8nGGRIUM4
tO+4u6OWkjV+ElwzhCNNwC0GbF/UjkedR19nx6YIDrTWgtt1DEFqrLUJJ57reNS2NHTD6CDxDcLu
Xe19J2RS2uUZ1f3hjYmw5yqgUTAjNd7burEBxtqr5BHaifEfaZBM2qos9W6m2ij7JvJa8vjdQcSH
6crpwcKgpXWvNqS/vtJ7W6UXoQMJn0m4eyMXrscoxXQqj0cEPSOklTZBgfvBAPJboksxloaLaumo
/EG1FA86BPuA157RcrvgAaPWNOVGr5fsRMYzVvH2kJ64W7xGJRfC0V/ckY6D4F+CrD4ud47tLa0K
6BMDohmpamN/C+XjvHrN9NI8VN7ka9lI/bIc9dOUYpHGDtzCxJcn22UGWHAc6tKOh8qUBWjaVLoH
ui2GrnjniFExXBJAFbBk1YaYNq1UNRWaJ+AHjp1pH7fSSBy1cJtEVQM+3C5muG4vkDViFA1HE9r6
uzlb99NaGDsIyA/L0Q9jSYYrehkS6Q96U5vFqK8d4YWUNjkpLNsSrGtRHHzrhsXjn2uMrCFSeR/l
9BO1Hs5u0ZHJ7D/RHsWpupsb3W6yQjEDjbQavGyva03FsxfRKnF9jTlWrllT3w/UY15NEzOhfqMi
xczGdXUR8c9mLb2VydsiBiTZ0y9POruTzF+TV32g0Xe8mv3ilinBEWa5RX/1rbutokH/6U+Nf7rH
EhXuOUfiRsf5Zi+kna9bD8v2Fx51Re+pknAuffm7tskRKIDo9zEcplWGlsnnx23TaB9Sn1xSoE7c
nNNXE20/c9QCR7orWEWNm8T/8/EDSK334rqbcrHYLa/tkZBMO9PtookJH6lWaazcyR/bw4W5JYuj
yMALprOwnCQ9QepsHSbKvIgfBUU1PjHxpvHIAwn/fqutgOuCiAnC/cdUUVEWdIouxLcp7HxydK0E
vqHwJwFRw/NVdAFPkiSwh/x1K94j8w5ESbovsNZy43AWkKjdG+K2TyOM4pExastAsDe1B7UjYH7d
ZFPzYrVa9B34pwCZUALrHl8yoVagOWA+6RrYKVR2rx9S4+JOoYKxUmJACsxq2Dv4aWhqh7esItNB
7Zi70LddriuWkxTC1j8NCU4S2YobFshyv3sgRht7fI7mZEdDR+EQxF80Qr+nTh1I9pXmxXpmmi55
jujY1mZyUs7cTm40XatJ28WMHQBNyfeU5pA6aIKawN97EpyP6VBq56lC6iZpkA5YYMSuZDP+unQR
3RD8s1aAyykUTSXUTeNCb5Cs/GE3VF2EF2b7GfGUclzc3FIyBpIV3AoclI1kUAxFyXCZ9WDzhyZw
pjKvdriWF6bb5XSDdhr4afAG3yiHak+c/ezzkK9uz8JerC9hFeihqwTF1YF8Tk9srqRgPEBgQkj/
MTD10zuGPjrVIOl0iXmnnRjFkVKPIfmrCyWFT5A+doe3zCuOvLQhuVji7bcfHtBqYY+aSRS91sGu
JIwGm4A0V4NU3ooEve5QwrDgpXW7niN7nCtl3jaD7Pn1/vKELW+yXcyfsGgDPVk5/frncsC4kPFy
cHOLQELipgEmTmfbv/97himhtvdnZn2Xo3i8jeCSWwKWCK7flXwyLJGGXWCi1LzojHAHseAaV8al
+oKnnsxOKNQwB03ieR+LiZyCPwQDbNPR1amZRvF50MB+QxcMaJcxuNFikMtx7N8xuwmOradcy/gJ
ioYitCH54kmwRdh5TPowwVkLDmDAz7X78yyl4PVzEQqzMvsgIj/CiuueMC69gf2mf3uH/oWPNlv7
90KIVmkMPIabiBbotf9iPVleopj6qi6v0WbinkwvDuFzHXdI/JBmL/97u6UJy1J809Xeo/FAScNG
DPiE8MVTCr+MTrEaGYMiXOWcThH8ihYRiHyF/CRE67WckwLeLUNonWr4g8H4Oa0qd6khdwufv5KO
xEIU+94VX1Eho42T7mdgmy7aW93/hXkwK2iy4mOIIKGy24xyZgnH4Y0++P3l313lSNeNeFSV/pye
Yv86OIgMygiqsT43e9oRo1EjGXz6g6oeFFtaA/O8HjfCKWjrPOx60pbotQ9bemMf5dWl0qTsmXYT
pzXWG9NFl5Hn1QMgUOgjXl+Dvh68aVal+8L3kSCloviZ0GisMTumqeEb9QWr81xgRY7CsHf/6LOr
ojmd0E83D/fAJFnjKkYzoFdPj4eCH88sD+iOS6vpufBw/2rtpdpsI9RkhZjrxVDrpGB7T2xeEc5e
+oYZ1xPpgD3FT0bwu6QAjDd5fs+XYh7FYV28jmvHRTdTrEpCIpk1fWC0HqUerMFY4uD+OlN7+hdk
H+FQj4ygFgbe3uXd2z8bOl9cNGifNqJBJqOpmeFoQDurLAY0ihzpq5AcPMBNFPUOy1hAFC7V+slP
o/LfzEoNtvJX0l5Z6whNVm8j3Jc6lscJ8IL87Ds5RDv+Fn0NhtrbkUI8uqUdBQWZ9TXsiF+ljay6
1E38NjGbC90ttes6U9Bq+XMNdmVirIP1s+klQxQGqt58XkLype9P3O74tgnymdcmGVHgv+0fOrF3
h1PfknPkRlQcHBACgVxvmEASv4OuAjB2P7Y9VbttizhJtZfuoE7hMb1SpF3rTr675MzQ1WQZNi61
2Xzlt3h7k2ih6UlLjDPlMpLF9mRAwUcWIwUyEWCvNFN3wjOJNcaiBh4J2VYyOdQSxJZw5AxdPEsl
75fXEPWBoEG3r/GG35vAImOk24zzXg3R8oyzPb+gpbIDXBBKVkHDkbdEv3WgiYrBkvRKa/MMZ3C0
K8tOgffLHPZOR1zrgohAcMLymndCCw3k66IFuJ2xO23nnh0In6YFW+p/Ry6lPO3sTgfjgny6RO4S
ohmYdLIbYknui7lO63RN16SMV/iiyiv3pW8qnsm4zsqtFtivCLHeTwdx6ZnLGtdUglylGlf8yC1s
X2u5ScP6VLU4ozoxz4UI9+qBPHzxOGnO2cRmI+zjfpAxpxeld+PSLPIX/67ctSUTVhrg0eawg5sP
Q+tLUY9a/m89PPZVhvOeqvnAU6HcgkD8XZncYG4qj7cOG+XKV4uHpn9R7GQGYRZXt+ttCUUWblWA
sBQ69uMmr1Ku/7lsJeWm0Xb06QmAw50Q8xRpC/4yL60RZAahVDIwlMdTQqPIoqKvTwqzKK5kTXDS
7H5M8dLfJhK4FgORTN9c5VaNUe5s84fAZnhg6Cg3XSwMiilWolCSijNmFCg9UN7apwO0cldy6D7a
o1X6D96hBB/wsqAI6o/XrtQgOUCzIf2GOdgLJUxYW+7TEMz5weugVG9vAa6sZHykbepxHS+yJpt1
ojG6fqy7CdfgHkebcy/YYTjmhrhVJ+8Vevu1hFSEabz+TTHBs+5yCpVh3cPe1xkD11d+HUC2Xt7S
IQBQ7y0ZE3G1+3ALCWJHoQ0FjqB4oLvsIcNUyHn2drDoyqMVj/Ye5AsVbw7fIKYQ/nKj0n4Tw9FK
P8MGw+Cb1S8izK/cVF4avrxcetA/UMciH3Y0IGmdSKoPl2bZ5dOIfHrVBD1DV8ZETJZB+gfEp+dK
xQ/Ui/03s8VFi1qyxSVUvwJ1ybJRNsRcNjw5oAqWYnD9vSe9JRxSS7f+9/rH0hvWeun7dR1h0xkj
bwJczHMp5Da8QlCBIJQimIlpGIzyDmViA/fjThvZe9mrrTXIvZpAAG3/3X8eulCfNzVudBqZfotg
iZXNTgyeASGYgVwoODhtESuiXPTu9abRWERaiWPSHtxChbJ03t8CJ/1QcZ33VufMk5kXuSyfXM6S
/iZLacquYthjMwGsGbq8rce7k71MmtEWTeeU9vr7mHELNBAF4ooGjzpiTz1gUAlcgjyaKbxRxYXU
/VeRdR0INL+7dxOx7iGAOrEkPktmUQGxdDagJROlV23RBLu/wkP979bPL/bsSqVWjz5MWEivpaZw
giSw5G8sW/mIqcfpnKwa1J8TOMXAA+nizTPgjLhOwBXSCLXKICKhNbhx9A55EKLRey5DGqdhkwJS
I8kIi9sOZIqnJ1eyfAM09pXkaxy5WiU8yEo5UPfGHh4L/pxasutAxX7GTIPQSYbjzolxthfaRWBz
9Iw2BhpLFG+c56xx/VIG1c4C9FUdQcZFHuEJLnq8r9u57qY/18UOVkW/Mc8CMOdWOUgzW4Ywx9Dg
F0pghqDoB01gB4+1xa40yDkWSMOzuDdLeIiwLwt6VKHefKbNhfRIzuvEq4CV766P04HOKDmHDS7h
40E7BScl4Y1cPQlbAUZI3t0RQFT+lwqcSsCUO7GslRKpE9F1PhMyVXOIkhvEtS+x0oksiBc0Qmyu
MUr4I2WvLRzKWvC8R58xQirU2Np8cEAqdwl9u88KsdAuuZSufJo/AX6eTL9bxTO9vZI7NTZ3HJID
sP8I4OZpahuANYzGjT/MwLAsbbiOGntFkL3eG/EoTyB3riLmYvH3yYBYK7h/cYfqHxO0ooY3mxd7
y+tIVv8UvQW+7M04bEvbr7ZEGWRoUy5+39ziX2DlvPRH/axDyTsuS38B2Fc+xGErwG3wBsVIr0zF
LWcSu2b5E8IO4kdPXZDRAMQrSJSspry7u9gWLNqQicOheE3ttZGnc3On7WCE8CtI5Iv9cmMId5Rx
vP3OSLUDn6hgzsw5iUtAaB8HBVMjHDoWFPP/GHiTR+S2IatmWuUJ1BzSgEab4HhDitjuJI3NS2LM
xPqybwfwSlbz67jXJjT/Y0lPAiH1aPkkfXM/RRPI3NMUdIeyHTdY4BFD2m2si1Xnvbois59MT+2M
NKSWZbqfbWlk9wuJRnykQb9O2bCk3fM60N5vo4JGkXQU4au4dMHBj1yQ5zMJPmQT7Hilh5ukO12O
+PhjkU2fb6fxqZjq3CHdmO39tlsRNRUO5wU1KYHLTMncGM1ikFdbjn4jmqY7i6UyEYPnndCQBpME
4EOhYUBCEvj10xaYvN4FWHEkX1430XqWmjdOPGvcvadZQK3HDUhX2Hajr19YepUAWsbL7s3tODMX
74qH83HBf+kGU0nDJ0FDGUE/DnE6fBi4cu7gZpHLLF8ZDh5EO3xs7d2IRf9f7WvSgOH8kbTcpBmQ
VaCnLv/e3ThGj7DxjwgiErkluMUwZf8pGXI35YyEq+QRIZf9aAbLfvkOLK6A2hdfTIV9523k0w3V
b4+GMMaNQ9o0hUmc/nOqtQtJdP0+0uCVNtG+yN3PZDsnN46msGe8+MNYDk7aLRfEwgvk7YcXfaW7
7TgRcZiwoCbaEH7eixBGe4XITwr4dhKJTq0hC3NUxi9yq5pPU+84mU5SSYjBemaA1lRDIyrH3qqb
0LFczvYwO74RsXvxvg3rUeNauAH11egW8nrioe8UWz5sdHy52VB00nEuY5ZLOP4gmPSP8SZPURLF
jj0JdfU8SKhr8rL5beDKg6InQeGrWGWIWUSawbK7px3f67aPNg8fGzXUnyosq21KCatU8QJkpZiG
UPL//5uDmda+v/0BhVWgfivd4der91X3SsBGuQYBfBr396oX8+JihMXcbHHhbuF8DkU7VZ7XUeBl
ha+YFKZAbJPP+00FkMAcxR0urd2WypzP8rGTlVxHr2G1U975sQTUv2TLHVz0+A6nSnxqncEYYXeT
Io+veE0R0zKIkqtuva99rtBpDY4uiyg9aUjkeylJ9xIwzaXU9DbyhnJmlwLJ8bRjveMWOblQVvkE
YgiQsNYiesrk/K1QxKPJINcjxaMWTv7c/XFKiNNEkVphtqs1h9dmVeBnE95Jsizdgg0tWZgtBzl1
Er/85Pdihrz+mjsdD4D+vRuLHCIPvKn5ix77oKJGWuyTQZvpgvULK58yku1RgdqUFPrsUMHu3hrt
Eq38rlspnINuMRcIhlBRf/bp1y8Mj0p/WlVOUfR/CtodGwRutB2z9AChShnRTC6HjEZdxQZw73Ak
QlqmZPgchfe+AZL9MWheWL7yQUbkA4y9Ea+lwOjzemICDS0Lc7l7I5uH9WFqvbdPeDkmErJw2SHT
Gmn1A9CTRyw7/lPWAf1yjeb/dyCN/fUgj+BXY/7jiJTdOxfUqVaM6YMq58YzraDWqrmxEyv+6ZgN
gUfuzUZfzdAWgwy2jWRSgvkPkLy6ptn9WsqgRkbWziCavVklF8vCGl28K45C5LAtuvpgryXP40kN
AWuR2OJd0LPXsI0saTWjQm7Va4HVZcVrQiefbFW9WVsSYzrXUeiO32PuJLJtobKB7SPbSUaGEv9B
ylfeOmoZlnfPymyB5QMbYXVepQW1ChAIUaTXx72BfjBd+JreMFoZUftazbrtFPMPVnC5ybmA2LNY
k/s+lpDuovVYJx3pRs8kTo965E0S+FAGuaoYxiyXJH/XuP6NHuEntt3LYXMlU0mnqwnc63WNUoIz
83lEHOWyzG6Mp9rAFwxzREhiq6WxFJk9bD7we9O6ealk9w1XAO86B5/voXqMMC2hH0LvWQvVWiSa
mcTjTP14S4pXyWaq2oIuXi367aGOoG3GICSjUxCnOT6q9qURaaFFVDD9Iyc/T3ie6kGuE0Mr+IzU
39mSYkXR+zWus3OfcJQ+nef4jARGMgNKBbY7tYBtHV5d/R4Mj2pBo1bu3S3YBvdNwUcA1+PrptPp
moZXkr5uZCr7qtrj6FpGV2i+gEmzAl5b2QFMnDzxbkZxS6677yZ0JhCLcqJIgcL8w9U1d0tjqoO7
zb2kjw8sQA5up4Weu/mxpJjvTK7otffQTIEiB3Yj3BRhYWgfNO2czF6Md8Iy8tEq0vTv4b349J5+
vbj8nSSZAtnuWhwCOb4IYiicDrLKqxQjigljISboYNQikJgAc1d4SMk9CrF0H0Rc/KPKTeCKmgjW
fqnOERFjkUwmqt/FmQ3YEgXIIlUFAUpDYnWxUsQ7qJscGmt52LXLiXQtA3NnvD0iWlHHvRo/U7nD
cQpxCoeiYK0CNOxWdPN/mBbNjReVubaXEFQmAGRDPtzRVJHH546MosxdM/Bij8/cnPjJJqIRX9r4
NV+nlmdBchHR0jIus97dAs/byr7veuqImZIVLMDXlEqysTHIE7eRTUo1ChC8cFdfDAeN/jGYiJhv
hfsCcoQHPSosvJmnRHSNdLEAW2rxLHRYNTyXEsdPqG+ckwLxwPQCiaA88is3EE/99nNRoYYwu1vl
3ehw/YvJj/lp1DM9VotaDch8Li0VbGryA1Z5HyyKSH0Mi353UREfJT9AMZqcBKd4x30RqzM+Tqeb
U7ePkzEDKRPC6eKSIsP9++bDyLoGa/FTU4Y8+ySWfhjvAc36NuRzU34FQTIewTwH85Y9DHZ1uhQs
BkXHholbGG1kAyBLLrXYSn01MYLtFWu1wEOCcrYi5UF/rAmJy2yr7sv76YpBs2gynsCTRX6CYIVe
O5269vCjD1qXETfe9eDn32JoBK5SorHrqMsDL1NkQZDl5SgQ8d03ZEfrEOk2L9nD6kD61lQ19zna
wwaJchVY7hAWXzwDkGheGFDYb1VCJkI1BSVc1ckF5pg8ueko6E697yNs0AvNXuZPKXbxnn5a/YaV
RaoSUsyyu/crAQj5ZnJu3ZBlpABEb9ZHSullh8dOVSOaMOajI0lJVz5+GTt5T6MPgw00I07FDYlD
Csj2OfypBM+Gqg/yK6+hNKO+k0W8FmoDP6rFDQgG+57njsZ9Q3S1k79zIzIZ4fMo+S+KFdq8bJeJ
MxWq1UuF3CfpvzgFeXtc9QbnfTJQNWl+UdT4zK7dAR36fQf4BZzJahKcyW/fai+GIU6up/ogCw1/
b2vULGCl64/9cmQGXhy8p68/zlzQnKDcghvG1BFA3uFEXOYupt6lOw0uuPjE/3K7rcU4nKfMWj+m
Ma3dekVSzuJCeaPpHNqEByMrzx8SQl1cSvYrxY8iixIh3TATbmEM+OeCKj51ZR7X9Ht8myU5GQ82
oXUJobrYoe+8sDw0rMDdPyHct+kmJtXt5iCXeUrgNz26O4dFhiGQDaLlQj9hda8WWoi6w8L93LUu
Q9XEog0DdTtZjuDSqfLvBtc8gHWt7bnVQ0JsCtvDZ1b4YTEev/1EaGBnh7iztUIxUsBzOTpTfghU
j6Zk4HYGckewhGCB0fuMvTH1punNBGMWKO7TNoDI3WJidGP71Hy729YtdzwoICqlYu5iQzG1JfV2
3L4A4lvuwdzmV69ck2AjrwIU05w9q+ix4+ulQ80ud1u0wsWVk8IeX5DROycsBlI1gvAxb62Ys3lx
6g4GfJfc4mAhOziyhqpnSpr0Oqnf3El0yRNkQM9isbB4D2PimjNKY4pghYziLv18Z2lPJdulr+xM
63iGT3HRLN4p4Cj7FX/ZRjeW5eTivNd6A00/q8NPY3+gMrgvAR7jUCGoeBrV3JsiIkyffPjDiQ99
8ew7f3ya40vXCOK+2fQcdd3VQpph2ghyrRP5YdDShNtv72rGbwT2yNPott44yHemLYH4lpFzKPEq
Zsi++pq5kwmNFAplMD5/BG3L/qlf8GQq1u5MZL4Or8A9Akr4CIYiClBdcF64JFXupph7ZP+Uv1mG
AGprTRA5xYo8EgsopJTuQPJr8DHZ3t120gyKIBENd9HDVlQ6McXL7pFjIRZJGUNP83+bGfo5yUWN
WtZd69sou4/xxj88WA6dOmQk0R0W1YjXqAT8jt1IZuMISSWQFWZAUwVWsAIshIRyaYSYf05LaXtZ
w+50OSPOlbx6hh0puFntxj/lZNR7rPATUm/+U91eDiBWgSV5MWcshk2eoFsQvDqpbZ2RYcHmqHBm
pOEqVE3x06c8frAuFoKlBYoiTqpHgAED442kuFsMElnvFlJghvlM/yQvE+0JiadxN3p5dxPHaeQO
5cnKrvR4/fF63XuT4r7SjVZQm5TlPid3fLndg2dwZlamo2Os98eLFUFmi+cCvDOotIwop6ni7u7Z
SJiSQlSJ1ra4mxJ4CtdflRiCFlMe2eZ+4pD9+6GuX0TpJl8KbBGMBLMecUeRxs96pmdULBso40DU
eSTXZJ2TQnIJHXpr/83pf3CTmMQLZCdz0WVqCRW462vv3bgxEQpb/B0bHZH9xkEj6NAlCyDPzZ5d
W4KneyUqZ0IhLsGjCB8r3OGdAfns0rPm3TPcbojZoy5pc8e+9HoAPwDrt3PZgulVSEzNOoeUphLT
e3T40rVGrFlc4j5tB1HILa1wZN1nvFFoCj5AQlY0qiOnDFvaOzLmkt92UclkvYALg6qMAif02Bsu
X5ElPQrkns4fngwqsljQvkVj39BSM1zCJ2qSq4XTj2WnjsD0olDkfdkcq4iUzT5itKgwV5gtdkxZ
cgiQ+BJmfpkco/HwHBXCaIIjcTHlTucra7omHtI2hetUSD6JLxTD8DH8bRRvp5QiZpJUi/MRVXmF
Fr96DCgtYpsAc5G1mYfutcUJ1cF0lf5Z1Q0RZjkMFCmyTqR2yt3fnqBYXBfQDx+2jzgXZngg7KYY
xS1j4xCPb1ymDx0C5QRC3bNSiHBUJfK2kLYP4jhSHmJvrrBHLkBTsvdnJFww/XM3vuO2pbezFfoA
EdVt5tTapsDZ3/oWjzCQqrQ5vys96ScBC1199G9iwjzSfnzDIVXKB60/PVE5XyvMaZSUf1Q8zFo/
RyCoj1m4iES19Sjs3NuXB5Q+15hgXma0To0ox2hC6KfcYwXlORlbVdAOPiaRqhVQsTcLTgqYQ1Ax
n5vJp/iG4Z9AGB6Tq6sBLpujCrkbD5G9iOA05oG3mdgrs0O4EtG75zO+NXD8zWRQJglgYR4i602H
714nGAj9+ac0bWnWkwCev8XDpnWU4u6WWmv4vLKTI9JPv+Dwrff+mFubAgRu0MoWQmJgVzGJNlIe
tcxw7aExSZnCsr4ZpkpdopGmKTfS7nJ47XYh0UxwBcOWamH1t4Bscc2RsJXIlV4xda/4/X+V/+Jd
n3QGJfrmtWHckDzsvdyR0/4bgN+0unrQonuEM32THc0eMYd9cs48wM+cAnHn/6Od3q9Qw2tzT8W5
ZOA6RAHbeiR7pVmOvnTg9s1d3cahCGIqHAHAx3bPuHP+PpL6lZ1qNr6kr2o855bcgJTLRfX7MJN0
HCpUlbA3Qt/xmyRIlNQoB/UXSN/lVxFcNzKP6fRBu9WcnefrDzc5HUBGLb+vtPoBuwiCqhHSb1Iu
HcgfXFPK9zpJvrilt5FLYaG/pvHUV5SSikIoC4y1rXsisgLkfdNRm4zdhXvXmz0bAfUJPTlu1qZk
SgAk4JRjrnh85XDx3wOY0BkbY2piokduvQJ5VFWurhYFWUJBqGY5J67bkx34ZpGptEVpSoKzfz7R
ykRJonrmXosgaKDuV5QNjOkZoG4DDk4flguRXHwZ9zJ38Y5Dw8DPmYUkd30oTNHGn2XQ0iFeQl0L
pqnr/NQ5ShYKnM7ERyjDvYLRcoPpTYAo6S+QcEgLPzwEgI2XBZ7Nd0+wioOjHzRYj1m5mxCx8A3T
E7VpwqngC6so+UHNITkJbytN+Y6/NRUq/PQXEGHxbgk7gR9EVF0xA+cZ+Ke2THOthSeU5vuxEm+B
eJNmgomtRXO8RNmmRoQ6YI6ZgLID/ekuznZd3ct6FLT0wSg0w5jaYv3g8MmshsWQcXVZwI4zlaGt
yq5aBZol7lJiTHiig2DZS2H6XmZGSnXo/5cA8KLwcloGgdPe7Z3lM7/hcrwosVbskxqHPQCzpeAT
2Ds+cKY9lkjnqyNGxjJSnakRmekbMWEVMaY2cxQz59NYdroesa7Qkg1LsmcN3xDSTci+hU+Eb5qU
tQi6zx88uYnz0O5vHW7kNFTRbnb5dsWBtkmBEkbk5VEt/atRQoDUII0+dlsbXSoLYsZV0ZRq/nXK
BSh4qxLpmFgrZ1o2U8Y+yByhei+ix63h5t0kL67V5aWsNz85P+snDZqfnJVxE4RWTs3ahusmkgpx
OgLnW0A9XHd834TjSXTO5PBaGxbqRznA/H5aK/X79h/+j+VWYYlP1/kN7orUlnV15PgTdSLRqzkJ
jGZTiZF968Eu1JknhQ7BGM9PexPtsq/KqfClUfh7QcH8QPrLIIatM9DFP8nVm1QMGOrnWTVoKQq/
SPTsIEfieX7RVLvbUloq6gJLbNAecBrzbJQqY8RV2762S4ERCRbdxBNNVqi3gxX/4kpkw/KFKKxp
Wj8KiShz8MKvxyogz4Nf0RrPxAC+HK3+Z1ObEruu5ZVHrGozwgZN+GAqT6YWTt3jBPuLPzqzBRwa
Cklx15k9hKpEWGUrZZk0CO+yK9duGdsil8KxN+e1H3TMYoDOs3QjCgdgwobPI456/hR86mKpCXk8
Kam8+zr0bHXZgwSa0Qu8JHJppkc8U2XWPKIzSQrdPW1YyNIOnEIqTomA8x8q9haOElTjbQOi2cZr
f757IPZ+CwR1fRO55vugKNfjOmoKjhlSJo9VDElg48DznoeXJIizmbyGFfaIS02R21AI17T+wDU9
rPBCL+eMeZDDFWlgHIyRjJ/4nFBEK9l5TAoIJHY9U5E4GYgYa++ugo8v0ZcPlA29Wxy8rZAVPwDV
1LM2hbgJ7iw3xl7PIKFwhEgqXAxbuJWY2w9zkjbOUw+FjtO6S4kdf+3AJx8i3m45GLukmPhOMa5k
MpUPRvXaeQiBl5SZlb1VpUi87R3HmRk34qy6zdhg7RYaOK6vct25w+a82C0pwogxUU/sJq1VpyS1
jwn3xHF3DjYURxSyoMZoyaGPiqCl5ilff6Q2owtr4XRQeKOOverARYAsgnWjxOpx3pVHNMz/MyDT
Y7ptEW4VaOGuqQvfap5q6tIeoO9BHHru4PWexw56AHAJOV3rSx253tUAQ7FUt89Ne4dYuydAh+2K
9mnh6jsmZ7fOxk9K6WL1PP7Yp6vJKWbQmEoFNz249ijeW/JKfxiD3YT58YzTWiLfSo896EiAX8Wy
ucWWe2rQMr0IsOPw4D0NXFiL/Uo5omsuJotuRHqUpO0FvdBl93NiGBQpz89eZ4mHtQDPT79rrq/u
8Ix4rMYPaD4r9R9N+LO+ycACTyIGvaYWoMV+u59pripqTCF1E5tmOVeC0o3Ei8NMBo7s09GUQcwf
FUyvpNPd/zElEL2XE00zH6L80PyLseATnnuWOaSRYBlojsOFljjqIZZr517uNFq9TmMIksLaTg/Z
aZ+6d+izAGFjJotElMgH9Kn75a0D6M08QTyMed+nyyekdImBDBuwJeUhsrIHLUjZVDEZhw858tZC
KxSbNWa4LrvlYVCPDyP8lUH7TMx1FyWVd3nBAYIy8HMDbqYSW4xIYBLWuLFwtVP4Sx+2tNOKX464
wri06S2RsjrRpU5whrCIVGjlgiJd5XdBVcY5eZsZu7ENQEueEH71RHmpnT7OudGOregQigeh//Sc
uA4WzHVm7GdL0HAS2mma6P/AJbGpQGV8rfC5nSN1IuWa7Ul4ZFuTeiZpb9bd46UQftjjrV16g9ph
P0Ho0ypv7NAezRCQ5b0JPS201pAcSmnnXbFe6xWVJ52FrtDSs/5w/9RHIucjmsM/fmDNjC5/SuKw
wfH4mGpYb3l2yXS90u6IOia/b6tOa0czSgS4k3Tp2EsVzsfAT4mle+wjt1HLdT/B0f7qqOvhRdLW
iKJ+5B9DN5hJzzGcKZl01+YoaSGEWr2XTFdrq6Rl6+o10Gm+HyFWg3MmpzNDL9PchlWEHiyRZkGP
nWohHNJj6+ww2MY67Tzhv1RtVCxilJQpknBs4sVMsiaCITziQx/Z4T0W44DBr7TpWAfxOKjAASV+
TqLYK3MUb/pzaXk/o36EsAhev4Ra0TMIdzQp//u2G9tlTIxojBWkNJCTX+yvJkdw79ObMOAfzics
03GD6Dbx+qYJVg73ILl4fz0rejS6qKTBTQAMQuWSlgSUInvEK5sYCbv+7Z0815OBfgRvq/065oZb
F+NiLFfbXg0H6f0egxZmc5Wufv9VUzJU2zvdnHDI6Mw86Mpr4qRtP8BgqDmM+AnRIL81hfqHWmip
RImrndTXQnIKXstS3Oi+pz1LpEQbV4xCgZobHPiqhdENNZ1+NlfB+9LiAjiHklho1dyF1tHAVP6O
si4D6HmaXIY6yWcpn/cBfttrGRtG7DOnIdAJM6V846MaE+REyC6gjrCTNCX4/WwdfkBTq2F2yQ7y
DMlzKK5rHBk+9wnGfTn+2EocDAnm5n8QcAiC7s/wSCsMX6RMI74cPbqUYoNF5umXxBIMr9mnkxeT
zTVsw6rwmtnqxB7OFnhBGya3YQqMwesloEd+UQdFPsMA5RYTLEodPYpVbv5X5CaTglRAVJr2Mm99
Y7c5fKGSsFDlf3X17CYLx6xtVk9/TWWVITwSEINXDWPEc7gKW8rj/BAaPb9B73x82oTfn9RoPRuf
r7v3K3civQT1Ex/6AGIN4HQnv7iNYOtDj+h7uYEFuxjQ+LbknXqVJE6M+O+Jys4G4in8jUEd8jXD
nEp7mzy8lrmFVJkdVA13JiOC2eqjo+GeNhien3VFXwe/WK+WhNpJCYtS+0PilxtgEu9taRxFhCyS
nR0pxlItEEWuh1nR24+lSHSK3WZioLlOVIG+Mu/UMpEJOssYt3D4Uee+dXvqyGTH5AxvuV9sPrCR
c8QrZ7tAGdkZIBzcj0xNwxYTqQnmt6RgD2QbyjPeBfBM6VeNUoxvTZbAqwJPUfxZK9JefAABbYZI
qSQUvR7Iu0jcDmMKXUvjh33+P1EcXEQUdemSCS8fac3elJStqvh933DqxUZI5kmEFxTCOOr/9RW4
UTnwUN7PHNjydEeNzOYKWMf35J/EpQHqIo2IyphGOdDaFxA8b9amHi48GEhSXckPOZY8+TTJrWzo
qZTcOGHrvg1YS8gR/hw3k/KeAjdtm6y29NBAdSUkDmG4lxVHTovwWkYg1dGaBUqkhUSXDTXOsQ/3
Ajbz4nMLgo1x1p0q5YTit2nnXZSXEXtg59ouvvjJprywGC7KiWmnajefMQz4g7U+x0YW6WEplslE
gzOxfy2F7/xyBkXzdohB/3ovbhP62w/OuFwkiv3VSkobOXNZmv5cCveyLGCdPDnQkDFStw7P7wYB
8ECgo/gu1ODcRLPEuRaN+8yY8/Pkmr4e8FhdBe76YwDykq5D3oPM2eg+45yv1wzCMX2kE9kpx9el
8v6IXXOOdyoUNVPfw3MuHxV1OJImy5mZhA+xvTca6IEuVr3H62RIcgNRwC6h47bWI6CmMcEhbHqH
pWyxnamoXwrIJzsgh392XATmscw7w0DobgJ3BR/FW2gKTKzR8ScE96UYZsuFa7/R8Ukai/YV76gH
6UJcAgB0vk0lYflsZfbctZzsFGlhQ37MONzbtZgew23I1CVI2Q4tsUgDXlqnmyQ1gtiJHQObko6L
kGy2MrG859LtRTsVoG+67HASceNZaIxSvg058BfGO1pBTXdBGdxb6zvYsKuubreuCVc3QKAgC8mq
kMmsoo2BJSLvxnx/qornwnk+Bn89SzGPmepOl3lwKo4rnAP9C0LegUKEp8BYVei6d/urze74tfyD
B1QaRuZ+SALBtuYuPUKzGe4taFFkLmtHQ7DsDZZR75Y+5gIlr9/vxr6gTQqAWI4o/n8+UcObXVPl
ZDBZxo7kFebxGJZ6G7uvUNd26ZQo4MwXucGPs/QoriDRncrOraOlYnz+BiIKCCIVgtV52/mgPk5m
oEQcd6DhnHRIRdNfoUNExnAGoGPnkrnzW8wWLRzFMWcUQJY+1zDS3guNxIs4no5t5qiPXOPyUeFH
x9IGSqAdGMW/PgeqLOWVICX5ud2auHyIoAVtvUGmLvWa7H2FmUhhesCfGZq+k5CDXARanlnL/gzr
4t5FhxBjsFjJGQyrHH1YJD9vXiE2ODAno/FlZtb+hMXmLQuQesMJK6O18keKetkJMOoXrkFwk3yt
pVmJUxVX9WqdpMAXQpJNXS2TQslKjq60IqoUKxagRPflKjxWYMHJ4ezYXxkVt5M2BeLZbWavpHkq
nzEaqGJ/JcJEaLwLHsgN1jWXpwDdyBgeYn8n7LxZN3+F5L5ZIDzHLpNWE6iclp9j4Y9/uMZy/rfd
5+QCHE7XeIzUEey+u0sHO0X+ftfAY5sqXDy3FeZ55R2tx5IbHsHRO/RRzE2XZF3VWP2wVoXiU/FV
4XqvWo+VWeUl2Y+NS13n/eiRWTmEypDsaYBgXbrbsgI3KEpPalC0rBczK1qWo/UKAkY0Z3S3snQ7
e7cx+4enJpTMSvvRh2S8n8/v3LxIVX/S45Nud5yiBIBFE/oooAxUUHxHh4rds7H7AiL7thfAS8Ej
141lXp3s2TfBPfrPZqSUzeSE4jDWHPcpKFkQOaP6ST1FOUdtmDOOg8zY7LfO/hdvP+h/M1osXf+Q
3cr9bgQabeTVZZFDvb9TnJSZki316OiDPBQUVwK73CfLygcrU/clMaVuwKwegXOvhvrAfZZoNdJC
WZnJXLPWz6e+IZifoMmdZVgoT6ZyQnxsWB7YCMs+9kQeIJNsOpu0z2g9E7L8ow6Tgzv3vtwBRhV/
k4EA7DE3QcKDGJvHsY0aX6BGJ/jXTVyvN9WRv9yrlKrX29MKcQAzLtFAYe4V7o1vqKfQW7gDb6+2
C1Uh4aS5L+sOCJIw/KEVSa7YVyGjfzdfsXXhx0blBKoXYOxyNtBmqhXYl/m4FHWhJN1GN9UDon6L
kuFzENk4c6U3Yge7ErbdJ5ExspsO+jChYxzyTODxMiNeps2zrEocYM7UwSBkp8XMCVfPDaNFqL0Z
OGB18oKRLXQBFUrt62G3+DOr9mpLaHW0jzwIA8FHsrR1Ay5E7WGsXuKCdGGZYZPYtI90FwJl6PFe
5Tld6plvj9FQOASWLR+ZLdC0EJ4KPX0Sh46HwsSFg64yr6fkGkxHgvmrH/4u3F3Z8PUeqAHDmVNR
hQVZjcgpw5lxCGKjogkfsNk0lNElzuHYCU8YMqvHO+jmF9BpOlm8gtbhqESicRLDiPNqES4k6Vq4
LvsdHCashzTyNi/ZJ9zdNAp2LBecxvRnQfP/fjP/qg7lciECCDa5nK81pEFZpH5w7CUgHLLzOhWr
dhiyhhmMmO8yqJIkokv1Ctw2BTADBa1rKXQEMqZnciYp2dVa67VYqUp/BI02wW9Fc0eeIKUVK5hN
QEgEekZli7L7OEnbiLSok88WmiSj9h513Op/l3mWejMeA05BHLoDmVq2Yq5eyIDZdq8HsjUrwn6l
vPiVDWNxxcLaVHrO4YkkY//c326XCXNqZ0kDmJdV1vB9oxLkzgf9oOYgbm6LtfWxkHt4ezclin+p
Cuse3noHO05NGM/7/WwfXiTgh9qe045eByAl3QvKRYqBKnoPjibCEfc3827FdJwRD+qwceM/6KXL
esZmxYD/diY8MpSamW3cbnLZUplrWRC/+neyc4XTbwQnPRIFTZYAYmoJsHTDYT+pGjOlumCmQ3D0
S82lbcCrHs8z9JsZlNaTohQK9xpuNuF717foTNQ31MJVTPaylofynpvtZlg+ay9GM/6p0TQrkc1J
vBNrOWBiOEUiHG2CYNooNqQXQzHnrLsn3/B/ND1fJYGFz3TJTpRZj9jhczkTe9JIsyTnQN58YP2e
hzRLTJ7LMjrt67RcWtc9d3+2Momt6E8yZuxZFq7i5G/A7WtFc8jVhgiASDCiue3oY6EQ9wvyy3up
8wxqpi/+g21e3yjSsx+5PEp7Bh8Sou7L1sbLR/UfbCyhvzoilL70aHT2gSF6hEYMVjMnzud16utH
xyjJwkVqYCMbBb7FRJBx1S2XqvBXnLNMxSeF3vmPThSIu7M32aBkBEkN2S8sHLODGdFneNlXl46f
MhqhJBuJAGNRl8MDyLcUwh8QEACs1mLbpO0jnTNIh5DwXptq1QnGuwWg541Xlhm2BtUxItQ0+M7s
Ogy32Q1wNtMEcXXl7ojabJl4C86DUnwaMGa22KvZTnEQ/xT/bB/cITm/J+EJmoM9E04CYJVWrSb4
JDGeHEP1DuHXo1QEvLoPy8LAmirdVfUTGTpChNWoGFCgPRZV9tLZw2Pu6FpAmZe7u7gOrwT76RKV
8ExN0NeIE/9CFKwQPr1EXCHSyOmrYgUem+V7pt9FqPs33+9zkjBYZCfsi/JzaIsIgF7i6tVkGhMZ
7m7x6CJ6my/A0bNAgwP7AoCPkmKsa12au85cWLOAnyx4wSnC5sQth0p5VK/3MxbwVAdpsmk5pBrW
SriOZMi3KBIsPowJPWH+e6LI0gX5f/vwS5izKHWcSFGqzMZBhj5xCWZ0TSqCboOk2JhD/JL3jY1Z
hfcDWw4+YPv6yUqbyNpeLjgZOaACnxXYDVhmSp4iJgArP4mVrg6KCbMgErtev7fh+hnibxAZWTlm
nA4qOvVdGNLpaRkUitPwYsgQfYCNnf+y9X7ssyZCUnEN21zEnPE9mMYPMRYcmDgTfe0mOwVyS04L
bMTliKHbsq4u50fd+17YuehqmuZHPyvBOxTJekSB6nXrdkgerWHGDLcy/p8soamolsEcnbwLbvNP
VABXrkzEVWWJP8hu+1CklwN56ZehtT58O3ZySjwmZsZEX9U7ZG0JisW2ecgfgKV8kFpVO6m94c7N
OFBDdiBLGPWWivwqP32I73Mhbq7rj9ewcQ3JnSEVtg/fQj3/JUfNnxCv7x9bUaS1S7hb2aT10iPj
Z4I+kLF8t324eOM+YsKoSOWa5OFfqoGRM0DKTm8+W8MwTbh7D594KZTMv6KvwyJ5to+w7t5Op9/p
HydancOf+XR7apzfGZBdKeBJTQWx4JsPXAKUteCjTUe1a9ZwhEOgqtr9OGUQD5n3XzkoFyjY5muK
vibFPvw42aSTz2f5UqAljGMYyn3K0H9LPvL90jFW8LnTHYPIHsNY+zfCRSKCeuQGlyRpdLXS7yRH
w+dbrONLoM7PlCDmKB1ojQPhzKdCSXdOgM78NZTC0bNBvGk8TDG8rs4HERZkQT0W+YoHDYVAUCDD
2PDJKkQbE1rmN2ujL3bhOqUZKNmNuuvk6bvUojo99OCBVy/K23AqKZ+KrRd8R2Bysf/44iDIlLtn
LYMRuxyJmN/s6F6Onej+iH+tjyVMRXKs1QUJLuURNowZrdiuVtnEb1w3OAdMcmxxW6P/8LVLCma0
LbEkhSw1mzA8KkC4fNXUNatVQaPAOBO3n+GWC5CZWzvKR1DNAOEX5/4WXVPh5jXREzR0Ehmd1q77
K1XCKHSmXgu0cPldzwZAvb/alyWJc7Z71RaycoJxR/HmBUITqcFvsy4UcS4rMynCjTpXBlrxkRRA
glQzgMgWTk1IZnsNFgFHDrxoTfUhhYMdIwR6Ice+Gz1QghK/2ztDk2p0lJjrb5QD5wILYLHEFr7O
IlUxyH6lXHsbB3+E3flEevgZUuGfllyz62lV/S4RCs3R09DpF4tDAtqT57EUmuWwpWhbW88WvGLj
stR8LouI1e3hie54Gjv3udHfgYSxE5AuW1prBVpub21hn2DHphztvmodmRAXmI2+KCznhLzRs+3i
k9RJyzDbomW5evRP99uJPysGpWY2sr+E6QREcB3N2eM2WAHJ/GV8HYpKIhfC7r2B6/4Sa/uVxjY2
2vRo0mUORgHk0nvGK7nxmAZnKt/iVS5+swE1oSqTRM2kiCwC4z/EWZ5Gsy4izcR32yaLSeOG4pYp
i6d3lAUBjlcTN4IKi23lNVjNcBtMZG0vuFRzcv8+aqAO4srTzIltkLCykWqryC9oSNbAWS3zXapG
5/p0m1IC4AY+WduHqdTWoMaSExqVNsIstmTYE1MAGMdsdPkXM69fZjDCM7ZLeOKN6tSZcOIuyk11
AulCx53yy8iWq8nUxk4RpIddFzRLEH4vQA6O224stxJMpDz3Xo0A/+lgTPt5W/r0s+f1+gNLYaxm
BQJd39md0os1bMGfkT3YkJx5FNwyQuWwBWKOcyvQu0tl/cxsJPsnQo/+nxq2WZE412iwwz1MskC+
DYCQZ8pOAogQU1RTVvgQiV4M7yZrqPlS6Z02w2xBgIwG7wOso67YmMdTkGH9B6/ZXjlmAAVcZOLM
DFuhJlbfsRs1jO9MBJX2NYsa2isXccLXYuq5TzjgnM0U8LXXcVYxFyKn22BCHE2eVAcUsJVr/CJn
7S7U+0M4KpIqLq/EK2MZhjZO5BjYgghcfQtnDaqdFHuQ0CqmgpC74zCjDvg7oJn5WVsTcIEW2B1r
wJoVynPO+z6ek7yyfny69hgPMhq2Z3EngDmpgE0lDmn+aCBlQbHs5tw3joGg2KPCOFb/cbAt3K5n
9v8pZx0Y08jLrdtQCBzM0nk0TzDPy5VvrikxgYbwEWNpSvyZLLd3l/EF97aZ8ylrALLoqWj48GFD
Fz9xhZYF9fNNFjkmgpNWDoZfOwt5QWZe+ISMbktr5mJkKWxwaePz7c81DKFBdCLd9LfZGcgHYPEq
gyb1/HANv5s1fLAb4rt+CthkipUFvNDmZPJva7em8PBKvs7eHwY+UDxNE/B4VDB2KsMQ4VUdgRyp
wwReD2DE3ovTFmKscv5K82DC+hnJmf4WzVDgzRuI+TwJVfwkVBpW+4sw9H56QlxT1CtEsmEzVHn5
hJ4nNxIoSOdTr6VFyr+HxQ+a27gD1gjDdev3j8Gzbzh30OZOxZ/2FXMdoRMqBoyJHPIkS/ff947h
0ntnkRQ9BjFfSwXu754cpME9Dc5OvMo4PJcQOzvfWmJ0CxlnGDmVTqkzp3EcAuaTAMfkrGUfMt3e
D9aEyPykxjRMjgWNgwgYnmkx+UOXUxWoqUyuAZuunoIhNO9DGf6ZkZcvaDlspxeu8vWqzHpEIbq2
hrDQWT96/CdI0eQ5oBjevf5qjkx3Eij4dd5xTwpA6YEAka9IAeItqI/UA58HPmAcc8def+BdXdUl
lVUV/K0rAW2EoL6QqoL3FAJJYkDK11jmj7iDl13FxyfhtD+d46ZT5yGk9G0Rx9LJ3GSUTE6B5jMx
HmBvllTTmfeI9PFmNYtAfNAQXiUQVB5CPUm3f+6I/SzX2MSVG9UXFhr8RoXZ2OEM7j1Vj+Q6d18q
Q3IrbH62YNtc604XBW3+ApFHcpcWKSXGKgooW0D1Gv1pL/20Vw7mMU0cpx63oTJCEDJO5whA/gJU
CWFUrpullGmDSmZLJURo79RgHbiBx8fHyIL2lM8tJ0Ipx/2GbLszMPhkdrswqsevmeVKqxAZTlh8
7SPW3kRilHYJ89L4XKLBfocIUAP2TA6kPkS5/L6N0yQkd3xfFqRId1oHk+xvO6zsBV74ua9Ql2wG
3jGzWGylFLv+dL5D9Jns/va9PUoNcF1gjjwOLPTb2UgkIjjnr9PaX3HIO0MGcWFjlFMwDCg438+D
2KkSNO9CgMFc6Ita3/prFIlc9F43XPBGFbguRxYOxkxrLd6HZqVq/5SIrmSrzwtUw/J4F9zn92xD
WYGE365TJN78OtpsyzdE7sUKUbkpiiI8a5agL8CszFF6Y71DGbeehU2G65MlHBvTyR9V6oC6oGsT
rAohT5fr8URlj/P84RP4F+pLIoXIk1tqd/YghRae+PNKm1PuyYk4Rh7H4hramUDSUOB3zd4N2uqk
3RtatSNKP8zkdER9zU0AE8kzXcm6xs/HeiKEfSVMmZUlD9iL6tBW0JwO5QrvL6cYe0kTeKE3OTaP
KiAEjgMw6cDcA2IsA2o6uzjKYFVF4y+c8jB28OjK9tjXQ/6gpWhC47vLRFaY365qSit2jCyveMpr
jFcX/DXuvKkuJUM7FSPBu57sXIGyV52GURttzWs0jvsQlc0YK3aQHlSYRUvtbPukfOUoDGPeD4AS
K9sq0CKmtKZ02ZGYjQQClCY7fnEr2XXWCVkr+361mNDmtT0JAEu6TgBR4bFBi33HsJ9oElWMytuO
ybyjYbjEu92uw2lkcZBNUPzjwrqXFUV/AXubODywMPlgJWjPnMGX/P0XrSb7xgGhqmUkVpy+Bawe
MC/rGWPemHdbmF2Ao0wFaPpip5MlOJCK1HDU2sXMiZ6sluoXTlRcLykd2gnHrN03O+LJ5LvN9nLs
YkTOWOng4cI5S7qzxlv8XN1TZheeAvFnU444bXv0LiQHSoqM8BcD1fsgaKKAjLCipVGjdyGhrISv
OaK3qI7NzQUEm6IbvfGYBFa5wT8WymtsuoBLosVjQrKUCEK5QrmAYk2bvaG1bmmbc0cM7FcSExtp
SCaf2zxWpEh3TsyD9hy48La6jnrLSBOUm+T7+z2Ubkg3tMSCUsVwLxvllBSJFasieWDmbg1bXE8r
arDPFTO+QdtFWWL/tg7cDj93gUqDWTNwDvR7hMxZu1mpDdMEATUQ/a46P3/LLIpwvMysy5Pd1wrC
ZU8LlKHR/KdWS7ACvNzErHEFsXYCcPDomes8Wq3PlXhCyslAu0qVE1ptQsmwVdYBAdx5CpqvVc3m
CWIT2y36J0PNDCRtqwK7qTx6LpZaYiGsTZPdYgBZv9S+5/bI03VX2yiXi86TMi+TPKFncw4zejYf
CojMq14SsvJWR3YUN2tB0yYuH411qRGDnRlqSFGUIWMlZEiH5m52O16Je4KLMgXVg1xSfektsoXh
Cx/j6+OCNGVBNacAtPp+xlGj1JEKwLtntoJgt2UJjFPoKnuInLvNIYRlbqgsMAJwmZBacM/mDHNG
qsNpC48bMMIqo+RfESPIa1C8l+wMqJBeE9RWP13OkneJbyo7mNZqzOWnCXzJw6klwN1jD7Nc5thL
HeDY0WiJ1uvXvo3RC9HY5g+F+i+Bi2XQNZDcwnCbIsuM2GKj3L23wCCpZ7L2UP2vIVTjeikJR3Rl
JxzAGbo2uJ2gb8wGJ0aox3jAiAHrhXnp1jeTiFQbtDsnWj+M2nhsHWw71acUKP/B29YuiZMLDVET
M7g4uUBI1U/b2TIcjA3knlvgT2TFl61rRf3ugG99q0Q7oGS2rZkaZpB6c+3+lzQ2ZzGWX9233dGh
e07jK90A4vG/FcmuyQcWfV5LVSLeEPLbXZMw4zfiAH4zw4j8D0yg5QLkGhJHSXZEmx5Gja9niAi6
8Thq3sVojine39q/JZJcs/e7uc9X1eIcc5dlUlrAoHL9ruRm+9bGOAdGKm3b/XAeHB5T8ZFnjjXc
Y6FgdZG2JWYjDggfzC40+MHa8cV9YLnHtH0DoeLXbenve/b6zeyTRgl1p1BMgbKrF/QRpGRhSRD5
4L4t88iC6gLPjFR+sM9EQJsndEgaSTLobGE5lZeOA2FMBiVWHF0gfYyXYqKFtiowgVknDHijtbQK
MFrH8XpYHqWnwSvBtOFaqVUFwUq12f6iL5irLFEKMgcVkbWTEer0BQuUxCWHfKbhhO3Pbel3NAN+
OZ+2xtbjiAd+GaktEvZutm23ZjShbwDRr3Zo++5WRBia6GyLAUiOI5WG7Xt/ivXVdYpZ5tM8q4Tk
axs3OoZfpkUjA527rKWir9zCtxwZqu1BGKAgFtbPTmJ3yAUh/AQYhHp3pJLnrOiRzZKyndhlPf50
ioofbiqRBKeEFgz5J7Ma9IvgfbqI/tA9Ng7UaYgPrckls4aN191175HAHt2wPcWS8mV6e1xOlbBj
RYdZ2yT6PoCBmZsL6+DuIBM2aSGVxFPs79aox1UzZqMjO8+2DEa2CFNGmc6ViOlHgCsUR4Rh7Rmm
Be8ynOxH5L3K340Lpdi3EfGgGnKgKylfQ3Ew7HGcWKs6ukp/xw8VJJkgMctx48LfUV7JKwhlVdHZ
GPNSO/gm1nnq+P+UBqNTJQ+HYjpWZU5F6gUPD01APrRxvtd9YfmIEoeoCQaRo6EnHxcXUXBSFPND
4ofUV+eXHe5FIHGU8bxGQeJce7PFvB8hCuKEpKK2HzYGM8dgBhmywX+uXplGxK4GoD4xI4lfM1fF
5G1WsMdLRqBw8XOI2GP1Mz9qa3G1crT7Pb5GbTxfmMdXd6Kcc4f2JaqKsTGFL0UxzMuSLBS8VMvX
V29uu0CqYyKq9UBglLjtGulcWSJXY1upeLXKW+nPzzEOnHA/6YPzfGwh6EDKOX+k8uq8Qkty4oDI
StxUjEKtuy0lVckwMXwdXhd1Ne8XaXqWfF3GywnuW/PqFeGfgkJM4GlEw4d2y76Dcnhhq0ZR/+Rh
kZGO1V3ELd0I4Oc2hk1rWJKGHuUDMF404hL4j0514hm/Ojow6YU+BI9gfpStGAkdypKyfmi/UIwJ
3JRHqdxNkFYNL87om5pEclndq1vfXAudRDqNr4exHX920T6MlVh5h7yBdlSWiRtYIICM8gyvFB2i
rOtkJ/3LsvlDHSJCoKO74zdm0Fd/P3iMrHjNH/VsZ8pnVty5y7ncm8ZsY6Fwdtxly6dQSaSdiNGC
Vvkd9XxRdwSOWw43iRh7J2di6f848xwPtLdhayBHa7Ahi9kAAzh9Aj105tbS9XKJA3deYOjitBrP
Ob/YifmtyDvWFhJ6RBd2R59lJGfa9g9xXtD7waNQ7wyuDI7tp2HYdOm2xnPPmKAA8py3W5GM8K3g
euLG30zWo1cjDjy7Bb2Htj3RBBLXx07Lq8EyhkMOf0ZpFp0dyPqkrtMxQTFltfBbWNCmoBOY/Ftj
/zPMY97g/RSem14wyU2E/4kazarRfGvtTjT7BNCmv2pH6vGo3GviZxdWDGQgMXuV39dnpcKjSDRW
36Y0HYz4GYyoL+4JHJ78jnCjwdjshw5w/bLGGwH7hLUM6dNzbJWydsGV3Iwu8VdIS6+SdeFw7WOF
eAepHNeSYDLd1d6CWcBWmX/qDyluaUNAcZDaUXuEE8M8g55AooQJKKTwQHS8KxZxPp6LTg9kpG0B
k/LMmZn5Un7aTXeWf69q+JqgKzBHOEbKTv+qSbACF2+wPqTpG0fSRzx0qeh1iiVbSg2GYrJeYglo
iMIYAvIblwlMl9a8x4AVwqWC4VnOEM8GhymriCoBkQyAAlcy1nTntZhnS5Iu5ityjNtr4go4wUFW
j7N0JBzGyhoTjJXQw8uG2obIUpIWboJDd0A+bwfKBu8GgX5XhbBx/f5OICJ8Dvdj0+nn6jG4N/35
8NNgkD9wTsd7pBTxiQ2yt/wvdVfYrLayqAxo83PgClEZQwZaUqvZuhJIOfPcXZ4L/DcGgKHwYvZ3
kZKxgsO0IDm9GzkdIHSyndx9p8Wsqi8qDDE7gD26a+7Zyjyop4iI2KqXZoQT0ZlQn0+RJx5JOiUr
688T97AUFYu/jk09+6xUFAmFs+sPWtjwCuvhPyQ1JZBMABVm3g5RSrqWCMyDyMcQCMGjWgGFOF94
Pi45n8yN8o7HUSWeziaucs8pjiYrmxAVe71eNeRXf+DCK82l8UlVkSu6UM4tFolaBgGkoE2QHPUE
dcOr8xFuFur6H+O44dGQLOgu+GOwBRX5k4YCALEaRCSSfM6yw8K+2S652JS5wlGrVhJsEyYVTFjJ
8Yb3vzPpYQlgoKf3pYn9XiTyLWGKEUnNGTfcjXL27dXJhAZAtLKteTinB3spWT2+ZSzzd0OwHRuH
eWhazpsiB/49gFWK+M+5IYfOMq0on1MtOQaXk2PawJF78imAblOVJwjd7ySDtK7wltyunsDUU0+F
2hnwOXKWnezqZWiEPb+KKjcXeuKwueN9ahn1ivQc6JK/5pzdmalfy0hqyUbNGLF2SgLgQuUvZXMg
ZFVxCtrxeA6o6IVwLMghplkeWi2cajTluO1MjYmEi/dbaqvxbS11M3Md7/ow0+32/i4rQ73ph5XB
l2b7QzcQCTmUnH000czU7rbDc0AYNLPnKNUN8xb4f6IFpzcMC3PeaCJJnVnmGNzBilCKiUEYgi/s
17JKLhTKgO/lI7cJHidngK4elNnF+yYodQ8AIAlhqYiLQ3ya3F/Ns9lj0oZx8Y11deUHIw/Fz/Lt
BQt49+0w5ydyF17RxQgmMhGQTb8rN25k01nD6z6lMqmbDdCwBC4chVxIOwGXDt2PfTcqoqbEzm/7
ttYIvxMQKXS+NyqGdEBz2o8ly/i8jreoah5Rli9Sxuj3OhQEIseANZqPS+PuB+yys1VcYlKUbIL6
KpPIg9g6CBQOU5yyOhDxhJu/TOKk0mI5fiXMFtFtyXh0NO1gla1Pd5YMZC9nDWHwWz8BrTC6V5jE
/1C6bjP8MN6rR0gjnULvIsKS2ikUPJA6tTp2i/Cwy2wKJdN2Dx7/OYBIGx/aRExQowjOdhY8aeIe
dPgC5ZuL3UbkrGEzwbjMlbpQzGPOcocqW4VqiMiFfx4zqJh6HW5AmuWn8MBLvAFE/2DMiHIi9WWb
3q8XjEmS/fMfBoeDMJuQMxCbEwXtb849wdJusRgbKaIN5h3S+hm+ytJsOW65Aj/bhe+LySnMXpzx
UE4XP2fI6ETHiWvLQPAR/EnVZC7XUN4lirJbCRDCGg07qxT3pruo9cfmjmEnTwKyu9riSDyawgEw
5H+dysg4Cr38GDAmWB/n6h7SRPG+KVICBPmsQ7dLEfUmy429ejVWDbnmrigRCt6g0IaEEy9jN/hI
dGRgBEGz4Cm6sc8axca4yF8g0iDBbw50NBfEBdls7h8Q5xgqugAXelXFg29+3Eq+kjDKUSxY7SG8
ZTAF4aLSa9y/FOzFdoWNcfkgZ0XAByxnbFm/RZ1eK4APDDE62RgaxYUYRZHZN1j/4ljMGXozJUMY
A+7KVGb1RrW1xtbNVV+iQ5Z2RIrKWd6jyerBsFBa4PuBJjVzM19JfosEwywGjH2ersp5cc9i06m+
3BKayYKdWJEwFrTGqDy7P66v4s4JdzF/67eiTajTGDtw7ZEEi9pNFGGPRZWCFqDElKTArdU10ez1
havbkLozPN+8cDYJji8OvAyq5jiU+/ZkRxMEAzs8piybypQAO+34DwCSwmaxAMQKNUHVEVXYnPIh
uHmi3At/nI+wQoMMo/rlXUFEh6tJ4vTXvTNdRxvBbsw6+jR7ABYtoNQyzonkvrVsjUITo3QOYKW9
Z67yLfiMxcNSNAVp3HPn1O2p5dVU5jF/uE2VgETt9mDvgzoVRkXetbrx5FcezGHd2I5x/0K4woVz
waFvCAc42rUcZGx40nbaX/u9BoU0jtxHiKqu1AedPsPXgMeOR6IpbDW/Fgp0iE7KUFDO2UBshwau
AOqiQDlLveno6uBZ7B+KCyKjn/+BIRVjW+KXTHqAXfdduUp4twYXM/3Y4jiSC70648FZN/QSidAW
LWiteoPbWcJwp3VGKpcxWD7nkARBLzMgvZb3HEkT9XH+ZOctXiwXQ6DFOkV6esbB6waXz218uer1
PTSPA2UrfaReOvi5HtoqwHot4fUnAEBd5SjAEgUU5FxBc9NmSSetO/SxYb0qvbqPo92l2gcrK2Bv
dFUSPY08v5n5XdyMwN8a3TH055ZkxhPY5qDc4//AxY2Q6dKPs3msLlrzBgU+a/zLmpsWreLkTZj+
38p6gI8JlVuOozoAiuonn2tssTzpUJ6OEvpnxsJNxPiQKwYHC7pD6pnaRACLvlBYKo0OEEo0taeF
ne9JUMPirEyVNLI9mdT9yn7h/yq0X9WjT1KyVrpUZIGm/paq2PXiXRJ8WAlb0SywIpr06w5N3I4K
tfUnZt62A4qecNj0zpyTJSQTVdspc+8v94v4pB7z//dpqr3arVG1WcJcLfHhbshpljYTYfeMtSHy
74yKlKk4U0Hu0UAXaLzK+9YxFB866o6yQmE1786tF8JXaYtIlhJzQ8gG34ejsBJN4vXQdBRQRd+B
6yyIVydf4Bq+6kFgE+tu/ADbE/QvsXOatGeCVXlhRkSDIWW7WI/VtUGnE/mEj+MNnD6REU+zGySO
BbFLd+42MIlhB49Bz2c1V6IqNqlkApXyvBKto2k74LTLF2I8wWo9Y1KY1isVulOMdpHPTYie7DrO
vIaBKIbpftgnQonfSIZWnTootBxQsb3ZyVQdYT/5LEQ1k0K2s/7ls7eh6uW6Z79njLDwdRrqUBTL
i19QotbQTL047t3wS5GBjDXbWofIgDsyr2nSzmMDRUVoCkLemGoh16o98G2VJ82e57XM+vbA1TDv
LjcOcURE+RiXH2QLKV+0S9Hz3rrZnIbkgSIVEhKgHtyYxvlayrg9V7JPfXkD+rJwsT9PoE9ADZt1
nya3Tiy7mKMp3oZjL0yclcWxjQbpHpWOOiSHLEaxXae0CHxzXuLJ+C8nX2wrD/N1PoPGZMYnsZlG
17mx/92StF0awXP+ToP7JA9wZ2/9JYlokgKwekUxb6nW96ynOS6j4qn/WIgHmuouyjOKHbiNCEIi
BQZCETmgzDn6BmHshgFPiuX5Fyri37F+Ltzd815o/pA32RuPSKHe06z5BRLZoHnSTKPvq+BGWrmA
R+hJN3RqipVQ1QjVuUIbkgTMm6wOt/rSUtDezc3HS/jQw9J5U6Dh2XAo+sL2O0lUgeSso/cxTiBp
0paSzj/Ni+ZY7Wu17aKAhZ4K0mX1hCjsAcPAwIiECDBgClArC1WrHjB44wets4iXCjV3Ylna35WY
dE+m00u5ryt7tK1nVrL2gZyX/Z1Rv7lBteMWDCHG30VEPcMNYo38INHa2oA/YXIZQB7HjEHwAXMm
vZEaWsLBY2tj1gwJpEtK9RZ+qmlsDlIuzmVLq/6ZKiaSOs3LdZw40LOf4fvABRaY7BxMV9me35Lw
up0ZgvlA43DPTru/3bmMPUEhhFA7a93BBqoME3tCyGGnF9TyM6deJQ61ynbWnvXd33WKRdJ7qxH5
KGKjDyZdaR2cvdC9EBhPdtqdFeIi5dK3fPHwAcFVpupZzkWovHg9E+x5dq1Km7jMdMTBwKBnv6PR
cfwSifi6tAIHrhdkAH/13MWbOzfXT+5w880pIHhVUQsYdZXnFdb+A/wKF61VET7kM+P4dpnWEOKA
u7f+jIcfR+O8HVSGEqTqy4NXO23unRHtnXVyL2nEG4v1bfn8QaICus1/wQ8osbcrMS1eq5PKVHvu
qebFR8B9nSintpvMwc3CdbNW8qBgPmnjTIoBAuQ8gu9K58ZGtvfJZo+vC+wr/v9kOXF+LLWHKBtT
Wbifwj/eGRSRoSQvqfNHxahs5bTwLwlvBKXNpz3pJ2YLyZEQfC2bkAgMLTOlTTYSD//aTZlYsuGv
nAv4895vILj4OKQrjQyWYeLmnXdrt2yD8G5znfjSqjEkmdxBmKP5tCPzEd3hoepYW/+E+WDyJpe4
SRJ2ahSAoIN07WPxa3NE5ajgfWmahy4pnO1h2nb9DXS194/qVIPQ/b8IYnC09ZRG12ZotcL5RJVU
jNGXdUexd+KN3m+QTOBUvrPmmFKL0/onL8ZE/AaiGco6HnEWBkRrrkTPR1HgPXVhiIVlA+qCsPMx
8v+RgvmFgFS4YH9hbrDDhmJC0Gvfv+T5Zzk//M0N0iJVlPUyWe1wlfOndx6ySpxFW325y/QONfiX
vXrwz6wcHYpxhmxB/G98UIH9rTy5nOC6wWtubuj2waIx+pJOU6aTqG5K6luXqh1jBzm5uPuaXOHc
0RlCeOx+oB5trL2fouJq2xwo2qDTnjaznGE/H9cC9y+nsJlJWyvob3wcTff6yBhwoC+3Y+eHIS6Y
mKb55k0X8ugQHzu64ltpbq6B7nNrys6ppOAvax79idAmd9Ytanu1pev+JsKCsPeDrTbYwBf1Ed4n
2/b0Hqtk7mbtFm4FtaEHmgPOZf7kCFv2dJm+mpRax+w5rLCniknWAI6hHreCm+9Fwp9VgFM/1nF+
J9jbUgBq9tI3o0Y0swah98FCLw6cKXpsLlPRMHB2U4fP5sAD2wegNroRo/QrC7ofxz7vTyowZJSS
AFTN2gX9wnGzq/e1A0HfrhJmRIIQI1y9z/OOJG28s1yZ7MdKq89TJh0/6JhtomyRFBNdgvK6+Z8p
RVOQQfn2tDUH6OIzVO5J9/u2bvQ7Gg4URxlHAeMhlT89QRTj7/yofn2tf4PLg3ywJk3aLiJ+v3AW
zZNTUjp+/QsUAaBH37UrdQjxMLINTJeR8enAp08qgBK5kMCmzy6kPobGd57FdHD+06tteVHjI7uz
DaRiECVhSpj1L2n7O5YVplBHTts1xWAEp5qttKyg3EE1deaKbu6l0khjjItMI1gnccj53sW6PvFH
RAc8Ee2xSVhuohSz6LTIciMh0thzjEfwBamsDXibD3AfdqfZup5pEwZOuFP6cfYxIgIEDq5tOOSX
VNONnUtTzcRVzIsnl+lfwDAcpuKk9d35yjeOY30beqq7brX7pxeobdxRIsSGquZGE1tgLdOfz7Y1
HPKg3vILoXk6LUsSPHyyMERS4OWPnHfMy9gMxG2gqWHiAmwGEq3K0k/wtRjjZqEFUc/CHAJulyuZ
4kGmDT6tX/Nyl9Ei8tg74h2bYeLYyjOpHcI8CQK/xUHMhftqJRyZYxZ0jXslrPxMRyuFx54TyxCo
zhqqQRN+f9achc6eOjBTvjCOAwbuP24nYRBxv1MdebhZ3gKzFI/xNjGx00ZhvsbsftCMjTUpMV6S
wvGiUxsh67v+KMhY/KFbmgxqVtARKs6mMvXmBZH8P6MJ1AoBEvkvvBkE+cSj3D/WF+LQrnTsKTJK
q6GnONh3HbB17MvXDTNb+SfrBSaGEJDKdpK6cEqwx4hll9cCHNgoSIBYyx1g9UokdXiisXq71HlA
Lyv/seXgC++nj5HuOtuQ4nKkIHSfKEVijo38gIQlC8MJt0EZ+0Ahzes1CyBv4mOktpnZrt4hJEjx
NEgQOkM/gPamKb4AbF2C8MUnyG1uE2IjpoIoXGP0jBwO5S7PCLvgwk+dvGKcNh4XVWFOhHB2FGwP
joSp+4EzR3+4JXnEzWOCH4SvfReR/UjA7I539ujyJlKkSklBLwZIq+W3FP7EbtJn1YGt/OqEb5Ds
RMz8vg1uStfg0Q7rvcWdczXwBtnVDALj4MbRgQmUjYbERLpwtfvFe9NzgwpOvP06iQf9DyYCNvl4
71hjGqjxrSDlcCtENCb85/uvzJGvm2+Y6VyD+B/MT+6Jzp51KqGcx5G1+QknOA8RYHhBngjpemj8
jNxUJXwZUoVzD1Zbxq3JL9DXUjPsKA2me1t3zlQhwrW6jEFqW9ryfwqtPDQOTbqSSf3HHQvBomVN
nvV1hvQBvPxdlnMaMTMvLxtOfjwPG4oS/6viCss0MWlj3TUfAIT7zFbu9UgHNoUs5Pw/t96LGkCp
FYyaxPKMYSnQBTT4FxpQk0PKlyiXpRH26vDgZDuscGAaxaJJSIdyEd7gTC3332bFDjcgfCoULmi5
OSQsH0ceuN7ZhkEsB1//iyOIHTO4HFBQ1ZpqGrYNnDiJDRFwgU44FjCXyyGJ3yCwEycYlZpwue4D
AgrfAgrrj9dq5Z+4v9qYiBuupHv1j9Bf/9vTBMXTE4dfnLTuMCarWRUMT17CtIEppWNwWEliRcYg
xw4OvdYRWWqyLWEzPkwUQsjUDZ/6/pDhRRaGrE4An1tLPvNqi6mnrRWO95gy64xEguSwVudFu+eF
5MP5eZ6vpfqUwjnxapTaVTvjEl73d26053uqgaL07u7zGWICV5wP+zP9hC98pEFH86lSeCTqnBCn
6GJ8RWTCdHuoRzQB5XpS2mRe/aQJ3RsNZKOmqkyTTk1R/isIwVKCz0MPv9YHDOU3/L/3nYIETXRb
paKZim63samvGAIadQYU3hLQO8TCmnpykmPQ8Eyzgu1eGjmqevg8Wzpag4d9IpmFgt5bsOv6vjpe
N0qEOzvOpZHlmYErPh+bsvLEbj8k1Rz7Hs1JbVpdseyxFC/HbSDlXIv+FqElcoN5hCl16+o5wbtF
CK+qb0VpcQnp9rxf/1QRTCbNx3njCIp/fwhtE1RopZsiKU1aWGgEYGzx00Hi9SfW5qtIT1YO3no4
zzmr9NxKGujgenfNgy/2aT3sPu1kyWCE34NwJAVDJoPx9oVB4nkx2IUvrhAkzu0Owe6GAdnW9+wr
aiptmStRJ1zyhunDYRCuWGc8QveHrGvBP3STnyL6U+cVHrlOcvZjwME8UibAtjDQHpqqQjexiW6t
NKXaX7zTN//IF2qjBABwi7vyj4rTVxWu5nLwwCYtZQjI7sGEUiQKqcTJq4TZ2EJdOgzD6dH5LBPS
HTrGK5Tf/+jbSxAyxbc2B8cwJYWqvV6LpI3qipmfLD8JY9pxEn+XaJP8TSANorfMo/5O5oVTHdAj
FQimV0gOEunwvA+trTr1kyeXCHKZT81bPpKkZM+rA8HknLSbkzX+p+ndLaBd6G/lqHrRqgQbW7+Y
LDENqJDlvhojID+p7v/OAB3KgXAdVGm83ZWi0dsYppTBKLVk5aIZjF0Qp+jfbMyD5NChlY/T2vdY
Z8ZwlbFGSg5I+eaqkIQZjMSmPAU1GxZwAcg0rAYn24f8dEgXvlAbq4kbwXkYCk3WAHqRRK9EwAAR
tMALADOsa2oOn/vcPdyQpqINSEsrrToeafeQnuishfozAbZx3ZVL2KaF/ngukApkC/HeAYwFpXsG
QlsddUYoI5ICn5p2/pSkQ8tpp01wxjiYRBRvVEo6P7CNHlOsSTw4N3c8/Pxr8esGNmMQYu71VhZM
EhPh47mEwLemlTszYQli+B4Q4qGPFKI/+cnoVQRfWupAMxtpJcCXQwb7b3HTVxP6Xuua8pBovmHU
AzCc8cH0a9i3ihe5prWpXfrV+5HcaPjg/73yBBJxQ+7hoxa0nU51nt1wslnjVAAjq13pNOkuyUM3
IWmGc3Vi+AqIJ4t41Du7pa6ASpk/dp2kOaC9yKXwwQ8UNg10lrMQYA/Ku9vc+caKK6JVZkz1zfCs
mpygErD1PvHd9o2JlwnjKnY30qTO+tZmQMLKdBCGwiBh38adRLJOh1x8hQyO3Be9ayDrp0WSolGF
k06mNlLUfzDi22ioiHQBU3TrqLiI4N+8DLIBJADx85PThRHR76d0LiIdXFlMyRP8gBYXpBQUHSCd
fqS2V4AyPtAKVfREa5x+dUwugVU9mHlwUz1RzlZWoMNfdbmGe/F10ZwB2MsQo+rzehyuJfXyZywk
LXUatSVRL2EGU+hGg72gZNycyx18WppOC7OIinQIG01rnOrUqEBF+QL000KmWRX+68d5uDuU3tHV
H9kz2Li1tCf2+LGCNntfmvFLQPwqY0S5w0bnTEQOLLmM1LBN8iw3W7dtoJeS3axaWbjKnAhC4D+/
BRKf6xisKFsLaY7jISBPKwDdOaLsCU4Nm1SFwG5GDWZ7Klq3Mhthvaf47j3HlOkI84263kSjliX4
sfg+MG6h2GaqFcVJn+kXzA6B1+nV3mKQ5FouH113OxvQXym3XPDwORel7oMkMhqbgjBevmCODGPp
bnFcAUGTzEW+AjEvx5crvNSAqBWbxe6O9iqhKTm4st4eu2yOecpRpT7e3uXE+TcKdaZEL2jQgyjM
zaw2fLXf1wDtCDctatTWzmdc4jU9WFCa2HpKfGaQp3Br59luz8zgb9r0Sgj5HW5Xp/peWxkeglpr
eVQ1DaeQJtl6QnHCuaK46uTbMAfHU8kTzFnOvPWE3fUnjmQWMOsdteqOkkF4pqdNGQ2+kRIbjkQT
aZ+LDMawL+ZsQBvypF7fHqTsopy4MSjVm7TJtjc2nlxkNe7d+RlT0kSbcMK7N0F/F6g+gfg92RO5
EXypSGwqcyU+Mbp5HauwxctxpoZY+hCpmCV20dz0exo5ToI8ZqBjHND0590tAG3Z4Mp1xy6oMNeY
ff5pulNQOxwfFOGfiIsglK13DynytsOw7IwECv/tWjfcDSJxKrl6uaRh4tM3AkuBr5sV1vbbeo1a
H9b0s+1XF417zMHCOKZm6cDqlqqj4FRQXz7/nXFY568EF+PPnkOfkpA5Kl+4q+fxQo4Hy5WdqT+m
HCngD8WnqlLNlJK00xuGnEoyOdgi7m43aVpRKMaHgeBLQq6TCeIjL0DJcbNSx8hnKSaoJcdLq3yN
DWWPwRZxQifwYe2G/bbc4hfNRfaEFTjSHnYwOafezC7ru0j3lJmYjCCEVH1FlvQKVsBsK6+TuRdL
O99g/L6Wc/7fUgbMXIZr1IxWmPM0zAZFZFgStt7O8zegCHqCbaKEhxcicmGfkVhS+k7OJ/GNiGZK
CawSEPVcR0Q/wqr0sqcr7GFTIwZZMFD4Ss2sIJqajjLiPzoXvgSc2M62aDqzvTzwTz+LPTAsXzR6
8jcpfam55rerFHDg8UQDHc7u0de9HY59iY8i3EPx0+Y1CYWfJ3efKzjgNrcOhbKmxeOWQkV1ZBrw
nqD1nY8bGUHnVSlUHEBGFwxVihDrwBTri3r/jwNwnDz1Ld50Nwmv18X3sEGzvjm59MGujLjpo+8A
0z7YjhgiA+MkLE582bWj1Rkd94o9XFq23ZQ9ya+rc3ouFSbUVPBWELWO6cjGr+1zlqc02eixsOpz
PiKLqR/RZm3NlNcN3E90ESlFxgazUAnJSVw5F+QYMOLLzvf2g1D3j0moC14XGsBlN1Bj4+CCdoIj
X/9D/5qv5DIf1SM68vVVhQDwrVOyVL2ggYgUx2u1ddx+ZNYkh/DNtVE26p8fKWoRSE01ZVMyUbTX
Qqx04vRs/U8j3LTeBp4fbm02xtAs7D/Pog122BfYnohihrmwyBRZ8oAhxfy1CuyhpNbZd29jlkn3
QI4BOZc2BYSSklsWduNot2a7CvuMZ/6e9w/jlZQF1Fj7Dj+G8GViqVGblmZJSAq5U+r2dCSKEXnX
fTNUgA8NyrJ9leeOBhxScTGz/VfDLvL9DdZbAQ4qvPACxjyjD2KeZ9CC7kljK1Eh5dFmuc5MQVGR
fMZSAvLnvTia9ziClgqNUGug450bLJGO48JtSuPnhPwRApinTd0sC/GUx9rcZ9KKYVMgm5N/+SZa
kG490WRo1cHvMyhhWvPvtSymN5Xgz8++/1kbfaKMUrqhr6CYfv0/0u97NU3kIRm9YBYc3CiYq1y0
yB9rjFZyeK+99Z2/G/cIZupl0MtdaF8EEJVp2oszj8y6LOXEekjtXNeoWKe6XHhkGnbfZQToNA3F
MkMmPl/MoY5AdcgEla49vfjP6ndXgvPecCOVnERqvFZOzAwCz2s8ubW/qwC96xRZ89OfX9G8C9RW
KmYyUGvZFAoFpnatTDUoLVQTi5lGnCjuCjuTtmty5jkAX+2lzd0q6pGxdbkTQl93atx47Nxz1FhG
WoUYX5A6o1HUDAkKhFryqLGCuDH5JFijM5SWmHWmK5eW6MRMVUOKqgDgdQ7z0ZJFGhnzr6IYR6kO
K7d2bQXjKFZ6ZQQhz5x5d6Ja4flmrtcHgYuMk67pidiOKE06luT4JuVlQY2A5c965sG2WJ6DecII
WSh7HeLJUvJw9oyy7s63KhTDKq1d8a+7y61rCgO7sDQO9MdPQLjnJ3fMmtsRGEGyrve5NTf2ZDwZ
B09Wtvwcbf9gnMX+t0YEmTq+VWQAxXWTPdV5rLbSVxOFEApm9ADxIhr+o9deXP6oA9vGab51RjvR
scprzdHERSYhoCvDERzy8T4ZW3HRgbg+DnOQNQKl0uNjwamo9LIkyUBf7567Q7ZIrRBCHLawg8Mq
IsObRsyPD9dMFLw22SWxCIeAOmnHWzBEMlxv4SURrxgx+xa9lkQLmibjm36ZWzw1ozYd8WxNHZ/g
Ld01BsBtu4sD+r6Zk3hEp2BBMagECnUIQjZVdvpt7fiZ6Xag4D89DyGDkTW2XaX4cYtZ2Z4F50Gq
/adlsPcBg3unToc7koWXkb6mUaBf+qbc6TZixJDGamj9L+f2Wx/VrhkeFUrItvVzTuRmBaH7f3SI
IBPQvstkX53AysDmV0hNLBQ2jVQqW6R+VCZqu8VgXrLDOPkEG9cZkoL0KgI2qdTxuj9mLTiXZa46
BbLF+0zw4TINcls3fGMy9R9Ez0zxXXxOWPEKgw9B8GPRh7Hm519IXGQVfXxuWDocVI3xj3KLPjMA
BQOaA40TxA+O8Eab5D0bfnmdPlgJ38Nvzw1qjOOGURRdDYUoIMOEp4cxoIqhR2t07VhkB4GiEe/L
jTLKk1unVgYeb5wgZA/W0h2BNegFvpTN2/PSnKOYShs45ESrGbFCoxICEt2N6WSfhHyY+/+QjyP0
++mxtaRGZ0hHTv1HeBfFn070a4IcVNoLDNsVvASsuOFHurRSQVPpTfhTv6kVk8oNjT+SlXnr2IA/
nsi1S31/f2qqCbImQp3tOjTNbLFhxveKiOSSzkqCrehUkvN0AYHuobNpueeTfR0NemCgT6dcsV2H
lX2fzw5aYnB1W51XHhFgvvIIbB0qCC0qOen40UMTEIA2S6Ad+UnNtoPVDoo7USY5B6u8FSKVv/oX
KOIHX/DmF9It1S7A3JQVHGnt4wbXuusgsxe67E3yoYg7TnrHtKB45ow+PT452QcWqrPEUzE3WTFD
ofkgY1J9TYdbRGWV+y7ZQ6k+wJ81cUtxs4jrhRJ/kc+KsBdYmkkJ3H6I6f3qTibT9gSOGzn4Lu4M
QDwMmIg3kk1pO14Y366xMcw0N8JAwaKarafRM9gBZHOnNT0n4yNNE0pyolQzh/qxlmvX678p3SkB
VCpvWzwaZpv0oOxr5hWQwXfeTgr2YIQ+jBOOnjMBu4645obYv1BJ7I3OjELk5zq8h3OLrHwMYw4n
zIwXv7W5Uix1aaQ8AFWnUpULcYjSn9qQ8Gj6JMGn+XNz1agfGK2lRFd1R+Lr4rMqPKzN7ZItN25+
jKqbfT8cp60RCev2knj254YNsYYPOb4OrBHaoohesiiQ573A9g/LVJaKWEJjb6vSvsesHLbGdZXn
JWZ7mBUqxTNPLyoL52sa6UN2mDOo6zg1Ldz0TTOiT39JEhM5QGQ9C5UMkfus2Gnimyo+Fazx1JmA
+nnGgnBjBzV8QOY9JMGYVQ6Uc/PCLxijPijLKNrOSZbX4sqrzfDoSpRb026PXjKQcy94AZZLsNM1
jDEjjaIjBRY5CuWTT/txNXL2LGJ239Qu9tCXxHcwKYqR6QxPvDI0BSAnbBE0KwsHBmgjSCAqL8wE
zQ019rDbSNj0sJfR6dLd8gi2Ymg7BDGoUn3ENdQ/br2vxaX113U2sZmAnY4RL0xZOBIobhGDWtXZ
X67Ox3pDsYAQEDV48KjWt5HWAyQhyyD/FxvrZNKq1pAMDJCUwI2NfRxasr9GMirDBM0aYg4bUUl/
+tNYv7Y0J2ytRYiP/Oojh+Tr47d0Vu125Qgpd2TgHDp+qACYKAFBm6uvVJ98Go6MNl6tqNb3hk2f
Pe6MMBvXt7yEKxml+7axAnrW19uiqNX2iV/vB6G0iJGcZVcLGMxvKCniU4DoaZJMley8L0+7HTRZ
3YZtP+GqHe1y8ECYExriZbvSg6MXz8RV2vCM1aboUSCDvYnQzhrC44l/tFdTyIMcarEfU532j85e
7Ap9o+b5wwf/XdUB2GSphKhRCsv4zzEyPvE8/sUR7ZjBCBnyN0pqznKBV5C8CxbmZhoAIvxwOIyY
SL2FTPOTBYNq82BI7AOAJzm/42cRJL1pxXNiy2pmYLQIwcDyg4svaKxJLSKdfAw1Qljnsocs3Z+d
pmOX2nyhqCsf91OKQZdylV4nhmLIEApGgXzdRblMoPNNcvntutl5p4EBNeA9+4cRZY35S+dJs5Mh
99dQGFCAV4kLQJi5D32Xa5xYLDzIDUXZT5OJMaPv1MKNTJ14TRazK1F5fprpNEtu1wcYi1pmEjKK
TuwWHiJgxRpO9Dkk2PXIee3czW4BjrK4j1F4Ck7UoIExNNbg2nlKwYb5V6+k5VHw3czC2DR1lM95
tyb7apx4qpmBybFC9O48LP1FOX/THnhpJdqjNilCHjJw10nVkHz5UvHMqHFXp5/Qnv30BIDFfzja
HiRfTy2kyH9thKaFSYu5yNlPme0DSNW+4FX14vsoHCKUiF8xDo/5ir5zRZvoc7/klVVSaH3R3QSc
xB7okh/RUEv2Zr88gP/TqT/y5JQj0EUkAaRQgHGm2LRatDUFIo4Ujvg3MQQ6M9HMNI7tZQEB7kk5
E8CUHaPVuq7pV81voTGEST2t/HuhVIIOuHcO/NlgrOkBRxbafIuMmjw2XX+TO2dqbmyI+FXbVGPP
i9rjUnPa9t7D+CS+4OxVmZdMGI7+1TZXBp2UIkfvPaNhsQFP1R5SBSL+JFpkI5HbxIm//gA8xv+x
RpNGBJATZmR3xaKGs16tRicUQgxZVV/dHuLstcNh9NzIDMpjL83TuQysjicEMuAiyQSgWRhTo9Vd
1AU1wEAxhh8+kXnV6QDM/kYLNLkJnTHNIUC1QfuSLIPmGOrqEfWDW7giO7spACVpQESH4/XRrIfl
TuscZ+BKUE9Vr1lC+azRL3uALvvSFV7s2XHVRak2IHAOExzH7mKq2U62EaPOZ9C5UfbRSfFG+aF/
kMIbzm2ahx6gWpH2q/Uvv/KgVXB+ksMEimhX/gmjzwYXjRBzKa5vWY81NkbS049AbV6VxIbTEYlr
K8Lo8TI6xrisZLRrz2/tX09S5dC2g+pSV+XglrNajdD2gbPxnGaQIXUzsufj5dfUn+dUR6pseGA3
fmru/MjLeJMvFHFe3/+RKytVI9wRcn8xpl+DF94OLzQt82vqB+/DwOBn/aPiq9LqmOGtD6SB9Uh9
x2U8vzFgKD/zi5k3uYzwDsOfylqiQ9rciO8PPh/fXJZgy25HloZo7LI9lCek0/Lk2oey7FrKe2bq
cVP3e6qlMPr7nwRFW7gmygxy8Y90Q51CrCSF+n6Smu1eh09jwMiRJMu00EtSiNZH0N6FmqwRgHKq
3D6x+1QX2N0ki7mcZ/WmqOIiNSuIpfcJ6bMSdceFGQ6fgnF2BKHWTEKCRvnbE5hsf6sGd6tOcq5S
J5WmNsvn92VxB/aKdi+rcEEx6uGKsZ531KKnzWdcXGBTOFhSWuy0m9lAe2MlDDjjEaewbKZXlr6V
9Nxp2Y819RYkhOX+c3dVP98oyjp8OO8kUC01oJZneF4L6ttBnwhW/GyU1inbFHSTBP+KOlu2IN6P
pYPgb9mNLIf33o7+JnhIM2gCR/jvRUQdtzchfjEVm6W6IadgVl3Btf9/DRam+9OAijQk/Ht2Hpgc
VISdt1JL4On35EYml1sYFRTRLDll2pcLkQKBIsa4cfWUCAxBDQ1S/Etb6KVIG60r/vho97vAMWGi
SpMkm5mPC24aFd1+nZPtRv5zVGE3H2NL4AeYGVNeUwVZnFrTO1/jLEve6eoVt4KdbY00vbrlnxim
Yo8A+RhVhvZYBRG7rwYB6K698qjUGijlC2BscbzqYC64qzCwPktX8TVsfhW7tkKwjgcbcdfYvPzT
EfKPhEltu0mrOiIUWTJ3X/4MlOGCke3OAwkqCKgCl0ASaYVrSQh4tJ7jPr8wd6+jlV/u2Pz6xdzU
2RBLjdKrBQAAieC/Lgvh6bTNyyTxX/y4TtLiwWCulWAHKidhA6xAq29ADMB2UX2q01U7wKsFNcI7
LBKIColvEvunyMhUdBJGGy5QgbDlkUeZAg0YpDRh3+iS45VBzZfPDMmHAvWZUJsFqiJWWEnj3XPC
qZ653nn0CDt1i1aNKOAKw/5hTa0TVgAx7fTZpJJlPUPfxc4mBfUCe1KosJilhT4dmH8w3CJ5SKzU
haPaT9Z9kzUpigjZoZTdgD8MWPkcYxhG9b+B61x5dpIfzLQQvV1x5bIIoOXSPzEwXA7M5hjGBo4T
mV90jOhr0+rQmx6INXZSR6TsQi/SrPSOqT7ANMsKQcUcuW5aG6jRkuzDSma+N2YBK43pzUTi9zG1
SWbhyjv40tTpz49S26LMg/QKGzeCKzs2eaJYITplXs6FwYgesQDtTSP27YVjLEiHUycv/9M5kTRP
EHLCkZs60z8OsF/EG+7OB/WbXlyEqJbnvTkaKV54RqtdDnjdAQPXHNlxVQZ1VPxzjbWlCql4pwLZ
KJ++XVLoBh6W5bGHfNUFplEKtjTjfQWb7wsL+tuX6Ku7A7ZyLAab4/92z5qLmC9Q0Tj76GhQ23eD
lOZyiT1zQ/CRALBsq4/Ev1NhmiWOraK28+NXaExwyi8l28kIWVQuhykMQsObhF79x0aVK3ssKUAt
y0qJoj100JBtChNnc7Ypg9mMT4/uaar5anYeomNLFb0gA5OET9IEMGlNnqqBpestnvPoCbuKhnCU
UuUaT8LMlh3HN11ze8u3Ca79+mM9bJOKJZwlglvwGAjCtgIW9nAwu0w0bOlRJUfWLaRtK9Vj093p
cHn9TYoKZz2f/dtrCunS8QGtbx8C7+kfDDlVsYLk/ns2iPKVm2UXL0gou2fEW0jOgawxoWpDusCD
ywv5lELhPj2L/v/BaWqyWuOPC5NuJ9/06f+q50iDZlSJyhFeby9O4yYkCEPQDv9IAGsFDoTB0itQ
7iz22mUyCXqCZ/57faLOpX3oDOBWtaflGRCSJl7TZMY6B8ENCCWxIOtJ3XsFNViRysq5hmLzzObD
HEBp+MjwT1bPLJDM3Hx9u5QYt1o/vLmD1onqZi7enGaoY+erAuKog0oVtpp5FcpvmLu9nkIonHgQ
f+4DeWTzc4HAzmIrDUGe5HUMKy6yKz1LUBmxRxjBbrPvNaQNsWcTzlz93hwAvJjQsEX7E95KCj0D
ZmIiAMOUs+ANRRVrSzHCxlNiTXovyg6VzlD5kyS37wlS2xTteF974A3bdxbjA0ePBFfpnugDYu7W
RrpyygE9fPb03jbZPWRI5gRJyF1M468XP+qKyNBCdjWMB0tyXoOHaIlXtt15OgTZw9ip4Gan9c+w
ZnYhWjAJMm/71gUSDCikGzNqVO4RV+ci8kUuaXFNkT77pNq2UTo8lcB2m29WwxYdagWhsZ4E8XJL
uTr9K4siV/ozA7XYH5Ji5yZHxEt1suYNozy8vjqcKi8Zwq+kDO7NApW6+czh2b6hjHJApjmgDNLA
nhXP7mSYdUmbEJqV/QGRW6hfqQ30uzDCxGAO3SCPowLW8M8Lu6a7s70nkAJnKxVMmS1X328ATUuK
lk7yDnqAPOVeSsMCHOR4QOR3yGWTUNsjLpd6fu1cp4sr33qpYllLesxzw4kqa6UdBP+xVJd1T312
9kSlsJHLijSm+CqMEaJUJ12nBi+MM81wrr/BFvSRC4s/NpoUfPYX4H07yINZ6DkLa/GltYPhWsc6
EBORbTrVti96kM04DOmYxJgRZJgi2mXbLv3JPA4jdBw348dhdEiQ+g5VqL4rn/aUB9xXAlxLsxts
2zXXLoREjuVEjFFG0ZhBEn7R4tnloIt6qjTSIQWPGYILyj3LZE8wQH5tzM3cccsW4z9QWMPMcbna
eQfYsqSSlBBwj7Ykm0k6bAhBVK8oXSjfIyE2SrPbgVR1K+ntDf051TrBWdTPX5LcsLljqqOtgLXz
TY/nBo3RSRVIjSQi71+m2jiTfbxxpu5RJhXZCjKXhpCvY+YyFVWQbVl+wUrcy8hdNFtoyJDXYLp4
u8Gwbi9dlnPCQJm8xwS8YDgFu+OcSGOb1ENJbAkgq7MMAuvJA1zh0ItbJPBL+BLRMwWil9UXm7Cn
l+RPr1RndczWO50CGAC74RthDmXTfrpWahb8H66l8XGyyYxwCo9cvkk9qpXx0Onu+kAbt1Wb73tM
Q4/9ujDO/17R6Nud1rFIJaLsezw6AHCIfCTc22i1cfp4XlRtJo0PHBRs/Ds7XaPZHn6CMOXF/2mz
weKFbrfO7jLmZQDCXaQp4tUECOns8IJwX2sBAx57r8r2AHt85UqBMPyGjRH/1pRgF78r0ycRlYbO
JL+JcaPxOtXd9unvCUOsZhCUQmxp9vA7JD2C8BvOpBo3YlvnQbSWxC2ZJhAD8JL10bskEk8UdSNK
fAH4x52sWrFbZFRTB8VS1cCTV5ITxWFV3XzyApz5HiNNG8xQ52Li3t9AFwsawVZQYlzjR5gKJLnu
gerLMufeY85mQmAXT3UZb0s0Q5hxiTncpzSc9raS+TL9lt8496h9o8OGGwww657w7NSVPVzQkI0G
hnM/zXWibQqUNQyHGxAtX4X8Ey77Fsb5u7P1X8tZL5D/DOFHBqU94WDhy+vkaiVvIAWHRYLz53jX
MU9EBQn9eJTkp/Vb2StcohFEfCAifDCoZIRHbv/CGVHULTZEMaSkCQkUHiY8HsgKOOEbVewDE7BR
1O6C0ElK6lgLRbl453JXTnlpCc/O+HV8hQC5f61vHR/B3FgEawSDV1+zEYTIYXCMWAi7W1qK59To
yeVWH3rGWknD757QqnD5d+qd5xOxYdEcLS3b209aSCP6eW0dDfkK1ZiVMU4jIWeWApg+5P0axunb
93FTFDaEFEU9ij7W2iwo54grRwtqp+fmNcn52iEi4Ife0tF5p3tHlESByJHz7EqEQPbIOjWMooOU
OMpDD7LJZh6/qypMbD/aLWIch4Gg1ZaDhUnZQ2MaxEV/iY+8td3IWkE01OpGMCRwlmw3Tyg3YQPM
Gp3fesqEv43PdAgUSWPRZCRVyqtWEdV899HPyXOerRk9s83b63QNVvC7zcd7F0rH/pIpR7zTm9Vg
t8rwWaNNd4RpamPUTSyJMr2c19aYv7F6beLyqnHmWWowOu1N/+/IS6Z3iDInJIgwoTCrHmDuJPqO
R2utvb+UnktZoQ2gTQYg5PuqwBzk8VDtfmGtHcVs8GqiYNaUUs2apuh72qsDuC+5SbAGO7DwrY8k
ppax6R4OYvw9mkyeZ97p/aqHze9b2XdY4MSHJArDqK+48QX9R9XnhUt6dDsVd/tiyG93F9rGFONr
XWkiMkQi4c6YvtQUKzp7W9vlnmMmuWaInh78/xvTjkbklbrDVS0R0AiZsJpcOX3ss+7O4l4DOtJi
0oPGb8Fo8bMhYtrhL2q3a8sbaV/0fAouwOse+i7p/y5q6OY26GeWI+WW4rhAv2L1+PeKRy6OxpqL
7ipmTL7A/QcrVKRHfTxQduSGqiBehQkDlxJTXutJ+0pVwIBu8fnjJ6sOiYiiQCNdZSLlw9Km1h6T
t+xYhOpR8o9sr3eLGbrXWo+HUoea/V5BivYzcDxY+wrjP9oDCosACKVy8w40PFBnaEbzX91o0zE0
I+tV4M9GOMJC6NKjN4XRXaYIyulN0R8GEQpSjuyVSmzt8uTUMYKSl9FhdliQThLCg7x3knawSgc/
UKNOk143nLsgoEWVpK/K+cNyC+N2PjdWijB13ZKHjSVh0HsI87WejgKBJgwtNXzztwWSg4y8TRza
lglIghUkSqPrmagfnzSJMF6ao3rjAnc/+elwgwiwzlK9VexP6U5g4fuEeU9mAUsV5FyiYFWTYi41
XXdl0TyBcDN3KPYpcOedlp2Q1fuBFaWPhN9s2tSwwNKsG3SwscyV5FqxMRJvY5Q1RRcVSJ77PkQ4
aAJVm0WTA4XA/zf+vrO1a77lxkPPrhBvzqLNjzi7CfVWs7KGMEB69qZWiLpu6DoO01pz4XPv7ajc
Ro3AW5pc2nDQFCZsYHxXyIbHdIQAlKmnkMppx+OQa2unGVhJkCTgCGBJ7E00Ebm6a2UvifENdxVW
FPJV3Qbr2P0W5A/duPfzf1ffAfh9QIQdDqO0VmnMnKtDcac/2FmmrTPz85GN3VgZKdDPcP5uy0FE
/avw91nb7vBgGrHhwUhNfDghTwCkVXi5PUNTKP5/yYmuj2sLq5DryRkbwvUVIplsJAKjacjvmSFp
owbtz43YidwzbdS0pr5sztLeACaUj2HfgC5h9yb1QXpuWOjzHJUnp1hRc1FfH22q2NOnC8+MmJpj
VFHzPo9JP1jUlX4RxXcb4Pva8fZO4ZUOhmPMbh4x7ekrav3UgvuNSlm5vptlB3kqKSh2olxkbr7x
R5ll1y9Jl1vutwHK9KORQ+7pxDdCciOxMex5N/XcfuBadqDCt4SroeYP8N5EKFJC59qsCQ10jVs8
2rhhygThmY5vQ11v4MYbcuU/UnnnO8pCRrUQs7C1e6dsoawKoOCErtnmt1vohMJq6K4xrJK8uVno
sZ9KvgIJX+LkwMNCuI5QK7toYF8se3Qle9zK/lk1ZEdwtYvqzSy/+7gANvZRmco8KhuG0DotRyGU
HhCH/kHeqHlReRyiQwUGxjxveRSqkBcH7Oj+zpM+syA8P4eptr1re9UzjIV7oBXJ7vm7AcE6S6g3
2h2M/nMLvA955NqQLNZz4r7SMDkM4OGjClsk+jxA28i7Tuv3Jh1y97Hhojpg9TpICxxti7Yz3GlU
ECN4L9K9lLRqSIn34gRWKnfB0caezFOmPbh+VKuqt24EDJkOTSGHJ2AT0h0mmfnJ9bFowMiu8Dv2
QXkCzctMYdavZ+M1neD+G/bbJvUcDvEtR5FlayfyfYlq2Z0p+5vd+OUSmgB0NBJx7/gsly6HY+uk
2lQLuyZnx5pPzeCn0GwoR9/cI0pVtgcE8EvQHy46zWH8e85qt1FqBEqayLNRtGUsYg/dSJp6Q5Cn
kW0x1S3Shwfu/JExFZsPI6THchYm31GSGzi2/HGoBCRYRmo0w7PPxVxo4xHYuAq368CmHqZJgeL5
s3FpVXe7rPKAmXCjKB8irYlMmfErou/SfE+VEoBZPW6rI5+yGhdh7ZAM7S6ijClCBOZ8GY0Kpv2H
AT+nYLztNRe/VYVHtgsOivQcS6/KTw8hgMpseBpHRi2tOyW7AljFRUvO4Lnu4LTjXTpyMI7TddkG
U1vaMWuMe0zcDy0miMRfj64S94jbTWtJBxDRd/6hNiTsNgyLceh7jHYqAmSk99tLQWKRUe6hlkvo
wNT/cb0GgRKfWlILLT3vEOn23FTcDMnHVoPEwz3xbk0oAeXvr7PvE0qNjC7L7uuNJ/pIlGNOPnt3
m5ZKG1IS6hztnYY1EPyMrgsynn8Nhoe+p4FhAt0KCyrR++TLTNVLUg973kHZdOxNY2JtsbGALKZD
lAvfyFBLQ61TbcGPuG5I8K4vt4931sSCmiKJpNVsku25D/wz8KGZ4lwksyS7vhL/SbXKBOR0kdhF
4nKrPRTBKg9SI8qSrvPq47Aj9g6v2/5jVovDwE6Yu8/IAUGPIKniK1TLa19Xv+z4ubMO5Sxg3cSG
maZY6N1P3GCPKZQ6TjCaZ+ALjg03yBye+JiG1mrN2CHpFcpuZ2S/m4ky60aA9cM+SluFyGRdAt3m
F3pF9Q8fawINSUO3ayiFoNz9f9W+kLP8+GNw5+DJXMXhHfD+8DnHHY0FAex0eZZkNNiKqiGhw3xf
lyZt7vTCxq1XnszPvT+6zsDAzyEtJFDxwQdv1wIbrZFUAmMoIixDBRqz6hSOAFpsR5iAHfDuTUMp
HQOXs4hNChfYN0wAuQtoiR3AfarJSHVFkG2TfXifYgCD+kOx6sUPc9pokob7zNXc491PAr0OxnHc
inlqZYPhtnDXMr++pPphmCMO8TVaAa7aVNYrfMcTuSLrO1AlwWZhudhCcwdf+sIql7PaiJTTVpf6
IEjG1cD0OwAr0dhBVPnWroQCvXGvqiTezr8eKYV6Q9tR2jsfMmdOLYgtWL4cTVXDKswvoV14/w8B
qBYSldOppWo0KJnpn2FBU01KuJHXfzveMqlBjsyD0VGQn2RPZT9gLzynRfBb8n7egkHfyIzpEhS2
b2DmuKPTDWSyYatKQiH37R13yVaunUfNP1q9fVcfdH8zb72CQmc2T9yPCMegH1AMbHZLGkKLF5fL
ZrbBfmg6nv9XDK3SBpZNFKaBMTmpRSpYdUWR8dSPyDS3T2gqztp/TfHklkUa36L0LOgEMiqv1ji8
079uN1xgyxK45yFPas5z6HX1Jlx+2+oh7C4WLsSXVgfUuiWt0Kncc92gqYaNny1iBnx9kNLKKebW
2YwQrLaY1ccXTSQsCfE+bNJ3TmspdoG5v/NFX5ngVd7F4D5hmgqLkabtpIyWtBfKw3GSHZy16nt4
94sdMbkgXMxGogeZKMSw5pMuRi/qNk29FHLKhYSon+r29g34ypoGyB6+OFmEQqGYhRSCYB36f5du
PkPucpGZrFRDuvC0gcwNzUTbML7tYcw/6r0rPSJGgOsLPYB5jFjL+lzrHtCguo2r5UVQs0iJhgK6
vU7FbDjMWyADUhYgXb96F5wd8lwaM5pBXlKlz5S0Nr0dE0JLHGaQQbx3X3ddLfz0yGWfL14g0DKZ
IdaXB2JI9q4Wt7sONkBlYEI/EN6A7lfu4C/tAZHipLiFoRhd86UPr7JfCaIdc9ocezxVQLylymqn
uG4VdCguAaM4oFTgvdOBG4M2N3u1KP01Ksf25SCJlSSsqUTCFBcBNPBgb/dyi1JecY9ug2gMJW7F
dFHs7JFOIfmEy3reOZBe/utQQHXomMG0ipCSs1Zr4Kn2Hy7j2uc9Q8Npcjd4v/5meZnVK/LHjnEO
gNywNUgwg31z5OWiVwpnYooIltcq5O95PJYeP27QcwHgeICrRb4V08w2QyBd4nFsIWw/qWmpFtGQ
tHfGPpOSZq04fClwK0IfHPd1GubPcDAsiE8Bzo53+x9+jkwXfm2I1TWvSCAsNb9lvTGVC2wA/V1L
6T3Ah7uwj/veHxwXlaLOh0srF2SO8I4A+11GHlgJq4Zt+nloA4PGs5Cjv+lthAan9Q+MhSB04sUN
JeRgTyPgnz+Xdb0XynhzAagJTJdbhMhxDK0Ol2O3gVfJmJP7/WRnU/71ABfiAr4kTdAg82Z+ntJs
QL0R9ytFwt7VWLPLKhRT4nMsJvV4kRa4iCZ6Sr9l5b0YM2u5BeSXhOAp9t5EhtVEdeFwMiiX4bNU
WaZTRp8R3AFvJzw9K4Itm8VGRoq9Rqhh3YDsGvAIBvLK2a82TJp8h8Q1hLQVudlptK7FjdoGpTWl
Vf9FnSo5aopiEhqBtDee9mAMCHj0wJRhsFbUei0APDrsgJf5CW4fgbZmyhrcyEmT3M85+uTeWC/Q
rXC21xYTSy2B10mAdV1Y5SneBSJag3udHbqJn8HLQHEpVgxqBXQH/m7TaJrsm9w9czHbpoqcfJ6t
ZmqyNlBST8CwSfyxTW+ZMXdvXKgPyOfqndkza11lHV8DHaaEEC07j47/E+z39WIMTbg+hoIZiRaN
IPMzVdQrPs0csPMPYOULsHbT/3AzV+3zkXg8BN3G8vD2FD3CvcPS2fkW1UoGxqcJIrAUoAULSyWq
+B2kMdLe/1yumVGvUcTH8dPpODdlC4IqPmoZ+s41BIS8LKg61ERTjI9cl20k62zWDmZRdhbIeb21
haGMGm04MGCX+JvFc2QvcSIY5kRPVQkI4czvUR9X+28d4X5ZWrJbYr+9fg6BY1OzUTe3Ks61BXuC
L/4vRAL7YUlhmDGiru4IuOYn5NRwWkNxtEH77W7uOEfBduep0unMh7khcjDpLgqX/59cBtbKPpU1
j/Y2XekwuIfTAGOQOJRD6fPfCSG7n0Fedx0+N3gvi1dPxBwD1iBDVhFGUCBRObQoopxV5p9X4bIQ
8POS2EfYOjuhqS9toCSOYEmThvJoiZ48hZo/1/vpHrWPCquxcjIEOtu3NvqJ1wq0HO+AejnZndZ+
VDgbJXaWRVez29mt5BzjX3TQYsMemPw+qah+OM0xgva2gEFWYE3qMsQFgiPyJs8AJK5SJtE0RJLA
adHI0IwhPpd9JD4B7jO0Ox3VJDlIdVsOIB28rzEc1g0k/rKcn8YTaFH+fF0Ap0MQceCqY2P9IUgv
fD9+FqB4MBpJGMxs8rDdAIeiLsXug0Ys3h7ShcfryIsRo6Cz9qIqasOzKRTC6djhTqvBzP4GDOX6
kPDnQXs4X/TMLHynTQVxQAMFuGh6EhZd7r35vLHUNOwnQiJBto3fJp63yjoppkloWvOaTkOYw7gw
Gd/4o8hgk6JcnjQOl2TnIhOZQfAZ2JEayorT8FYewoRjQIh5LUh73aeip1i2LvQa2tjvhp469a60
61+4iJ99jCi36slbB4cJTH/xKGOOfQMUHEhE3SHSOlNQU0pvEgsxk8LoHC8/0TpEVy/TYsbFx32F
2YmXTlV/Oj3XXgvt2ZPoS5PwvpA6MFlKmHoBs0b72zq8K86URZrxiBxQxJ0AQ4pRnECnqY2SPNhh
SNXn9kwVtJ5e7dfVjxZfXaR1KECOAWnTnAFtAraxVUTo//gjvpoc6avu7QZlw0CrjG22I6QxrVu/
BfSO9jF2KO43oIAXpzUWXUVQoqWEDTRUAwqTYObmhF1WeLPE5IMmKeAHP3GSJxcX3mN9kwNitMMj
Kq9uzz5T7pHdF9MGvcyvY21DnbpKAYQO0zcZfNhSw4NlY3OpufxuUtcHDlC+Kr0mbDtXGBZxuDQl
fYcbe8ubrEgT2jMskb17B2uUX6X4Z9DfcwANsKT7u6AVyViuaPf37WEHSpFhl5/L8oxfNPbziJVp
QbDp+J9SUAIamLg9Ig/7Ny/KHIczSEjEJM766w3NM3iMpOIAp/az1psCcE/7gY9p4sEhAQPjzg2A
qaKAygTFoAOXV5Hd+AFitypuQNBep7akUHc9FMLEE7+E03CACIUJE7rvaukEDQyx5qrnjgmz/KJS
bQu2cdvVli5MpglzOVNSoTU9uwaKEdJZ2dh/mLOoyfln7/PuWySPhon528H2+iikoMU0qMLD9+QU
OSG1YJwBFOztQpIsPwJJW/ntdPAH2ISYCQSOqpeQezhx/a4NZnRBfLZrCamVi7uXuxX49Zc7PXkr
A01wLFx/2oP4KP5qcIZsrTccVc5Wek9BfM0wt1Esk8RaXTh1NysuoEBr+sgxyk/8YIGsftekt8DZ
makZt7abg8Iy3ITlHOqu3Ih4K4tIqOJJ2gP94gZsRNxHyR4IPa4adG/Epxr2ofuZyHnTjzbNCHDE
lmBcrSIdVz5tXM4QITE08FSXPH2asTLSJnLB3JgBvIJju6e3IXcY6cWT6hcUwqmyFCMmQRguW9wJ
D2aROfZEcgWyOHQ+kKcFrnM9TShBG8i+j6auhA6jcNKwj070yPABCL+wS2cqd2gTPk3haPUDmfOw
tdVsZYZE617qCfAjkGqiitgTrudJoBa9Qeg2p4RY66fxUD1OSjYqO1w3D4M1wBDODA/9ObmCobf2
6KjTRFkDYeEL1K65UyFhKZ//LEQb/U/3+cNK9dZ0ryoAL2rECVkpseNFDKsIkV1KFBPoDZQftLDM
VCh7zo71+ayZraUQs42wJq3X93LbjzZymD9ewx3JIdLJYRV4tdr4U9gyLDPsqd+uS9/2VCDFLCSY
UeUxAjxsSNGvcMnkI6PgilCr+MNtEttYj9332Qw9A3/oEWhlxeasc44k8s0XSFTrEIUe89/wgDb0
AmgkxFI1I88A8HSWLtHFXSiQRKeZN0tR2Tk4FSzYyyRyNK5Z751irbHdy0fr9yOPEtntwtoefrSn
yuwtOf/+QmGQua27chjvaruF0hq2Qm9WuzuTmp48V6dsTUsHzIrwYvQYmwXI9RJ89psTaqSap30K
mDrQMf++cGmy2jCUCpMeAsrm/ALfhreNSGc1c+uDfyS4GGdR6ogMrYS2dXeHqcT5KlJRhWvByCWk
cvf7L1nQzJfXShvyoJjmXWhBFWuwHA/MhTHMP4dd5j1vYFrKa7PDIWzRrI4P8VPnwWMdtehNWK7U
mwYfR9ozKqy0B1nqR40lMKMgq/8kirEKQlhG77WjADtVt+ptSL1J6IRtQiyldOejciEVgQLeSaaW
owYoU9QGWVDuvUZ9KIlmgAZVCrjtBTHZxfByk8wvHiFMETn8znx4iX+FLWSkfPBedzeTOZk+e6y5
qE4eI2n74rTDQKjM25B+kW2AB+a0Zqv6uNWeNLSl8eipCjS3Gyugg1PkTkhTHSsixsyCf6+Lxp/S
c8pIXQh5JLznG6Ge/iisBn0SWWxMCi74bjo5bLc6BzvANQWWPoZYz1Rseo0TE5CMqsmz3/GhbTwB
haakRaFI00SF1LBF81k1lsbsm2L4O+bxvlrhK6TCe4R04ZjLbX3Woj6IqdcDr3Vm+CmVLqGQxt4X
fV0Ory4hKY0FP4ON8QaiYVK8i9GS+/i8DuWFuIygOY6SSsZuDuONjB3r6CEzDHglhPJCIh50ZAfV
DdiHfjPaIs6i5EfzxwMR+u9WkBQJvgOAdkcoDU0KDHHvtJahYIfSIQ72tyF22jDZvJ3YwLuoyanE
FdBYZinB9ux3ynXqHtKMnZAir8cZkjpJR2vguhL1WlTwZLMl7KSCpxVDx71+6PFBR5DYdh23xefB
SdoX2VXR44GLJ3AtK8nnz/Y5uIhyhYXxTN2IMPNiuHD2xPGpgJZJX2D5EQzGH/MRynV45D2GHk6v
hxR/LJIjFq4eqdus2E8LzscS16/cQNV2p4Q9v+xZB3rdBpAPCwvPAH0WvoUb73lOQnEsW9buDxTf
DCYLn8FRV10BnOnvCAyJ61gslyjJWtkvp6uHBNbogpAYbbi2LDKmaQRQ20TAhhb1vVTsFVymKe9z
ef+WLxiktbC6rP5HDBhJIat8SRjVdB5G7XjbUCQSwvJdpIkNhGa93nvQkt7T+y7G0/2W3bpVFkXy
rlUDnZux4T63MWFT03Q2/02xjdA6H1e9AH/GWzZRzxyu22JsqA+BatOV6BGSHrypkoCVCPWtdBA5
XDU6BbkxQQaDqvIEzPf8w1+mwpovilPl2l9qFFUuaE6SN5mQVwKWKrygQZXjxCKKxgeTf58Ygla1
mVAwtKgWnzCG2nDCqaRGsJEONINkFJBaFW4+ywxdWxfMZUsa8928nbTUOcPKljn/rBNVztjw2GxJ
OK36+FhNsGgsP6H6qUaoQeW55DKxWrGnIrYHWsO8o8SIA+eKTgg2CuWSjlbT7m4F1QZgefOrUsEi
RIZ9aJiY65lp2QJmsIcx6QFbinNazRkpRceSSXgYXcOinXM37/RlyrdPncH4/h4arcX9fhg84NhB
9Mx6yoBDQWgzNNsqRPMSCyofLhfLLnH4M7/UOqm6KuHT8DFcXUOJdCs69Y9cu0Gi4bVhvfWZu8M2
K/FYjVc5OH2Av6eFb+1GK3Lk1kTOZzRtZS8LOer3p6h2vv6ua0kD3zLntNn8OeEb1TFASt3Rn50R
vpNW6BitC+N9/PWw7xEB5QNXUUwQtW8+pJl/u01KaT0S/CBTlDwSkIBuxWrzCO/BSjwUSfNHLqBt
fKHCUBErSu0BLfDdVAkPBQsiPXX02fW/10LKRV95UL0/rc1/poRwD1LJvB/HkwfdFP1+ZY8gWxIu
SBUPEQ1DfCQ6wpsTSO5U8sBJmxpXK6TcpxMr+Lf17T+cjHxLZhS9nqVEPZFiD+nUpIcKU5ZEjbgK
J98NVd1zkBnHPBH4rZtEaga1fCVqBldtw7xR4x4fcli25XbyoL0TPnfycXNyDD4wJB98tZDb/wXK
wSSiC/3e+IZ3+3kYXPIjRy+rBbaRzDTX9lTmPCZhzB4M3hs8Fy9iDBupK6cvTNTNO3Bnm1St3Yqh
jMhro2QI+JNpPzj5WkJ6GQDEA0UWPkqQLIAeld+ohx5Ca8/so/F/VZmryQmdKDu4cJ/IrrheT9MF
Y/mqku/fwi4HaVJcMEjHBBP710CeVjpC3bEpSddqBtAnBdVkGNoKvrH/S6BMRIssSV/B8L84QwN7
tK96T+kyq5OKiTfzhX4W9nOiHUwBxDh2DipELvPcWhk/B2hHgKOJ+od8IeJmqaUH/raGiSpl6C7s
v5UtQhGO6G7B9EZEE43O/PlgSpbxATCxFLjeUthIdss+atJIYK0pOu+4Ul1TFPKA/6B+c0O5dM9y
92bAqm+o4Bm0KPIEWCAzAS1jkCkR3XJQ0jJtaolKxWX3sr3qaMo41K6RRgVtx3s7BJYdvJDiGhP7
SmHbmzywnJy+IjIjftenIf3hXHMwBspMb9grrKCSdt4vhjBbEttshctg4jk9VbgJdyV3zTN7QIFC
9wnCdc3X+DDzgLUwli4rNYev/9PLn1AQdfamstzOySyqIdG93jx8XhnwnIxX6CUuQmm8Kec0KOCw
zelfyRrcMtkZApXXxB6rCv0AxJAT7wbVPHRkmN/N1Ci3dXt34VS786uyjZmnESK3JKD1u1VqyLhF
/K2IwEHy3/5EewpPZ8Y2b9syzG9EB0rmPyGhjv8Qp8AwkaHN/qMEd6u8Xn47kl4MBQINx1BO96aI
MH8kHMH4dUUybGfXPVonv5Qfppk44zW3rHWZLAuHMMG5OccWBBhC+f+gLOUwctDgkXc/nEHBlss3
lxn3N+yGam6l/FeauqE2CyGsPvywvsMpxsCQecH2wpmtTcw7VDsO7XKmuzvTGlkh79n2ooorKTmB
oRxG3Kl3L1rShrZsSQgQyEBQWqccWUXmck1Qg82ehjZl4hG5rv74E/kXDn/8UZ6EtczQioS45Dz6
lYSstwOgmHhSmzSnBk1816g16CANyjo3tMuQyt/fgN8rvfTbwk2Nq2CMbI9YP30o5cxR6bBs5s/G
MOYe2ISo8TzYsiDq5z8Z1IwpfVFyaGHcFiPWoYG/42rN3NITER0TeSaCqfu65I3z+4jhPppePQQC
jOK2KgR97jS72ClK2CfYRqqW5xu72TYh3LBKv0xFd0sIWUYtqBWUYrF0xLB0nOEdrPzjn3pRi8ql
3HYK/jzliWqLRrjG3gmVP2qZkT63vVcxIJanOoVVn/pft8SI2u5QFpYw5+cjIt5IWK2lxOXBle2u
ktKQ9EW4X3/WTKTW2QPVa8sH+9K+dzm666iDMlXYd/rCx/jN+0IPBdUcXSqNqm5CaJKJCXjV8pVk
YMSu4HMR7oNA+lpCzAPvBDY2eQdqg2hG08QmRIwgJiKPCWKVqFSDMfB+ExvI7AIyFda6qzxoV64j
EbXJ5PIQnVfMYeJahbtcWRIEEtUSeLaKPaRGll9h0waeRmNV06ByPjlT93Zwjc9NG5zaQ4MQflVK
aiug65RD+BjNzMgtqb/gAaGJjMkV5B/5xIPa6y9YN6sVVQh5jvvHI1jkAZ0w5Uw3OFjMNJ9Jfzz6
ocOzhWUEMaj+VM+FduV0hn83F/F1qObgHSXPwvSmxLPprxnqKqmM0scqguTVmfV7oXXp5uWgEflu
SRd4w4CMzWyAKACNBKetPGW8S4tVXHs0NpTDEXGEhBk1YteuFXcMR4R2j0fg/uZNJQ5N1XTUwnZl
sqwKDc2mhIwbKEgSCKQvjVnoxZVAPHkA+R9uu+3EZStu2/sxj4QZbWf3oCJUSugGNp5JQjtZqvnv
tUpLBAR8aczS2T8GXFMVFl+ewxCHXglxiRoHzlM+QPi6xlwsEd9xr1FiSEiLnr9/xFNpUg29v2wg
13yAxnKGHDaEQtf6+8XS3yo7JCIXvPfh9f3FjS6aNKjn8IvACyQrfm62TDcc3VI58ZheWdmiwU0U
gInNqmnpfhA2g49a8g2mbQPD0dmCKRi4/eHstB3pk3tYCBrXolMn14KJUu9aEjDWRFvhbYZM5Z/m
6q53BMdVuhCUyljnsz0ir5Wv/fiKYfvYMtBMmHi7awmVg+U9qb6NkRZdriAG4wagBPtOgSb6eUkd
YHC2clRaPYMypBVN5fBdQKuF5aUbDYe7TabiImRBHNeNQrQAE01DwtzXGtz7r8MbRtnsheS3jf+x
ZJzrGybtULWahSobldBsas60Z6ysgCekwbB6Bmfu8GU6su2dtRleSvTt81dvr9w3nkzgqQT54mXC
Biz/GV15PPYrcaQKsVoNx6pLvzmMEd0vH77HcPrSECfWC/e/sjzRx3FO88fvACYW3UOjOQZZPmZz
GsV963cKkkxZA/wLsnZ3YzaBWWMKzMt2mQ+2vIBu7cBdqc7jh1ct6SJtwkjptYIik/g+B+Lq1etN
fIcc3CDDdEGRT+Yk8lcq0RkEZ3/k66RPPFcL8hRV8Vp+RY6k3fGw3OSfw4Y5fekwq/3pKmynPtoo
cTQfMBu02Pr9On4PczB62hmRbriaTXUX3HihBA/HaHQdn2+kmyJHzRPGlVrp7mDLb4ILovhenqWT
FhDKmWZ0ndtKbjuzMyDSykRqMS2sTmdEMWILPviDIEQqElS2lhf/J5DBzD24+IPX39xCSFvnGy3W
3BbOPKwk0h+hTpnSNrO8LwV1gJI6Xl/eSIYaRUImiLxTfp67yjHyuWfQZjhu3k5X7IvtQ5GZ7n13
neqUpyaPs/ZqCFwu2vqfQWD+2e3UZ785WxARJUM/L74E5yTFYIjZvdbS90wXOIqqyX9ZkO7UD5tF
JSSdr9/QIhkuRQ4V5sKaXJBVk1M+1QHswEXVrSpTk3wTtCbYTTD/x1aK7eYvL2oFsmYRxGZ21ppJ
JFuBJMcagpey9QUgfwxU+WoLBCHlKIl8oKpWl30B3IWG+mr9tDoRaoW3+Dg3vAy0sKwuUuSEuWsw
TimK1fn1OjwIlFizq6CFwK2EDy6xL1HZn8cQgCC3PUsfpNC7w0W74XMVIMZt0x0pzi5xe/zMN4X+
FSMFvE2n7v3yrJgemXLPz6zLDaAcGCMsd/T/0/mx5ISZNz1oOTNOVGYQQimpU7K9r/VCieZMFzCQ
UdsEpjwYQKrNUYXD1Fa46T05NYGaiuSZdJ3oWIg1i0X+Qbf+G14fDVE5lXCLTVecvzKbB/D8qnKC
bJ0d2JxFNCIndTbhi1lxMR0/o2vo1PNpxsWjuzzntXbyXpVJ29bkXynrlycXQ2yWqUZK8+TZHzKs
etrbxiE2utAY/yzsg7bL6MvU1K3bRonj1sbvg/fp2+E82UkoKoCKtLPEHb+JOhITrAzky/yW4eU7
blqAKBMPBYMZqhP8t3Nw6GSImpTbf9LlSYSeYZsEDbN/RuI3TnCs9VtX8Hy6WD52c1Hi8z1g/vjJ
GMJlDyIhTA5/FxqUEFcJquObN9BXnPm0Ndyt0aH7hcYahoNmNg1ClI7Cop5Idnq6ppTN/jEc8xrW
sv3hfu7Tt+FLeJ3QP2FnW29Zj7AARanUKnfdkHXRNBXVlX7pzj6ReyjGVgOo6dnnzT2fwwxG9fva
FdJIrluhwkUMKw4Q5peaw7Jm++Ox8TwKI8bp8xeoiw0ij0X3SvPo64/g4NVLrMOSWdCmNkEGQ5IT
X5JLW4e7P+lz+/UxHCpDNAwOYq4MjpbA+ETTTN60CGosBmhqsAv4ORkgsV28a2/mgyiN3K/TAfXe
EC35XCWxxo7XxCWmO/4bNrdGjB3Jz04t2dRvc5ZauVHZ82pjIAzO3UWjZNzPrNeBN13OxLq9bXgd
k/ZOapR0MhvRqi/NXVb0T2+QzHsNqza/e75GD9Ijg5tYiADJlUDe6mfWuTeqJhWnkgUWY51Lxm8d
iScixHuVMi0wluEpt0P49PhhqTjovnoSHGZZu0ZMqPE8tFYioDPNniQwLKFEQQUsxdojzuAGoZi6
XdMjZ8Zd/JIMnJvLLfwvgNak1gsTMiMhdpSyl9jYcqX+/EqhXcdxNH2C87nruOU8JD4+NTsz5DUY
ubtg3A8Qls9tp1kK9tOIr8HBjX5ZLE6WZsA5I3M5UnRt2itc2hugIS6i1ZU8pHUWVtnoThE1RyVm
SGGDAnxBeObN2XuJvKjJeArN9Lke0AszqegqUM1sjxIfxhx/lKw0sifoyIt/EGYWwfpcEz2DfaJp
iMgDep2v0TO3zbE8naMVoXHs6zUMy94arjHYvILL0Vw7jnT661sMv467HXJaqxmOrhjYP/AHyz8X
TrGXycXiZNZ6Y6etThg2VpAva2jIS5RJHZVGBZTUlfv4RrFwtOKAOfLaPMxXlipyRNLYy8d7wT38
4WqfdCsX7J25JXSrZs6lwQOCbn2P+CwP5UClT6gCWg+d7el9Dy2my6Jjrf4qV4as+Czn571FiixJ
Q3kitriZd+encRWubRJHEwN+wCWKp1HgtKA6fKxYdQB/G5PsWM1YCEG0tit9/Q/bAWx417azhARV
hkaE4euPfCG1JsnFV/CR2A6itBC7bob34S4t36DOIK+ftc+PLsrDF6oylVzBHXe5tD7h/LGKvxew
dxUlchiLLi6bUYaxAOdsIcgiV6sDb1To/aRYM90xfSAXwaha6YPYuaCkjcdRhE32T+fBgxD6Upfx
YZmihOtxXQfwmE0Ws6KOVM0sZ0PawPqso3xyycIlkziorMVr1hKoOSWJ9iqUJVuwZe/z4FbNTZRx
06nLe64JZM6H42i10Jp+MxSB72y8QXIIQj+RE46xJXKtQ24ONlX1nqq2ShdExypQBP+w3kyyrl4J
BmRuA1deDF+mbANCwg+8UVTPdtgqATu4G5NwKXUq/BJPNayppKEnkg/6HP0JgVJGaiRti6wWbZoP
S1Jkbumjq6E7ayySE/uVoztGwJqDZmp5VKVZG7ehJwVOePwbM8fA/Q/ufvx5qycEA1WAulzPUgAL
Wqu5CafinZ+Qlo5V9VMp1cOx59alwmh5SGucY0fu1fGjsH2y1Nz4KRoFp/LWM3RkprcULm/LNCB7
RdFLi8PUZWkdA6eLdEMlYE3z7F4ZSy16PbdVFuzauE8tA16TqhwSWrIhnRAv9JdkeQLR4ks6/xIG
2nBLZhw/jlBUgUQMJUcfmNr0wiKf8vVX7FglASjF8yFr4EZb/rzd2GJCesTZVmtSSRaOkGNsQdRh
6PTdD2uToVSjRiaLaOTLAJ6tCwOaTLtJKcIZ0pNixsj6WyQWlelqW0Ow9eQhKUsNMHkCIR+WSp97
bf+5NjbeKxVTjgdHmmN6jtQiN1QUzE9/enDRK04ntfWQ4/kgwwOInZfxTkucvWmIrzeFmRDgsZV4
BR0ixNuQ+0eCRs/xCfrMLGuP/7JqmGAPlcx82fJYYfjL2edHiJReeHCKvwUhmgy5bW+K8uA+IrbE
31NsTwlO7OUknvTRX50jDMGBDYRAzg5Q820ZDp50aPzpBmsUPs/zsbFqc+M32Vp1aBveIgVLFvEi
nXwfrDico6JwBA2cmpne9D/1TGOhq/NgAqxT75rJVeZ5nCyDrRgAtr9HHNiHCzG4c5kb71piz8Vr
DMe8v6QhhwIH0hp/lhJb4znqBwmuwCWgF1ybjdl3yfTcXiFIqFCMZJJCspeLcpS8lVLYCaJj8eh1
KTh7zZSJinF3L2sN7DKmqAfQHQXmh/7/JvoKm0C0CsFdrWh5f91m8N95s0vGrXzS7qd3e08y8hC2
WCSNBn0Uu4fkp+m8lZn0NgCP0IsTJdHcMQVFuXd91ad3L6UNfI88gXfXeV+c+ZgX0syVd03g/Ge0
XTUdD1eVRMTEAEZ0VUEYUj6dB6XAZF7nvAWcDFOL2U0ruaxpAtogiKPQEjspLGuc1N+EafM+C/Gp
6Az+PqwebDoM2E5fzZielbQEvDIT8cDwobIz5dHZo6D2P8UTcIB3g68womy4l6djjXgTsvL21Gce
AS6+VBfUaT83svx5ITilhXqNCkjQctZssA3F/LxKkEhQWlCe8jK9/EvMAm3RC1vM0+13qIPxIKV3
w36S7ZMz01WoIeU87tv4TpgijO4hnG1rSApNaNlClggJ6M09pO7wBZYALMtW2Wo+weVyQ49pTkey
Evx6AZ3F2t6GVGDTVKR9CoawK2lZQF1Haiqa0H1ss/yz3S9FMdXrUgmfmSjYtUu/bHdN+mwFGrDo
XDKD6NMzxGFdH+Hdr9E8rxWP1dd4iR/q79Zs5I/Xxbh+5GYCYsd6rl4LA1RrZeJxSjGCpgQpNFo9
18Mk48rIL8QK3z6IOzZDYRiVYT4Ugcb5OWabulynAgzJFDlG65UHVF4hnGZpUxtL0+JsSwWkgHxd
jDQQpLipAW9W5aR1T1ZQE8dYYSM4UwuYZ6oyr4yiuVOSduFAY3aEkrpk8JMfr/alNhQOFCktyqUh
8UTwpKCUOBytL2UZl3G2HY1XPbBnkNliQ5f1VGDox2+LD5p3vqDfhy4iPqGQfuIkBWy+GtfYUDqn
LySJh0i3XpuxxWJ5OkcLwR58wU6QOR/E7UnXXq2BU5oGJLFgPaWuD4C4iJVG73NGah85a5s+zcGA
ng95frebMfIF9Uoxu+MgnFrFNUd4WgwqDP2bQL4Bw6El+Yr0T6rR2AY+Apunh9WOYsfwHgHD3G8C
aCBVkBHraFB4H9sQMpxsVJvdBj29FyJtbSmObdy/E9BZaIAMmSDLDwho0NmKh/7BU3+WMGSMDkrV
XhMtZrTBXWAkllYHuyyJZzzMySUBTXM7pmBOrghbUXV/F3kw/eTgtU9d/q3aYG9e1llmboQGet+a
O3iKLBUtkOnYZlCcMLfd3qGW/L/4wGk9s8FNLAkvZDDpZBBQtaQnpGtECOdJ6crOMiq7Rm/byFXH
5yHAZFQVmZZeq0ajIDMzfVgXyfmcOBpoex7fdSpsdAlGeZT2dH6/Ao1cPCnMimSc8Y1jgQei9tdR
l7eqBwyZhRtRhsaAXb+Fk05swk8Dw8RLOIhM9KupcfnvqPdOGlcXM4cx15temGLSS7O/sqba/cnJ
wxYM0jS2Rv1C0f68MVX5mV3JowPhi8nypqgDl6jxNOjB+AzVTWA3qkRS9omv11lc+3z9rwBRjJSj
kajWQeUIPrr4fl+ZCDULERdjHRIE9bdvN5m68mBg8tRKvDrijyProPd6Dn2T1KWBAIcaMvW2Xv44
iQ5py/bpyUHiXzT9fC2JJdCnhZsbXZJvIEJLdAMon25ZITJ7M4RP4v8d20qjF286k79AeGMk//LK
GA7SjglS32YLh8g0Yz2iE6gQWuDdjeb3a4jlv9kuzZ6e4eFm5ZPR1pOCZZI/IcGjy1XSQIrh5oSv
tA5e8JFdKHXlhzgJD6ib3SPGLAwSvbpf53knwtU0aIUUnApPWSN1X9dBEa0wPGkYF+jIY8FJKsbh
nBoAX9n9ELG/qrfFsGDr2lA/oEUkBOq+xuZtDbIBfJcPPkC8oUNA4j9XJrd53FC0faPYEOp3Lpg0
eKOLf5knbC8n31nVn8bgdLiwevKOUNHwBnC0x7uYm+4Q6b4jqcXZ/ky8ot8zyI6LKfga/9ABb6cB
Kfe1dSKc1NVb4mFsGDDOXh4nZ8Cygf6BH7yIs2EfIhFnuPdX0akbGx+8Ae1K8+LIurNmgHrD/IF6
57E4bIoJ8386RgudsBYjguuGWbNFqVdMiNCMcIUFJAcCBBNxXSIkZixZCDypZFjenEZvULnOON9Z
LHkiC1s02jomvcUpVVSmAmxoLclLndWyb59C8aYsjJGTmvdXotECO75hVrGnVRGa+POvGR5OJ+9C
PbRat8nJBRpFPbuY20MQlzV/kPeGF9OpcDAjjRHqDDQa6ETGa5w2Zhm2ARzeLSpPHmXo5mqNP9UH
FyVx+9r7QFyDr5WW4IEFGSgRkYyIFuYyPsDFRWeh7imOdNU6M+pVhbzdTx3UnyaJV4H5kvl/0Ya+
XE6jycgeXfeyiNLEHhUJm5UlIWw2kizwEBA/xvbXc+RxIEYRwonQBubkqBCXeuNfgFZ+lY8ijcR7
+CfccxC86BVkWgIejfIh+hP15yvf3OCTa0PZqXZK2bMCrLB1sg6Oj+1fFDH3au+8yQARHGmUqaML
V4S5RZog9v8PYErVkY5Sf7u1u8TZZMOugd8hdLG4b2uvtbU+21x5SFT3oLUvQr5HtikI5r0yy1c8
xkDaqSylUTYHgwJANzRkUQj/BZY2D5RTVzANJCt2h6FcY3kwrELI4+pyxaAol24/wOBVHYlj/RGI
TggE0Ei5OVbWCErmoWL3+JYqHahMQ6FifTqhVdA2E5vOlfoG0luyr++u2c8YiXQOZ8MeH+DnUR2u
Ej4XXBuYE855gP5o3ljySqYqSEfQpOKZQej9fF+v8JS1geEqoZJWPjNk+D5Yr2ySEZFItEytSugj
QOXOtnI0AFZ/Nsv8SyfOETedP0Ysu2RGkJlm6kQCLt5G4AOb6aepI04F9QTNLe+yNUJyECdHyCrz
bGITZ7sGKXgmXGQGAkaJLPwkH2I41FRkMB4a6kKaaKB0qmC8VGtdDRL8yXyIFEFB28NprtES3rDa
qISQYALCvEKW9HbYK5kqknvYBHLjBEFEMImcLundp/zNaMjHToA27wstWBDQIGRRrL9K1+ELl7sk
mmGu1DaF5JYqXNcGTzLJ8TN4OOWM2trj5txi/+1iTouPAvsp1Umth47+/zLG0MajhK+7+Hta9xZ1
sfabGEAX+4RlsQhrIaq9FsvdgOyKrW9uBHwGsKUMi9AIlCe9Az/qqw5Ia9pCetcXuFOKYj5x4SV7
K1e74+hty+83cDrNI+W2cxztm5TwG9+koUr040yH5DOjsZ38EGr3a69W5oH2k8yqY3kWWWsTJiqs
e3cHff4J8uWrlXmu9WdlxGUiz3VcziT2/U0zH9vNwwsWd9RmIJ+N2mxU5rDVWBiyPYqGws2WGoR+
FTtwaqdHNe4T3Bpr4BPvY3FXbwQrhr+P4nDVd9OMK5vBgXUIp308e+g4JJYhAshm1V5nqQ2db1qj
mPPUGCvw0HVk79tFJfdUONiuhWSbFdPMYGUVLVhjv/lBdQjXH8r8HFGNEiKdei20K9z3inArsnEQ
bIwgDNTRHDEey9Rftk0NO/43+Eyq5hbeJsXQooIBWYgh1DGCCnaN94BE6R58srTNwfG9IHwfUNX5
oAE4ASlICQTkEX0Qj29ZhhfHlPGl2VTMYG2umuoua7Z3idEW09CEdS/BMUtyqkjGIM3hb8Pia/es
80WdDIg3Z4e4zrMJKxqznep30EdWtpfvCn89d1jBxOewjvV1bqYu5aAx3nxbhq9FA8v46Q3iPoVf
HFvWwy5mXVbaVrkZoc4RRK42+y1TyhDdbh0bjFo2rz0MTJUz0X7D13ujv7vZbpxCpWMMM5qtzFtw
twVlqPE55LGPsKNIFe33oRORlXMjbCxRTgTIlD0z3TyQbKtMBN4daa1mEBLUwlOuEubfgOD15pGM
iB3xJ6TxJVgyT0RDYi1FJLBMwpqmMByJFpfH94LxBqhrVHIhFExWUrhfyoWeIT2hVBmwtjB1Iu/Z
xhaX5jYvWc5VOrN6gaq3eTsb0gwgCjrLEFXFvqVQaeNhPGblQW3xENgqq86QDwf3xbupIeys6p+h
o1ZJfzry0zQiLTq2mpDMAcHFMFSgtuH0+WtMByj/L1+fq2hQU51OdRqRLD2hXWj4mYC183QByzID
YPRZcWHDLjbrN/fSiGb9FX0eiXiMNejTSBi4lQ1UvQjJlIqJH4z4btd3WqQ0/oA1kMXFjVLZouiH
ppm5c4SDzJzZPqfRma3/9ighWBGDmfF6VU4VKH5iEoOhpUKDwqW1Bytn57zuqQnH5CVvA0X+LWsu
inyOUV78Fan/4hzbRgvglLg4X6lEeTpSZFWDxU0IZH6wfcJ1JRVc29vJeJKSh/KUP6x3+GdEkqiQ
vecAM5iOfLYBEMSlv4tY4a/3TZuwwyBt43A6BYRINg/DNS4UQiXOsrTtwP8JLL835Z2Ho+1OpLjh
HmKJUwvkv2wlPb353SHvjFeaUHWRL9EuHifeRTNHO6Y3kNvPPsprzXJcSMeUZYMP6HCYMJOz9xvQ
OQNq7Iv88Ic8T4aQ5IBWMjcT/SlfNezj3r/XRgow9HauROSNwHyqNWWlUvRMIbvXx+jPI8h0iLhS
FlQxVMmufi64ImImzA5GT/CHfgWDgLF+bZyKKGu2eo9SH2QR56Bq7bn64RZ9WMebff4E88t5M5cC
+TXDg7Hx9jh+tb9CauvLLksXD++7heGPGMVE6SHd4uFl2jg/jak3qCjpNyHvJ0xT48ezUDtTuE98
dK6htroo0HqG/F0mGWoTsPo3aar6RXRrWJlJ70MxF/8q0KgyK5FEQjzaohc5pcDSoRTWxrQPDHt6
1UU+rAtSWOed2VvR/AJLNP+YD4Yj3Y9O6q6RI0o6jaPwBIJfqeiqc/eyQi+JdUr9EK1kdCAqrLJT
tB8d2WoLd3pJRbYDdnjof91gKRvRmSFhDCHmn81KIrao0dIm2IxtjkYqFBoGPuilfe6yRb4n3Vbi
KRMWdFvYQ61K1EHjRsLdUa+jloySYk4P98Z53y1SktXuLE86d5Z+YVBiV5yHoDu/tLO6EdHY2ptu
nMST8Xec9sUz4Sj61lPv6a2OGG89EL3vqk84PXDAhKTZioO/4+aWjS7IvsJx0cHL8XxPonW6KVun
vMu3v0PrpOkO05sW5mdfkbykQmsq1sHQIXDOCwanWaEUurIYkW4PBr12TWq1Os4nRYmHsYburFeQ
oUWKCvBVd9Fy3UKcpA++mf9tIOZBLPm+3eM17XpctifkyD+b1zLIzC8fcI3fMLGykUuiHkHKr6Gx
M1UQfWKhAx/eODVNRd7B0MYiZ/mMHDYD3hNo67iOts1QPOmpSc3xwxImsjujaFyOhcybM1Joguom
pqY/b9iwWbgdcSoVwib0nYVe40hGuo41Y3+JOhQNdaBsddAgGIHuimbIPGFFb7m68rzsz1XpB6RS
UYKqStzd+BuAbVQyCKB4HqMCUVWENRMTUcFmlfIEbX/Zyq+GG+e+2EeyWKsCVvcEonmcOlmKSLys
IXc2NEJymwWSvuUS/QEZ7qxybkHcMLYcVkDWlABi7DTxKPtHPtwCFL8C9gcm9OEGG3ORijsxyhnz
plGJ62vpxcGykug6qmDfBcmstgEhA5MrD0TS7D6BDI725YZa5TItYKCOC6RVXTz+y3xl0ZMeWVyA
w4VESHh6QY6R/YkMQu92xzRo0WLRSHwqjZ98LN3zkFsmU1sWU65aRmTefWNdl5YxSJDvDcN9i2OW
Yx9vFz/EPubexw7+rEyaLZF2qYfrVak7c4LsAkzoCPO0loisbnvYKQBKLMCRhcc+JXbigM4UsABd
+qU5oAL11taKyqsit60vX6s73x49He6pZjmHSGdmDDet7Jj5Ukr/U+xftzbzQcwO93FRqvMFmvou
xNET+EMbyBSaGwIMhLoRt4U4/JG8J1zY0upR0jCe6TdclA/4X5vtElvUJcxo/B82NUbXFlYeQNep
8QWc1FgT0+tdQhVl30O6gKKPkydpbb4XTEAINsYbbde6zShkTAdDZ/YJx5FCXOBm4oSB0GELhF7/
vncGVIUx/YdVwdDBYU1M+iDcgQUOdrFPkiQ5CqODF/lXRLnjh6s38UL1pAUodDAeOkldsG3ZU1aZ
Am/hr9GmKTjnvRHFExrLKco4qJs1HN0iaQCxeKeLqSHDrN5tepcWProZul3w71aTG9lxg0v2lcxS
RzmZ+WhXO+f2CfrznWl7bC2loOtv+tS8MjsR379/P4bj6fnvW/VIGIC4I4/qn0fjw4fYmSbWROqI
kYtfYBKkPwQ7LoNS+dTcBxH7UlLe9mQr+DQONgQrG7daAc+bHbVPPzNOnXBUvxgE/9F/4WkEsz+t
ux0hMXDF/HHLmnqzXjjWn9ifgo520DCqKPjdeXVc1m25JO1A1MbXl5DSDih18T4anRHotPKTleqZ
WjL7GP92VWA6ZHrIe/n2BwdsB982HKb2nRj85cKbgzKs0Qm4hcx5U014+Kc/TsV+Z1E7X9XXYO8r
bFIGrlrL3D4eTjFHNY5H81WcUPUZkhNZa6OwTJlzVQrrMbPBkLbEjaXthqm1d/Y5ywJJzbJBKlci
BtoFQlAn/j73hFilNWkIMLg6jgxZzKAQVvi3/lGABtiK9Z+pXYT/w6uwykKHD78WS5EFCW7qqGCK
iJFeJ6wuehACe+UxbTmS2JtPRQTx83yuQzGyM2n4LeGw5vZXJCQPTCqvYq4YD8qCQZCtLqzmFhdc
4+nWomCb5VXooK8/d+bl/J1dskuXPD95+bvp6LRnjDIUkII0TK/lzWwsOyVwkY+rEo7n1DZBXEul
YD3Pdi8+CNkM8arF7JfERx5sBzmYOZOXOUiR1m8rmn1yp0Wx9My2IrfYqu2x569XYP6YKG3bx4rm
NU6O0ARBamqGLx7eiqhDfMYeXPu0DjJyDxiscdIruGDZci6lbBmwSxVStzVXmOENIZ4CXf2n/h1a
VMV7w1/k9TxmwK+xrsoNunQZoF/uX0BkNdAqNJBPR5iBbD4uDYMylsfSS0P9LRkrozCcVhjlFA93
1wMieOcthgN37MH6/8Vc+/PDpK8Shyl46pLdjbuyot2ZPUJbbfDgSKrrQCn1ojMP2cF4S/JTEcD6
ugZR66ek6qNBmF3N1CWhdw7IpBRujWJPitfaweI+wofTRogv/p/GL/mSVWFEyiLdgXI7j3GMMyDV
TlXGk9o1/UYJAlpUy886dVO09gspTTK26InT8gCaR5886XfvbdyDLFsN/UT+CnUnYWNzitWwQnpT
HiPPYnoGLo7n4ywVzV2reiA2cAYGAwdbZSFsmlK1HtvpmXRmHO+ZYPkSKtsMSLJhNZeSMRgxIFBq
dfaUZk0n8XOaKlgYbuZw+IWbb1T2CzbbQKIcs0+gLcvci59JKJD+k3d5LWp8kDRDR+nSASMW1s4o
xsdVQR+JNKur02C/GyEa7ubuLzZJxxID0fAV84Q5ckBi+wfsA4HLKt53zB8M59KY+ahx4SRXImaj
hg40UGW22FaW1zOjKdkUxigiRIX0WpAhsL/ctAmS+BzS2gUTdMbcdhTEOmXlhEk8igwsCaJ4tdyp
0XV7baK3QveqTySQzAvkj99ynFXaLyJSeYw3aNL4OEuJsNAPRrfICoRLdLBgKVS8WMqiD1uPasmD
yILSsX3RYAVn81OqUvsg0/SnFYWUk1xAJZ8PFYIsR5dTLW9LQwy2DXBGRLYJoVKIc7ZRGbIodbDn
tnb6PowGHE5rJb5SqdR65nHGrzSrQGvHPMP9DWPz03v5NyP9Orlt4Y5NBWmyTl1/AbjpG8II0xYm
70tYKWxkiTJ2fXmbIAKqvWoJ2LTV/LFnQ4il7PmTZUKsl3kx1SRn/GBmwuRwDGzu8o+2Sm9Z1GgC
dB9RudTJOcqRNRuUZZ/AOL2iIuhB/TBRUAfmyhEw4ycqFFQT4Ki2acQNlZFfciC6FWmLWSxCs5hV
sD99Jf/9Mas5fICTtCA8XzpUrCf845AwCEnSH/iHyzTcnpH1Co6xiKOAGmiUfAjCAEI6p8KwJFL5
wbK+u62Swh/jo7JIkhDdAU/pvFnTaixKihQnWZl9Mm3IQtzkEUGJzgTysUlKVBG4i+fiwLtHx35G
5lrYi3x27hXjJCoPfbub4hjXXFIiyruEocoTvrWiBAMAqnIn7i42S9wB2br1oEpjEhUVrYzORHQJ
+GDJL2dmWIinmEfGhmmGRUiFEap4z2NWbExWDGrlWAx42c1gVitCLax0pOpNALM0Y3szzS3bCZAl
g+7dgAyFJCdhMviFyERBqxjm4AYT68Hg6C7Ox0TvpgbLPeGEAYbzEC0yhM/sBFjvjRPNcuswo7V+
zCOeZHpcqCZf0pnN7QAlX6J5v5te45QlkaLOo4pDHMsLH1R8Qi7aam0acoJibNNbLPRmRQE9FUNs
X9ofEhHCt1ikhQpstJJwnqIdzUAtFWSE7AVfjjd611Y5vw+EepZIPR6dxtWs2rDrLksU1M0gKCm4
BOvX0Tn0Fcgjsre6VpP2UTVCirt+lnM4jyX2Amr/nIeqVtxSRqlJV79G5owmGJcURIO14WxfEYFJ
AlYT02d+2XMB9HiB/palD34ldEhlA9o9rFqhsn6FwhqhjsZcPg93Guv9VtOWrrqrQSo3S/HP7SjK
WoZfGL5WiRelkRvDcU6EBdlSRr4qJYN6zxdxWVXO8qIehzgnPuDU2NqaCgJOQbDHjHuyRdRUGvf8
KO4PFnARYD7dheHOpoJKkROkRIHWECP/dAf7BcDUmEnMLD5SwMWwkUgAXY3EXFLYSwvyakFE7j3p
pd0fZ1T4Lij5hQotErQNk0WKKf1HnVHUFMTi01eGAOL6+KE7bFgM1auAH8lE7le1Svh7oeqQ62t+
+/1rBuaX+o9WPonqqBi5ydB+bOZhvRUVlQh9EUfPe9LGyK+3sGn7UT73BCSD+OtqEkPDRfDmHXMM
qSpFn81Nagghp0QFKFkVghKoHxOZ6/NZsKZYZ5mZ6iT51hMlsyEl77cQRFlx+xJykBBhhZi19MX7
Z6xb1zXu0P3PLu3q/ezOb4OQ5YGB9z7kyxmySrq6oW3DptfT8V9lwl24akIYOLxkHPJ3fy2GFgsD
au/xMkSFFOM3xPfnLd9LN3ZH5mOPT+lV6FgCFpiMJ5SZ0P+VvS2opcLFuwkCVM7AaeD5dv1XE7L7
0RML2gPm97hOg0kGU12pSwM8Z7gzpnmQtGa1kOLtEnnTgTs+vTzOaQjfZUXXzmVtEQBGjsf+ocMT
4w+Fb3ZZMbxTpgUMlpELjFD8i/ekpK8Q4ULwqrWmFWAP4PAfPfuxx15YWH2rC4rY16HithSbE23k
oFh5ZKP+O2aFDjg02nZdXNQeA9Y8PGqIREpyl7N1J2QuCqsNPyIGWFnGxRGWSB8BwgOJhaQWodbG
dasYKtunDsWy6yG45c75cBMYNA3g+eq96RKv+uMRClHiPB9yUQX2apW+d7eXHIVgOBEBONBuZpIR
5lTRoQoW/SUtNFAyMzU4Ghin1+z8kn8KUnSY+gtJwm19ZW5NMzxnlhPhXIVPHkD4u89B4SO43Ktc
/rTxqmd9UWRpb9o39qgwdsHyVKCWqjP5L941Rvc8HLViQHMUcCFLrSX5xCtFwFHxrG7fl9u8NOSA
eukQkm2E8eP0SNqZA/6pADUEK0mTvRtB3beG9Wvq2jvYvb1ASyVs4B6l0D6I4lEDZM5Zy4n/ME33
Kt9lM4xhUv186LN72TQRjIXOgKStOuR4lacMmpWod7yRH4SU6ni9ARfxWZ6c8QthNC0hGfjBJaR7
OHCyM8c5siboPpuuE7UndF7o1zpHALhH4BvM9DUGBhxddOdQ7m94qJsLvLnAS4muD2IRit0IWLkM
3IyqP47EUZF3jQmM746QI1FTqE7ZDZrXNhY8W014eMqroVv9AF1RI1UmKLGOo+690O00MlRkjHGU
wPzF9QsGoD3ZL5YDSjtNWk0u8oSSai0tgBcL/hJ+Bf+nE164vt2wXQ9ozRLFsHruJ6scxvQPHhlT
25IZqbHSu2A/Kw6Oe8Hy7Oujnt3If9ngQS4/a8G63WCw5f5AqC0GqYn517x2NnpBc0OMNdql6eye
6cJNgJXbPiEjz2dV02fI3OBuo2SYVT4VKFhVwAu/3jyOOxXtoTGfVUaJuPWlBrx/zxy7G6w7/3n3
/RbOYkGh9M7eSobpbsUg6x5P3jAb8kjkGh7dgHP/9uwCdzdLJ9yH1OcaLzjeVb640PUmHfnTuMi8
lPj+9s/0qB1jGhICVv28iHLE/1sdYv7Bpnph8RrtLdPrdnjKahtG8v7Sp9d58fDYkMgZd4XcymlE
fCPWNzNChA1ibNebNXs2UNdzIAywFTjHJh1dxJu6V0Dn1bmUQMoQVnDp74SU6esVqN1qTfaxgH9C
UsuYnWyT7Rk8TBqcLBcs29AYrtVDOZatNPKklkVpG/KTUN0aNzAtn+it93yuEnxq4Wef6q93MlLC
dTTdwJuHjSdMyUyJGGZ+5eckbzjDxI59QctlBwN0rDG0luHd0g4qpQYYIICqnjEQsN+HlhoViFyO
W42r+JHZ5QDP/zeyG2rARR9Q4d96UAlbRduP+XWVoZG/z3/HAiVPV+jZ9dEc0C3kzYIknL1S5kob
QOCllu3IkWVB5ORdbpCTkWbbPEzXFtED06RNvMS1qQ+TE83/+H9oRkW/TMzd024LNdmPFJuIVrUj
DyZTjJYn3bWchuPxlhePjiu/Y2UOwVD+5ui2miGGXAMhqOoPW8Tsji2zIMH3ozL+n7tTGWIFionf
fsIe39Sity09+/8qu0LduQVAdkP5LwTqM/RbM5tIKfjLr8AVrHfdQpveVen4xXequ7rI/dmQrX/D
fYmud0yJaCrDqinqMvyOko4edUZ72efSlDMXeU0f2Wxx8WQn6RisllS/pY1SI7CpTlOdrm1u8v1C
m0dhEykkaymvZiEpaST+cvhKlvm5GjULh6gKyxTZ3CWgiYXmjGQRJhANTwk+HshINcJ+t0cRcBz4
R9AloK3VCAoAuJF6wjaFzhH5R+uskfCXpQgKX54+3nALXPmjXBtkvDekKtaJRYH4KGFft+kUPEOp
+0eaAtgUlozxmYE5y67DMDDnn/ZFzSuQaQZIEWPEGZSwMU/qWs5fNhfZqEGm6tGx6qqhum82ebOE
UWmSHbY/kl/pAsKPlcP81qD5VDZgbdNUWyZRxhIao7lmb/vWpp23lDZAWs8MdJfpaTa4qIg6fLiJ
3o4VSs/oqBCp2XeWgN0DZ92dDQvJvA4ccsv7bgrScMO3NLDjrZ69NKQuHX1V1Zq2nl+EnArSVbeM
LeBi3rgZFhbgIzjmKgTZU2jPbmZhmsyNnNJt9iKkH/bKBn93M/QYF33sYhatdqgXLbmBohZ6pj1G
DueMEw7d9JrrHVn0VWyYabM6tGMyJmQWpZWoiPUZFFU6pBE348KIFXWe2BmzVP01sbtRqJa/hvIW
SwjCkYjOSzmqt5CQLlnPl6ZmRiOE9Ds5cMoePTWZu5lJ5yv25mE42SCTxwER+aqyRH8191K9CBr+
Ht/5evh0G9YjQltybzCgSvREfRqdTBuhxU5b7HAsELPtMbXPWmMjYjBj8LZGChTcrqCmc2ivgEUK
PQsDaEBuIijpThTv1N8dNi2HYdVraDDg5P5QH0IHJneXkbJTgsa+gBWNINwVr6iX61wu6g2I/5+g
A5xZxEGmzpLbxl6BWnT8Dh+WFtAFTJT4wgbkR4lwAsEOR6Q9cKu1wznk2CO7ELJtfmpLAg4Pxo+/
zH+pMDcObtzH86fI9grr7CuOtGCWASeTttB85OscC2+P5Gj2AinmHuO4iF1GRK0nSr0/1bBFVrf3
ptDNGVKgI3X53DRPN9Hcpa48pW8e3pyGNUqizOD9YA8io+1Rmr+1zxkOPtmfIMIqzod9b70x6CNW
ENzRPMoYa/PtdVsGC5/mbHKPWdgno70pKlFzYGe3NLJbHuO4fKqWZCZ+XQk7+IsASrvlSJtsViTL
BUYqJHVPGVwbQ5q2eA9iOc+XmrEYqiPKp9ZxpmlWaw7HiWkPIcRJzKp14ElkdY/RokHvzro8R2c1
beutFvGk6yIvt7wnNnz8HFOVETrVXqzwMp/a3qvq8rlTINRQuQMfAcKcE4+SUPzX3SytHPwDZ55j
9lZd/96hHT3E++057H4MNepsikTn8hNIrOK+gByNBo6J2e1xL+/hI/DqLI/w3FgEOkCl0RF9x+uF
uCAqEVe+1V1cWJMevBeU0D1xt+aOYvEeQh01kF6ONbvAgxkbNpm+O8XWC5A1hmFBT3EpdETn+oJr
i8XBtYaYRqPODCfLmFs2d85yD/W6gxplH/BkZrC0SCDgwOhKsSqsxfKG9DFQHgq//MyGLF92MPBc
O8m3w0yQ5zZwDnVZW9fbZ3rhLG79izbON9wzLXX6gqcHIIXCYmbUPn+urBqB8TQR5GunNhestEvP
3XbfJqzwOVUy+cRoi+XJvrHh4MHu0o9xHQnPiphXUonc72xM90MaxaL+mH7b5o08fQxCKb35hTyW
dwJHQOS07l6+cvSXL7khodF4Cdj3pFWQQalHLwMCz8YTp2ddGxggf7OTt7X0Opuw/gH3UkLFjdUw
Wek4BKaRCuyzpref/b7KCWXTtpIdkesCKxw2QwMafuC6IT36F6VGQoSRqevqEfJvMUgczft2+GAu
TvlQDROZw5Vxr+L2DiWk+5c9/Ud4yziU+1brw/i0n7I3lgWY8RMQRRQ+eW4WQFwnE5eeDiVWeFZj
pUKthDG2AJetSyPyvQZpz8HJwThqQw5epKQ8MIHvOc/Ih6XFFOxEan9XuFReXvP6H11LYftMrRez
1y1F1XCHNPJFQ4opQaEXB3OFAp+F9ijVw/yWO76h34J5eqELwNyHOdVIPUEKrk1PWeVAv++EqROV
LaweZ7ioCy0Gy2JbBtmWPnEl0/NmVeMjM8c2HXpeSS0mnYujM3D0mUifirCaPj95YPJfgdHs+n1z
ORqkhd8y4xELhdHp8emrwkZXi6UqkPdqioIs7IUu5i87bKeajHv1L6w6vdfphuC9c/GyTDqB6ZtA
rQ77inavGKFW/K40l2WZR4N2yhPi/eSkmN17r4EBsVD9WuvXwlLjcBHYDsWvPhMUDwhAaabla5Oz
o0tEdwecvriZB7hSSet9FTzBourRPWbNek8oflD82xSQVAQc0jMrpAez18DysLy8LrpxzjfCUpgP
gdWRtTN+F4IIy2BBjeFJO3WxrEKSqtfcruqGXmqwcdJq/CFSIy21F+Kkq0Zcr3xvLzyXoNe1sG8k
M3qRQ4AvPwfdLK7ppfNNkLSBsqO+VtEGGgqXAzhScFs1EHb0IZ8BKtdzyR8hfDiXMcLiDSNtaBp/
j8FIcnl34pzeVgGXM4IFlc0HlgHtIOWJ2yKTNbD6h9S4pPxJf2wnufvE3P/XpEgdEZl7YZNcM3Dk
iCRjUKetYRJ8EVgXVArJuOgAzyeN6GKrO+7+kJxVdWpbgrcCc0DSLxsJT1omj8JnJAW0EvMIQqoE
817zrOmdpeSGkZWgmTJYsSR6ZZF4zSgwGnHnVVTSjocH73ry75XdGOhzfZVJDiplQ1A3eNeouVHj
hBKF4Tt6YEvBQesoaLd6gr6npp/2ITWDhdvuWcDHhZGHMbLRRphcpSE/Yo43buGHLLlSBx4WsLdr
dSS33FTpwpdG/1AMKj/nHJ8l/5Pl8FJ40MQYNl7ufkXIbMhtxg/plPpr849JAVXxOJCbkYD8KGWp
FQGuq2XUnc+iqZ/FdrKRWMqBTBzAH11r9j+lXk6j+GIgzN8q/7SwV+zDCOQHZ0QvFmYR/2KTLq7Z
EmxEmzeFNMYhW9EbWFyQ6+0ZlEfTw/rLbahSg3aCwC+1pDW4zpuijwGLtb6hlU/PUR85I9D5NLGl
1V9A7eFrD4O4k3xZ24I476W1llFd9iLO9hUduG/V8dzdWTNr00rWMCYM7hU2K9Rcb0Q1E6UZyALS
T51OMHcVyn7ryqHkRpTBduYMDs+1LcAMUmAPmE3+w0H/2lFcmtOsjkR48gW2iVwl0lotzC/hUE8P
wknDCmKZPJPPWCqCo14bY/QR4tRU79vqLOC60QKLiI93Q5grbN6X5v60OcUzVQEUuFzI8/iPmB9d
HC6fgAW53RZfjQCshq0JJ6HINr5QJXLJtucOSAm8Eiq5xtkmoI4umgIKAZZf2DGvZ0/xK2qCdZeg
pXC0xhHc1AGVtmnd/p6JbGT6o4N/WMnQie+WIhQrVGBI5fZVRtSVhbjqCkNkH8XkNui6ai2RYHdN
d8NfWEE3uQRanDGkhH0uuclGt6yHG9dNaoHkSLS7ncx6/fjERdKayaEGRoH+xv5srrzHkyGPH86P
kYsksGczuwhwQJ9kcnzoZO244Pn9D3TGQpgWh3C/S15CsxGHxZnT0/3Kdj9VkF2xTPwWdmBaLwW/
zKgXuP5j9clDgpGAgTOgEi6YLfudnqZKyNBowDwwC5Ime7E3Eii1i4gsKfK5l/FPi2EOTc7xev5R
+i6z1xZfFCjlcqkwbkjLALeMXrDMxs5pGF7eTrivRPK8y1bEcqon/csvQevP3TRv8qsNMIE8ewKX
/aCx6a6fHdu5syJV2FAmena/wQElKTWHTUB8tXac6YY8fuv054WudfidCrEdsVh3Wv2UWBuZ8Wy6
g5WJcRW+axbcTAYVTFrQwzFWU79a1jYQ6qnSYxLVtK2rBxHvvQ8BsmV5q61cfcHNzSHZXu5i4HlY
2bLisvHtgVbCyG+mYmmNwBpJnwV60Bvb6YSv92FBJY/C4H0/PB/nZU0L4WT62uwCMxOvRGcGu9Fi
LZNdLIH7L9GZJKBz0BeQypJdWjjyzLUD/cpLze8MANPWHi4M+Nnb/C69xgY7gnsiAnW8QviXXzdT
KQ8g1XrPzIr0IMPs4SPr9LvEHV8c0cYf4A5DtI69M3Xunt3IqAaI0+qATwGBpaVQe4HXxV/7Inpw
X2JqWt81QklD7G3ivCiJ2GIGCDKzcYXpHIXyEoOtwOv+y9DKUrXXDlIoBgyTN9e5e/qfnPHZxlQl
nYpC4IhK2/cdmUcViNVsDhWmMrO3R87Y3O6CDtopKS4hvNUO009HINEUSIKK5bvAL9bxFfR70rjr
0hWTBP4HLC/RqawQcX//UJDglLed7+T7BRIkxaVNgS/cwC2eCjwKGfbZVW3ODABiWSxCHM1cMhPm
DrNs7TG9U3gcKws1VKV5BfXq+q46xAicxYw3p4YGM1mtV5of+QPBe9uRB8RIZzKiyy2w42Iz/m4m
WL0xBZ9XxoV59BjCSD6u9wRaxEbXfRr7UEQAznm4G7q5GQOKyubErpJjkj+wWU+tLnVvPhNwBzB6
mNw2vjnQTMzBiMVY/2bzXDbkR7oXD7qXQaxGZBgkuXpykfJui1/koy6HjuUCmjpY4i4ZZXj4Qnzc
egiUzsmATIfiO7usUt8bPmtyGCUkic6VTPA6NmTuhu18X8QE+LuLUtlPxOXOuD0I6ibyddv7u10R
SgqTiMyUR3xXJCU3RK+lz7qRVwLtfheB6K6GhbGV2iQ9enqarnQcC6t9UkmDodRmkQD+bDtqeJK8
HtX60jpui/Ux/udecALyk552HP74a64B9RZdr+0gN08HvVNVobHE9/km4Ccuypwmr1njwWhuFmu0
9qqcZjHzvPsc8VgaPGYswFS3T6DRe60/goCSDqRv1jGYxejnwzJJ1VrCB/gip+bPfAy0SRZMdTjY
YpZumFMX3a2fXaNITHK0rKO4SyzvZmuE7WntJVXLo+gatAdlzFyGakQHnCPnmvh/dtOUwEfrWf/h
z0k3km4Wrh+LICsWAYLR+SxzNmRQN0MPnndPRn4jiIf60tgkeDcRqveZgvXrmMrPdodZCzLFVRhG
bjPb7HWSlTqMYQrGW2EY9x2H/lNpDH2FOzYuJsTuEjUppmnrf7lfNmIoQXiukdLjV1du/aB2MR46
faCZb0PnUOx498EVk4nHSmpfnYGYkt5wWUyR935GKVBCp5t4/RR9NuyJiBnqiCBNjfHg0ilQWz/5
FOkYRa8CDeSp/2KdswsDji/kRMr17yl6vVNK5pjkXtJ+/KBt7TVKjJzw+eHUKUXtka/Z6R4wUKWa
VOQFcfmsSTi5keX3FbPDepSu8KFIXEvwTy5VD+dv9v0M3xT26DT2ljGKA34VHovYVx9uS2EiuZSC
0wxNAExdvs6AFHbAZtWXmXpAnS51B2plNvCW3dgefS2CtpvcrwHwQLGojcCS1F19tqcUri6quQzF
uZolnZdwYEEzGuOIxA5IGPbii3pSTPdN6dd8d9Pg1HI1sN3gALra0NJRMBdxsp5Je238mJJySBy4
NPQ6Qwgjtccek8zUEPiC+Wdp1p1AlKfJ0iloNAY4RkCA2aEi/R3euRWeg40ZhwsCWxanuZMNkGBT
n0MtEevUX+LcF2PcbyRe3WoVafgYK7Xl7RIy/jsimBcrYQRsjXBVffTGN7v0qityxRhna7iE/P4V
HI4ipYnydg0hoz/Vx+tFRgzgbQawoo1naJST9tLQcnxEVdD9YXRqkyI4j5dZ/7KCsXLzxbwAf+/o
XhtMmBO8ZC3h1Fc/9ArIO25kPRWqDSBtValrh9lsEsbhPr0jpDkBLGykcx5RDrurKmWBnQdZHz9O
AJwKzfRLkpjcSyMeDDUgrHFamNdgS85DXT4csE+I1i+S7/3ybvlXBcr/yw84ksv504Im/5s7KIbe
JizbuDTeKFDFh2uEGjVX5w1RKrhX4HXQ6xI/+e0xFW6x8CJwFHE0IMXr7T+ikW8K1TFu1Mel888t
0VEKh4UEKjNRq0uj1TqmUnaENowJDI8zrmLl1Nxrg2mXJMs3YMz9M81B3r3eNSsoMC6DQxMKl4DX
HVLa1iBwL7mWFgcOP26h8O8C54dTsg4oFe7nHpbAq/dz0kvnpVuegRDeHIZPhtpmrO4CSs6q/9pz
trUqvAtScZjrgmg+K8F7GxNih6aGRTc9qfBY4hb6Y6oyK5u5/BVzBgMEAVtyk8XrYxt4tWfVx9L+
/AF0qtkUgni11WqV9OljcKVsPU+v6TAh1g4LD02dwLaLdeyt2gys9cjp9X5gqiVLLo6fKvM06Q9V
Iies7O/7XmDx4MZUr3eLy/MYjZ9nVU8+tWNCYk+cOnBvpH6MQkEK0isi4n1suf+oj7BvVqf/tG1E
E0mSBv9k+NNijDEZwQ0uhxEUE2FLlvq6zCMxYJ7hAcn0+8sBfYC3ZqS5iNaCRfBSfHp2PSwMK3bK
+4BK3VdSpvBgZZV1fPCOSbU4l+D8EHJWrwnVR3qIphwXNtZ3oEnqHiMcxFf0a5YLxBI8Kp6aJBFC
xd2jEyctnmKRS1lMqwH1xfQ2fi1yzufKst1h7qYVbA4el4cWJfvmmfgUj3KvC5OApARoxzd8ys7x
nz99obio1wZtgQfIZnLH/dErOzDB10QZ23xE+i4kURfvTDKGg8m/uEGXaTNCXuWxqbeVV0rMzEw+
6nfmiSxBooc40a4213Ji3wt0aZhvfMF823b+4xffy7rbYbCGQThOpuKEcib/3CPUU1UBZQjuPqHM
8TGoeZCplFmmb6N0wDtWGwUnyfH0skdXnp79zyGvtuRjCCF/4cfXLKQq6u2y4vsAyNHJBaaoe46n
ilmGEq6AviDXFvptNtZBXussIUF0X2GpOL2kDidd9x6i7NtBgvu/p7DCjpgvofQaa4dM08uJRG4+
Iji1tCVarDLe84B90LmhEfDrLmCUjR4l26P/ImMUg3IdDalOpHVlqxb6VukX67ZvUcKW9AoBNonQ
7Z6sxdKyc5Gzw62XH6jt+R2sFEnlG1+i1EtNWPblSiFeCCB59wmgAzGg4DHX4c25L+M9GN6ArIAx
4c/ZIXPLlSc59D1OifKUb8zBnScgg/36LP5kPAZCW12YUnIX149tRrel+Lhn4ton0XcCflZtR4+d
cjBQGAjnozdppqaXOezrhNaBjcR4t9HlxXh8VAYfvdSPSRLJITDSo9fOIlhm1gaShpkLZawI6/yB
yYSrKDhGStsyO2aexbSEkz03+3KSH3RROq3Z5tvbmvwkVDl97i56mL/rVtFDftFuUJsHAh503575
tT4b+jNiJBBrM4MhOy5GY8PyhJr5KDG+VCx2pjmOTi6XUKQJPeGSArui79EdQwB45ejB2eP8ei4Z
3CZhhN+myCtRfOuM2r98WDlifUvfIFfUEA9oiOCnaY2LSZ5HSiUREI+rRIpEQJQIpztFVU90pBWq
XwACnaVpADY1W47zE92KieD2JNYCFlBpg/d4+stdKBpqFcIifoEtIlk9W32tmAzQD35ReIWqVbJ0
jFUCbdXR/dUJ7J0+mCtWC0mzd0jTIkRcOUnLCPhTTTkRnJPRFJ+a/ILbCQFRXJt6hdpZENYrj60L
pdViiLENqx9qJM5H5RYYsFUZqEOrjib/tuQZxqqOw5KxNr+bFFFvNR76u6RJsFyCxRm/xFK0qIfU
31vqKuaN1wQLATuJEnCElYo/Nr7o8GNm8etDJuE720OCrvHFUnSNFHTZ4FLCcFCMqG4MoYsfdvim
Fs4WZ73f6pg/Cy0XpNRodgABGFE38AmXI5JW/zTXJbO43R7dj/HZWE5EP3HcsznqjnMU56Mfvhr3
FNRFWts2lLk3OXTXTIe3JFcOtVEENwHa01bp1vb0gHThh5fFJabFWb1kxnPfj/Y37Z8WrgexLeBh
4xUm8oIPqqB8IWPaWSInK0csa+G6THL9FIY2obd3o24EaTxqpzLizXEcfH0Cd+Pmaqxk1W7zCQdi
0slH8dPrwcKZhfl+rie12UZe8LXCWf2bsUIv6lNoar8T//r1/lGEpNaMKZVtMtSqdF/qknF7LKAa
l2hklvNeKec6Fx7MPHT5pi/vifyAkCYUPMyGykI/ZyIXGh3enapviVbfkkjYPiJp6FR4o6K/I0i0
Cq5wwcpeiWQzvMjCChBQwlygvMLDm43zVVQo2CaFWRqJMyavlfKq3bv0OMgqWHkwfzRFkWKG+rM2
EmURCABfTHUJJJ9k+nC/3vKR6OJ9PyIfJeo/odMJRZ6uamIuQSiXzNqIgPYK/gEDPIWwl0ZONz1E
l5UYO21O8yOuDgJfTgNsHk4qs2dndRtjcXVE7JW7GI7AOvKz9sftN8+uKsLoy7RajGb6okfHwMw+
OaVc996v6Yo/H2Wu+XNUvAKea043YtrLVmHFgS2uTS8d+AlJOT6XmDsBqykR4TZnXchbEEvvUqB8
lbQaoegA3ONtSCvYP0JuosZUgyyEgd0wAIWrcWugDZvSqOQMbLFah9IVBpNPbO06wHgqyu8EAK0r
imLcDDG+bnTshj6SFuDkso1eXUEAmo+n99jhvYaNdniebdlsW3EmCoBkkz7qbWcL4rcN/kMnQUfR
ANnPzMakHHPxXoMA4stOeAV8dJrU1bUU3WfqncyfbzMZZIvJkIHcIokt976pFUl38vbCRRGfn74u
Zjkb675d2faurLuc+3xsS8r1JtRRSVndVBWKrHFAa8qaoBm9b0mYdchf7oCrqdmIbvsqMH74ajoA
Y9WzvZ/ldYQXquYjMlR2inYVTAkM5QIn57no43AlvHEKZvbw9d/BkHkLtbim9TyI6Lumm9zrmX21
zYDlRZmRXrMfN534psMylD4/K73Optan8fqg1GtBFYbQm0E4NrzDjwtG3kR5ZybldMawq3gTFTFk
aelU4N0WkhFMaCpZSyBE2YCOXqEvHTdkIx8TpE5mZ2qWeA/4o4oEYbwTeIeqD/8cIWpPmftShsUw
PcOx6ZW/SSSfeUnkdt6GVZDMM30qNst+RzLo7HGfgl0OyDwsXD90EyqjEcpL4IVtVuKYpiO3vTCY
VVY6O2djLy79hHZynB2v4qBplN00czR6/mpHKqyujQhaBZtDEBMpO6DXZpEtWtyO+5CSCWmI3ETD
jfTTPaKSAPw4HXf/++1KOC+6IF4Bm2i4D0A6TSUqfPrT8ZifHbGYlomSTV7cZj3AbLfovqNaRnsE
SNmOUxC0QGZGKS94fjLAx0dWCwcjy37k6UoIYuG0S4bgDgFEHz3P0iBmqeNcsTHCsLrsT1nJi4yN
KJ3V0eRdKd0WBHrEvaw5OBpW4v28r42YHCWaHThWTpIKEF7OJFNA9No/8r0OdvrbuR97gKXg//ui
F40T9eIrdUSrHGh+1iht7Suc3oPyX7vL9CMhom0bSPFMrpneSVEJou3Jd2XWxmSk7Z1dNjzJQlS4
JTlxpPeaxrCHZbuu8DsJwEa76Jlvo+zu/tdXmpcgGY2ntXS+bQvr4AjcAvqsztWZ5UlgmlvDfodK
UXBYDWfuprYJG4XuTE2aL/ynBM39UNBj+HYfrAxyQ5E2hFvdIzyFAnR6cmQsoYmn0FZh0P3/DkqS
9kderfQ8iR9AnRcpGqCYrdw9WZ1onK8NG706bBkbD09uHD9eVhGrIf/M9oqgOrSXdf3kIqCrg7wM
VcLeBNmDv6cpTqEVNdqKOT78ayZTrz+1DTNJP5xAZeXFhWJmnAGEscyK6rY/L3A40xmD6AknOZWO
r13ivmQpkLShvfBCvxt2kM5KieP5BX7mNSrWe0vHzvxsm0LJ5WwdndH0kC6oAjAFsXlI/eKt32GF
S/+Ae/pa0gTMLXBbS2Azq13IEie2ZSuF0gmXb7XJekHQLALYGb626LUHW2jP6vIt+cZ9/bPauj5j
utfbbrht7Hm2Pjqb8kKNdJvg1wKW0gq3Lw/2EGiYV/Ka4n6lRglcZ5He7GMlmVNDyas3gbuI4VzO
rhCbflR26aY3ik69CiKDqP+JsbYEys+AwXBijPpPfwZLbBFM0E7sxwqlnKUmP7nlRceUgRbqwgLV
MYtxJNmlMDhuSky/dPz75BT/M8odzVCvokTV3lNmkRmihGKkJvLKDeE6Zvljx7WZ/7oqpG7V5OB9
wjP2XlQu+pFDk/RpmZS0LejDxGNiZoxQQUsIjk0MNPGIrgac8rb0z2Cz8yH0Lm5sOhQ86FeZD2K2
yu9mujaZKgrrRVtUBMFPYmwbczIRs1YP5/CgTIqrVoBjJNRdhPTIgZgBHmfoSbVTYpG6mKklysu0
hp1/1N/8hDt4XVZX34DFH7Nc2AEV7Wq4KGYunXxorR/jDoJFdhVjm02to9poobbKAbOT/bXyqAM9
juxG8YigI5buR9MSTuAj1411dBknifF/NssJA3+8lmkKQmCo/i2ATFEe2595MyceuaxGXx5UXJW1
L1WJHHcTDLS+omt7sVLCxjLnHSqx6LU8PK71biaXMPscGae7q58rMGSOUqsZIWYNepRX+w6kqMLJ
LXB5fIHFEOtjnT/yYu1qFQqLBkJUhIiJ+NT/zb449kyylD96JBLZeKp+dQs8ytA/5PskIwNBCQDg
jiNFFy88XSwgQKe0yQdoLgUp8EHOIWEUQa3PGCWAoqoccPB846DLwYcYV3tihHsWfHWjoAZH8q52
mV3azB/MQ6Yg+Lwdupr2MNy+0PAdulCOSeLNqyirqAXHNYGqDmU3cK73GngGo4ij1aOFPGphTyTf
rgx05Ouz2LHkoOic4kSjqKa5IQj7KtHVZmQok3bAIV0TbRC+uAlLx8kCo79mLlIj6D+B+zrh1E6r
pDraMCYP6iQe+zzCJBUco5UH+FQwGs0WUnoMcYuCVd++w1YG3QBdFPH6C/HBrS7/5DuZ4TO1RrHM
IYnhKv6ZsbhoR6wJYSp7mIzdFjteOkZTjBAw4fYLHiAHEHxP9zHv9A10AiCClJsLVpVn1YtprSbP
6Jrnm4c7UrUp/B/VrLo2xUCMGULv4izaXOEYTdOvHVaxXUgvQrk5X76Co2l6uityNECXcYl/dRHN
C2lJ4Rjq9wf0lzu6uP+yutRmn7IjZf7ybTQ6AuJd1GVuyKFijta6zBvNd8yqKo86B1+lFn0pE2HT
mVn/kgT0wDPx4me7Teumhyw2/IFNYn+eYQTaMbS2R+AX1a0glT4gKfYSBBgdx/iyriYWaOeQzzaH
lE96TH1MGdWDOXJlShdPzz1dYYk+bkQNPjAQi+20hW800yPSRS8h3L6nEZLbYh+UknUqqHhagjXS
R7PoupjVQpdtH8VRe4Vd/ftKbvpp8K9FhtagwHhN2mktvAKVW5X7mWT9rVzohl3ws4bPVTsLL3Px
UMJ6nNVn+L4e4e7MI2QE3i67sGk1T812bb0JjLwjGxdsAm3Nk/KGnkRPse81gRSYUa6BN/Eo2vP4
pJq+5MRoLaEFfmdQ0X0rmH8YoVEvmiYk/tFU8Loe54fM5XGOODi01X/cSG3FMw63uwWbKsGqKv1M
6p1UFmfde6kaqzgM811Ppxmz1YMu5nz5gdxWl2NyCkUKhVPvrbPd3QcC8huE0WM/xjq1pMxQQ90x
vkl7qNRhm7s9wPg20graofYSqKj+1QVp02pXYKI1R0oHeKCN5h93PIQUaFI3v5abLQ3ngjpV4o/v
9sy9w0wK0Bpv5KsmmIcEotj6g6XMD/3KOIYZUZF/35cTQawQbM2eeqA8z/1kwChenUfwwr8aOp+f
Mri5eYC8fG615DAMEv7IYRbPy+QLjKhNuSt/u+tq+sod/MAifYH3zkcSR+iuJ74BRpzrCcB1U9Xx
CILnJcT/m6tcBHNpKPA7VsJEaxe7n/ynDN53BoOXo2FpKPpjVJcyFnqujGO8RVVTMnGEsQRVIUt1
WIwjoFQKYeKt3utiNMQWQu60pIsiHU5ZeojCw5mukbGvGHG3oDuCMfaDEerbjrVSBdsi8wZQRc0A
nIouAH7WHsqvAX9cY06ntTckkG9M8xzAvGAxJ6vGw8NBKsczwrFTZXo34UtiZT2tJypg1h1sjrh1
VAAREBMIMrEPbEtfXvg7nnzk97CTsW3bV1l5xCTDwXa0yYVID0Ga0rka1YJsdooeEfRriob6GmoE
GpWSrs7Bl5RpJ/lQ7o5LEmwcOT9idrVBZOf7CwBg+d3H6riHQ+aR8R6i/jyUFNg289g8ukSt7VBX
wApaLuWWhmiEZvC746MbynUTcjsaaVcLM6nAvjedqnDN1mHzRGri2HIp59kGh9p2EQrX2jq3LRJU
N7F9gGH9qEtQSzov7u6oXhFXRxdqt8lqXEkfGJ7B/RE5TrjDdjyF3914I/QECeqQGGNveCYKjnnQ
UzRQQpET5wxjxhOh3Af5cZ7qr4BWCwK62ux39Pt9SZDWgK7tYqs4pxOsh0X1cDYLqxYDR4TLGrge
XaCe3urZ84JXvSu8KYbAYBmcHpB20UPrembUk7ackvKwB6munrdRHmneuYUZfj6FCciLIsn8LAxW
yc8awr3HrNLY7NdJkb9FyQbhEkPf1rLon3jBaANaURyHldlKedUD+33I4grFPWk/MuqrtrNsZliL
RfIx4V8qYcFh1Wgx10RB+NPhuYw4+M/iLsVtfBQpkIFjahu9G0cf/NN5/+JSIUKo+3TdQCRp9+ih
jvtUHGy13zvJXRXNuV3xM//jkVCcURntDP7gOsYSWCPQy0rD7izM0i9gJzpiUjFJQkORV77vdtTg
RYLLtHxwDOTg7YXzXnB2yd/RzooVxeIRWxnES2pyb0vx9Gkdpt78Vn74O+ZRzFLwD4Y3Y+vgz+Tc
gZhV+vSimFP46yBWwoeIX2Ws1heh4NDJoyelpvPK/QWIXXzbc9IQtCuXxAxNQgnMuP9RA/Z1JHIt
Mt8piSzv2Fu6YxQfqbxfTRqGDIeKFY2tsKSP6xfq52hZ74gZHV6TPvO2cf2l9C30IlnlbyW14moG
eu89my+ZrC4jhd+/dj/b9njHhRvM21ZoI+EkA/Ps9XwT48D3Xwi4H0/7P0XxFrNLWfuKTJC2zg9w
aq3QIpLF/Kn2R0pj4e5iqM8XnZueMw7Qhd0/tf9OGr3Rvv/ZYnaRYq4KdaNHeNMHYvTSUrb6HRKx
skUdW4GnqzVoO30vg0PQoMx3ibjbXd9fjzwT3ncZhx37Jmyyy9LE3kXdHn8z+GRtQhyoydn3UPN0
LAMJ6kdj2QlzUL77Io8B9LwXNozcM7QRTxDJhD7il0bhornkCOPYN4ofhDCvPplSIWJnW4MIaB6m
9YrFk3ayG8+maQ3Ky1uHeZxiqf9XVnDXaL0K9jVJkTy/rxYpIuni4iISVe7SDpYLbat8lswn06II
OpkteyEGJ42JoEh4KhHoXXc5bm6UfTFoG0YKz13Akyd2zpnT/Tmceqxy3k7UrrREcc+dTPubsGFw
fCVTb2FfTSbLmvwyrhUU67ybN7YfbIintnrqPCF+yhWQlCOEC2x7kSgBkp2lUH8iFFTw5m77jE8S
3vF3reBLNySMWyQLxH3badq8/craDGN2wOgDTIHsF40E+xxjHhE179wQpwpRATehUdIWL4SNLuS2
UUx0s2+bshtiQKHGdFO7/dSQzoGIX+upTjAIN5a+MTRU9W/fFGUxxa2fyNaPlAURPqgEbExazvF/
wYbAwgrMxIh8yQKFjTex7kjOnAT2dHTjOhfd6pKwcTzrVjrlf4Rg8HfEgT/+hkR9Jv+AOalf6JX9
Uz++URhn+bfCaKmXf4JpMrp1YkDxXme+g1puBh9ER+jbduRmdotBmgbRrqVxpZou6apqGmJMs+44
jqGK+I+gLSOglqsrJUcJa5RR/Soe6A/tVKMqMd1VQmlFpbyMt3R9It/LC6+l3sUybu3rpGqb9x+X
ULBrkDXm0NqvqZNurLOR4r3x48SYRwr2f+/VPlVPar1BH+nE+avHepg7YWbowyBVBPaNJRotCQdT
3a2K0TYd34XQGlWqp55v868E2dAAFRoUFNW3klbiTrBvIU/XTVPpaUyc1j2Glj2iBjsGdowqWW9h
k18zQWYni+KIdLL8nUTtIwkQc0B4MRdfBt+5mYS+wC6q3HMXnB2k3GifjY0LZQCc7r8Ms7+4USeZ
3YH6CtXcCnUf0yIm2CZKa6bLT3/kqLVsZVwMeN3Vx6WyyYwMvIq2aq+Q5hdhc/Kd1es8uofmG66/
QhBuJYbhDqOfq2aCEkj4gJBnIqIY6s4c6NwqHMVUGC4GzO7wD3u0sa+9OxGkyq8UpqhvSWGjqery
OUcasRTiIUVJyrioC4eoCxz/9qpjW3tZWP7B1H2ngxWQkaPs8Y8Sf/Co1bdJgfMm0djvZxKP9CSS
B8S3LT8RQAj8UHSCLfcuGAvVOXblydWsOcr6nWXorIZR+QGU3JNrM7sk4stM52eXYRcp6Kd3d9vI
eLGyNbCBW5iLiKxCuemEzMk0qxdX3sRaHAawcVoOaY54cqEvzx7G5Yhuv+4FdnmJxM/NpSl2QbyE
CAI5IGZLMsg79rPmHvvTizhcqoNemH43E2sA3YY3M9DFs5A9MkaTDszVluA+p13mIueRu8GEja3+
yhbH3OC2HLsauU5in/lyCoDEcdIMfW7FcZi1dguys0z9ovwATBl8FPgbZLm75H/zeh39ZyVDcBXd
Pru8fsLGzxGi+AcKWwkEzltruiYoWWP1S7l+dGTbt3pWZQ2z6x6KsCkx70MWuKPZTrRPUBoH+qaA
dYBQ/nCcakhrv8wUMv76ACV63Z4eNG2UdPniAWpUmLW9zOo0Kvj8jDBEnfQkHW9cfM9OmoJD8Qdu
KhZvvXiopOw81A0iyA7qFmgkHAFCYHI433+QlRhQwxyISy3K0TlFabR1FLNAsZZBj3xdPH1rCF/6
ArQ7tmzpHtuBWsJNufJHyrQKyMp3aAUPjO3+8PVNYLElIP0EbFhoawfqiIZcpgA3sq+jG1/7urWX
VPPPnFIjsJb6Pocy2sdLZls/BF1y+8cML63CaGQUC4Klmt7N8cS7QRo0taX7NP56N4Tu3ouydXYz
LMgzgkK67qqc9pQfdFNiBnxjY/UuZRPaTp0vvglJWN7eFYzGtaMm99t4I9DzSTrhAaRd6lY/V/Ga
7mV11+Y5MCQ3uTVjg8Sry0ZENTmmiQu2e0yn0Lgh4gYoGKlkft7LzP2iK1fhpF4f1Rif7JyyDOAu
F9pSZ6XawRSaQde+AQ6sdcbZ92D+I/TRlh2I1kY96vi6ROUn/JcusLdkGoPIxiyr8dfiWVLF0RoX
CUmCkD7c+CU3mSSZWEUVzxhQbmvWBFa2t/jFyeAIpJRonpYa0PRWd+v+FuzKiqhGP/tZPZPuvLk5
/wmXdSHRU3e0RxhnI4/G4PiaUTD4LXaavL49YEICjw9En5M7Jz3blDlPSRi0gvh/FdKakDXBKvR+
7i6vsEdbMl/+dSJA6RriFVvIC68NLCiA8UBZCVIiGpZC2PJErsN3IOZENBfvyrF7wIPBwInnVFIj
mlmnTuZoSTUsXgJaxECNHQXlY/xmmFLTLsI9/AKWxOQ1Q9RToPvPdKHvroqm0Pl9b92DwtrWqRkQ
V/MWqNqMGsjJsUO3N40iid6m/q5aFynS5XX2PleDZYI4ACnuJ9FYJRnS1TqlX4DEtOy3SvFzEABe
PxZLM5vbS3AYxdlJCY5gv39K8pH0tTeLJS/FLEwO32i1jsJ32VXnIL9paYfu3OoA6bXOLLzzZ+88
ua8JcbBSZNYqbmmvsGHC4dtDBNvGI+GegS8ph2OtR1KhHxOs8So9I3/xdyqP+zM+8vybBwCgX4kp
X6dUUMBOWFUcSN+5oxP0d9qjf+8YP3msQqawKeAbtuwMN4gJKZmH+nx8Z7u33xaVo+goE2Kmq9tF
UmL80pVpSlAvStP/lAkInkVIpytWmkGIyBoAjFgMPGKqwAfmJ+EvEsmdTFlbVwZ/YJQliZIsWLZ0
ecWMy4+XprpIilCli591DGEb0hwKSyaLXID4QlZS+hlRudQWnzLY5s1/GxCYr45Jtr0AJuRyhC5x
VUIZMpcGBry0MzprxPSWtjp6ZdXoIvTP0lSKF/2EdGWQFEtgEhV3YV3619bRHoF1AyV75KoyrFrh
RBiKOWY6kLWewN4BUbFWYC7l5kiMW/CQCexfFosICODh3pz3M3Co4U0tsOVDgyTeEvAUltJAUlh6
r115jSGf5qmwVWyhRaI9XfoBQh5Nq/rUWipXuQpN85VAH/C+EJkw+kffmm95KH50ri6FBx9ARF4W
R+Y/1mLIAXfagurw6LxS4Wv+LAbQcYE+PnWYkvsLaeQDTXlq6x1MxoRDBCzZQHlwu7YhpQWvVRAZ
ssv4AN7qwrjf+nBiK+9aBaJ+e11yy8dtflsm44OYg+gxmmev5b1rYblfOwAM/LumpUXsOS1dsVIP
D4NSX5/h8I8kb4S6K3xzR18y98WNlRd5Kh0dteKx+RonD6QuyqDG+T+xk7+P+/PjFgXmRSzo4pgG
6bZZV2HmThGOlt/kVlgnIeVkeihnmsJQ+A6sjqP1gcXwFy8cO4zYIDsfMoJFm+lw7wnzUdQWI3i/
kfJOkEh2+1njpsLRr1TpFebVEeV3wtBup7LNO/27jWrGgY5rAqMGWiN5TD+66VOxY5HBK34iao9E
5v4GgCqUR3ket6cvzSsj9j03Rn9NaR/oynXNAD8gDRFQGNXAlxpUL01cx+PnzWi5UK+xrHpZmEhD
E72vrxne9Lz76q8lzmG4YwytBOzkBnb6GHp+oIbh8TdvMWoOV2KvXKyxAR5Vx/NXxh6/Qni0qfQZ
eb0ROS1AFHWSHwPuAR2VMJ17oEtchyufPgp0I4wioSm/+pMLPvETN4+EIHWTmI4hMqQhkLkqdj3M
hr1cXjqu1KF2Sp7mOwOpQOTrW9CAkd7LTBxVhdKxzF8hkdR98lgSGQ+yjdJcaMa7RKA/ahCbEzFb
+ZPVS6Fy8xwNNjbl5QFVKJS17itwON9Y9VcYqZV+AGvnquMrOwKLl4z0SB2NtpVDUjY3rzLyEG2V
opTogdK2VZsLj4/nDWIz45lS7Dh+gqWHZcdVLlgxdf895zcagyMu++Ar6aG+Wbi6HdgaBrrx2a2J
aIh36oyNql+lePlCQUKv2tc+LuvZRRLpxhoh77dsukVpc6a+Gt8/JWgERu7YGv6V+NuierT/cAkl
DmnH3nnpqvoots+ecpPha0K+7csfpIhmddGwbo5fe6ylN9OO9inCWvLy/RAICo3gDGImkyHTpWi+
oTD/nWUX+7bZyVdHBhy4uL59M9YgvgWcChRJy3L5CglcXUyHDKo/PlBNltAgzYOankg7RxkJw2Rd
ud5zie4NV2NIrVVvxnDk4+BhiejaxYTuUFne2nfe4DH2xJJVE5xYylVrcQVxehLCzSiFb8KXiTS3
RLB7phq8EOp02eIyYzrFEbuuVSfL7ayNhZnyfEFBUMr/BJ6Y/KTsOmzWlwZnvnxmAENrSH/cuEOC
P2Lc1RNbtYrVxPgH/sbQP21bPnZFFyzcoc+U4ceGO2LcMotyRZHiSu6CqTNX9npLAjNW+Aypci0+
FHP/gCMu12S5s8cBvzF83B/UonTMXZcxEGHShyxjVjSifX6z8ynrLljOQkIRpMBPwZCcXBnDMld9
07ZDMVG4sySWR17khktZag2LpDMOFxqKLFyk8kQD0AyKjmj5dqcqc0hZjJm7GHJbXrQZDDIZb8QA
y06sWuDv2m5NdZeTpGmM0iGkVAS0c195IF+Bn7sQD3t5l6exMP6K4DPiVK1lYJ9EaUNuEtO+dwfF
sNfx3JzE+kuQLTklaASDiGWQunIcMkE/yKzO2KWxM6nlAPdDIjYbFFcrJsuyRljM0zrDYPpe4zwp
8v6suqkv6BBtMlL1Sw8maIZUEGk1pZSz7W+r3WJiNs1M5Vz+6bICLolji5DRMyJEFHAF2fHjmAJI
Sg3RHec+xK7u+PzK1nvCpnyzXDnp481I2x3xmMsEAKy3LlSErQ9SEwnIQNbDblADMjOE20bUKp0N
M6KXrnn4eLmgf3EbBT6Mk7Sa0LKo6afSdf7z+Wgnu5Y8fpwRrxnzmVJYM7MoBMlYXeLzAfIY5RQp
dRQEhR5wCnakEhwAKlkcawcp9dVNlCtBBNYj5CpW5pK2aLG4CHyj9JFQcVs51asXE2YYWZuSgE6Y
ubp20HJ3E+jufzBQiuFZnsi+EooXEE8oz85WsHe3Us1cFa6bNWnia07eg9+Qc5jYaC/6LnvgAXo7
VEWXcPLMxteIHF0kxJUqXJKCRWU+i051U02sBsvFtkZkcPcBYYB1lMvAWDySQSWvhqsh1AcJ1Ujz
lKP2NIbUBmD0uT2S+FqCCGTroK3mgi0vgaVTQj0RveMHo1+3qh7oIWmpkzgAPBt13JSDEX46gcp9
DQBLgGPoRDjmuZciAoqg3xAFIW/Bd3yBp5L2Gxsp0iWevHz3Z8Ki4mThKVV1RB9iOSYmZuPXUiUE
++5wKaiIVncS3vstIsFi4tNO/qqPQ5p9Pk3ARy3XHEJGQqvSeAJ3taiHaVS5vc2Jh7HIq1omfzlD
502qPcuG027BDJ87eYZz7fgRFbJ+K3P/Njs5s1RHTg0FO+kYjDQJ+6qGYXMlk+TKJLR8u+waTY0E
1LUp3PcuvcS2LZmmnNmDAnwGrLtXw18kCQLzcuUN3lLhKEyTbDJvdAyKTyDyisEAW5YrY+pyVTEW
/COOW89kJDboGbrmeJHKR09gIzZO/u/i+pwHwff+mxaNkwZkF5XPp4aZlp0VseBlkbzTis3TdzOM
LtI/Z5Drr1MFfO8xBwEjQ7IbRhG4BvzE7ki2jAIH72wWiej4FzE0uGDYLfCzDHcNkSeNR/VFlcE3
9FK3VfBSa4PFvh6a69O1qDNdIfJGmk22yeOCOyedl0NyTF90sGJG43PP3ywz+1U1H2rGRMKSiLo2
WnQcUNAxseawUQ7tPX29UdTP2dWgfdjZP0Tf4vHTmP+lT7fbKeRv3Ha9v1J1ssgi+jDbnSQmVQyv
l7Ob0mDC4o2M9s2YvEdaxX16qJDNCZJ9RN9lnIc9Lxyqj3IwAvQd5FNMDKGJtV2oIFtR6fuhi5gs
40OAKJMtubeoNp5is7EUIXUGjTMrnH51YcfaThdXmppAP9G/nvRLgDIeS5pWkI7noLRbLsG3xh0m
XwcVzIh7RYHPTKOSmFweenZnE1NiWqIRTPT8bpedAzJesMVznH/io6d11ogopKMBTudIby3x3KeQ
6BEREkW5NVO1HnQPJYzqtKpzDLkJdARSvBZRfzxwIC789zgULYXvGcBfIebdVw/dkSGhywQqo3yp
2HAY7Udlt3JxoQmsOx+Q8DZJGsU8CMDfJwGo0SPioX3B/Y7YkRYVULO8OsCFsfDt9nkhmy+RtalE
SuuiLjBCk6FjOUjCa04CGWS3DCybpT6azF58WmpN7IxWmqv4vvIqU9Fu/ZDPIzTdAERFet9ipeiV
T+Kgllra3q7hxaHYWY4r3HIQJMTqL2myi+zK4Bok6HaVOnK2ceyYm4MyVGHOY4fRBiXZKrUeDZMo
46/sg+eILmi+zAmxVzEYB3lubq6VzXh3DUX9ZRJo8DyJAxF1AjC5gnlDnJR+ONJyMN1+425GG/SW
qAel+/Kydi3lA5AvaL8/N4iuqp/nAszq2XED4USyX9sUy3ozatzxR3bCx5+CoOLOPU/+ZBsY8kb0
7KPv6rrhugM1VboWW2RH5lFXA4dWAEd3tdsN4nDGycmsF6MeDRj4eCYDH/KotaXGi1NbOTri/50t
2dVbEcrRIQu+Twr2D5CXWN1/wyHfJPAk1Z1NXtmZpCzJd/cAmdEvIPXLSpp5rPvATuh5LRDheBBG
4mwhBe4Nnb6RjvEdtIziMFi/obYp5TSYvMfmBFcj3nMEJWNAFYJAf0cFEAbKZ8TrEdCP5ABhh5Kw
QWxB2dakpjLPlB1TVSPG8kQ7AKUdlfl0Jhafhyv/sda/bERNTq9dPjDS8fyPME6AI5GmJp9liVQ5
ArnReD3wCyqKR6+1xknaoscCOKbxp6e7fSV0dX2OQ9zREhurLpBkoyAT+O7PHTyZdmKT2PC3n8ct
XxdGpXBrmSqmcIc7uaqvTl2fJqgJYyQGwd3ZN04JbqVu/xko04S85mOD1I3onST0D+y1STcAuf5W
GIQ41W5ZeBf4xIZZcCE1SAJrNdxCPij0LR6+RBCJh4EpaByTliEZ+kzMGbIhVyw5/C9zg9+KFSGg
zpVOHueSO3//bQ/DqvUdQrlR1uYsJ8i+mf3FwNdOl8ZjaMNzLzFqTdMEQ267259rfJ/hHuCKo4w+
4omddB674AIADitXjz8MjwudhX7DCsc4K2SYo5u+cZxrYkVFjr+jWTmxcWZuWTTFZex26t8/th8e
UZ7po4hbC7r/gF5qGQAqUWTX8xD9dxNyLkr0+J95RZDeO/tbDwacALwiiWK809AWwwlBcSjajTwg
qfFY+4uyg6yl83KJ05G1edQOpnBej6acmUA871LGmFVvf3kjSFnqL4wW3LC71r3Wbg+SNdI/58Hg
VUTDuC9KSs9Gt3Jd0TrN+wRpaifdjA8KMdHyxOBvkDDNp9rJKyFbUTwwhoQJxsBf7la7g5VPDjAS
IG5He5WQwaxRqbflzlPAq9Kqc3za56kSx6Al9S6Vlilc+o9keuMQfj98ZI3+I/tXxcbDKyFFCSRM
mMg9sJ5K4igk7qoUm0TcFIwJy1dCXJ794eHSOvJgXwgNm6k2NiaCah8DkD9EGRs+o1Y4YoMBPlX8
7wi2D4sV8yZLqfBYo+Am5qJNi8VZreiuULrWIeQFu+wp6ZnqnUUojSyO2BMiXch+amajx0DA62wX
StgaLKo2EWu0ihttBZBi6jo9EYH8Iz6ZLTvgKfbpyBYyh69ghLKQi4gGWOp8gL1HS5xNrLBZ7V9d
3g46VAy25nYquuanLfCDhT+R2ojlXhh+WyikhCcc70Myptb2IaM8KUgEn68Hb2DRiAkAqdfQl9zy
eP/KnYB0HT0KCZxQC3xuHZ7wpLpQlun6pTT4ieWFr9maza7vNX44i9qhLTO53QwIUu0FOt0E/Ti3
tmmfVkx3/hH7/hBo93/eeZeQbiG4BJLG9FIzsUwQ135ALXZL35AKtAHS5mYnjSE1GsAiAIdmBeEM
pCkX6Er33LXsDP/V6Wwg2aw6duaAUfdHXHsyisD2zgHAXbkodqSSVgVIBBexUhj49ffUH9H5QEXs
q1KisBTcoXetEg6Nu81xvkJfTfbMYkoi3lvyxjLheX6bFAsn43srIlXcHXAE3n2JctxboLdvI6KU
34iTnP5OgVq9VgVqGGvRYXBUKoNG5gUnI4dG01QxUGwOXRKWAh2S4tS7D4RsvKPWSIo4qAUVFsbW
4EMt4UHEx2nqC5kA/zMGkOvAQ/ZWDG/Verb5W9IGRV7P98Ht1LNV3fjqcrDGdqA91LyQgyLmpWhN
ROg2Y1kcyAp/9frY6Ir7dPtrXLvQPM+nys8y2OLhS1eQB8GFe/z92tkCmpUpIf19dtv8dsYrWTLy
9QSpZtN6SFxfnBw/nGfHNiB7vZO322rYQsoSf7xT233G4tDVRde7n6uyh8xwzFmV1hFxNG0BIwJ9
tjIRw075wQ1l0ZlVkcz6cUq4naWAOmgbL2PSyoy1i62BcJblk7reTnzWlPLndffH85dt1iajMcOr
+CeaS6Pwr6TwHJ5qRywF2OYdxPHaf7wbP7sp7im2amr6Ogczn8/8v257z2NSSu855+HrT7NCPZcN
URjLndPOcAlGXRKQWxT6tjKkD6C6qgOF1LGOe39Mmpu9lFUlB9sz8cMX7PsgGp9hEgfXrLhEwOzx
cDURFRYXazGx2dB6SNFlFCFGV0vFXEK64EQbtqXMtwxIkRg0JAk5jS4j1jJM/wweCYrtPmTSoh5n
WYot5skTzca/OEwSDK4WhvapTe+MTBImqNs7H/y3+q58cloAaFbDT8F5wB3pJtd/3FgQtnCScc9d
UqMBMaAdUkbyUXVaJ5gC/GSdqtLyNSlaHUZu+zI7H1ZKY0fcT5ipUTtO2+h98lIF31POSieN3n+S
m9rjMDweb73ZjeSoOrLtGa+9r1RTsy04ecJCbFnQkx3+lhz9Cw/ttNClUgULlYC+YFBlZtPJxgI8
Xvn+G5pTCGlw3YAQMn5e/W9ypeL1GHUU/nlIUOKNO43eli64HxgrXI+XYz3waEGahLOOVZTnZgGU
eYtTOrE512BRqOJXaAccPdvR1OdeWIFD+kyy4nOPqmVqg9ghSEWzRke+GdNciClbK73+bk8/kQ15
1k64s9XYO2pmH4Td497+keyFr90ZYnBdeYSBs0tADTPP+Kk0HVD4I4OBab4Zd6l06uYZnMJ1x4sH
waqo6hBrqW7lWejVGuhDk3uTOxJuc6ExZwVFKOdvRQRYnoQjcVwb9yX85cOh32Vi6DDesqR0Fp+x
si5K8FvcbhKqoEc98mGNA/sfPpRSw66DupSxtcW7e11DVJXvfzYnxRzC5lB5EmzYJX1BoLy3gMeM
1InCXSM9J/ZR8i69oDEziQNkUwyNbppzncXoZIMjk5CcreTFkgLjnKqfoc4KXqqxDKyHt6s1ZwM3
dUqBUN9mtuCncI5K5oZTNO6pvHDvl1TXeJ4cc2LDbX4Mlrc6osXIaBvW1pr6VKviRkl1yf6d31XX
tl9VFdDX+PMebjAODCmW1V09QPBIom+1cjfJPxmdqEz/M0xCoNN0DQHp+aSH4lMGvQZkT32yggNA
EHVz+HZV9YWzStzxH9VwqyXqp/4iYWR1rDovz603f9LTyFhgNSbnI12KK9N7gs4t8/qecPLfyDeE
+tBO0ayiY8JoQJ5TeKTm2RD4aH5pMG7abAMkDruGplq8O1+rcds9dqHJ/DfnuoohmGr8//xxKWf8
/NgH2DQL1pOu/Ti5q0l6bqgDlmS0BWcOUZEcJzpEGpobZL9ZI8R6XHMaE+rPFZKkE5QiUU19k/Z9
66ZW1TViW0FvtONaU5AX6yxNpG8N5GpT1WNnX5kPB9O3dKbghakBWJKApSajRLsQ/RurS4wUM5qU
PjhWNoppL4rA3S53KDEAudjurrH+RDltcRJDNKp2QDJl77YgYIhOB8yIuEFsdt39QWIVX/0H3Ob6
BGFqUACPCkS7PXl3HyPG2qtCIo1x6+Mr87o3+ZKL9BlH6XG0e/RZDikl/7IYWPhkwyX3Hlo47vzn
+pz+ntC8jfg7CiHR79YyY92h/YjpeHyEKsuIgmOvWisa+6WOcWr6ULiBDKIMC8akzCEgVwRywJkT
gJ2a4Hi4KFk+a28Nu17r4lE41857CAJepme6dwUnzJSmaayYYPeBdfWJHpuwHA6BmsLh5I+F21My
f30w9uG6ExGC6D5jErvViuTO4r0Y+IZQc1P4okt/f4+daKl7AzyFxtiRnX+1nr5FBAPJyUV9rpao
fRboszXZPZnCT4H6Jd2cxSgv4UOT/siT+3zOpKaoxhcHT2Xjs6qvVJIfZCxPm9673hMOQjCxSovT
brUE/BuNvZMiEpQc7BqrrcL73S4xRo7hIp0Cz0iyLfclQrESL/5HTPnUaX7QVu9g5S6JwSFXW/+v
1H6xJPFeVL8aSDEPUEMow4XnlBPL6A/oHC/EMJeGhEw0iE/MuB2qFBhQc+npuqD2CPT7fyC4NskJ
f3Hqm7CfoWB2iqsPvV/LMVxD2SSuZOgGqtRh2swrVfS70eHtueOkBc0hlf4tpQ2uWCWt/+yb4ho1
Xtw4qrPkW55jMfElYEmAlYC043tNyM5nQI0mQw/CKpSYzPu/iLMeDk/SMitJVPv/B7U4fFhUzprQ
eIvsG2S+NhuyTfez2tYCXhj+IyV9Cv7fweua7jnBn9v7lisdehcpbQjFOEYUTwG/05NB1ByxUp1d
VOM/wgg6uZMAGWCtqLJq56D2fQKNEdsdMpCoREYCLTcJfAb3B/WLTwddGnpSIgizFz5cHWuiNNYJ
ZeeHYNEC8Nsxc798+oK5Fkq96ZsNFydm4m3ROWlDvZgyEDh4Wd8AhGgGkrEEbpwTOSB+49/N66CX
mId31EgaBO1aygjLtt5zuX7ECD3JwyF2Wk6dUy/E6RYz12LaY7S7xmpY1vQKTggw9qgPp5PWn0QN
RAfKZKyVMRwW1iTqq0uvmf7y3bKZjTNWVM9EEyTsQrqnTsbCBhJWUPKAQK4NAvau8zEbcfZZmXBD
tAtFS/2/sRwOdWszNrMLW55WhMM5eIruBIahHkRLuYzSoZyO5sWlWT0SRZsusWFDHiev/db1QQgx
KRA8cVqTDYUxfjUSBBHKIwCuPsf9DgBQFCqyx9GRCtISelC793zGLUofIxG0TQlGo++gjSwj6U64
tHzJI8Mp3zAZna0SKbVCGLBmNAz5I8iU7LLhxlcfp6XidElih1+VL/uUigiVaGyanW6A9yT96T35
gT7EeT5RoaZUJP+RMDrWhr7+Z9LPt1uI0KIb0vLN44DPchTcjsym+8Qc11m9bNTdiHdR3lVS2WvE
ZyN4yEGqOgRXj8PsbrrKNZGT2X/ejTACnKdEJnVi/Yi7gicKAy11b+nETS6uuWQXG9Kf7SzMwvgZ
FfwrMWaWBF5axtHSGJ36OQaMAEj9BgeqjIxoRy+1ihcx5n8R9k1Ajc3w4kFhHZFx6jnCAy2n+onQ
0jCOFLUIOJ3RDjNCy9zjviYTIHC4E7UGRGguPQfncv2gCBWIgaLSl0oi7ynJ7/emx5AC8ICgnr+T
9E1Ap1zA8OdEXmqwHCf+V55hlu1AnDyafx89KO94FJCYm8FyMg1bw8q4R9xOS2DZXIcRXKPASC+H
iQHp1kzaGW2OI4WYgGzyy4BZM8T9j7DyMVrWsmS6EnOconIhmFAMfwKRlSS+Tbw64yG555skwgOD
pxtNv5n+j21dTHOiQMdLVoZdOJIXf3s1yEW0VHRDqDV2t+VIVO231sSGNfwwTAMBEQOrjDibPgEK
SWfh++eJidkou/84jI/HyYRUTtoAjwDWo2UR+8ASREr1gfXi7QN77zibVlIH+lulJmbAFEupdphM
Y2MEty0aa/4q9US20X0ETm6tjGBVVsRUfO4UY3XK5reJAl0oECC9bSJekcUqPCQ456Pn5Uudv9ir
ApEvJfBnVBF9alUVbqzyEWLlFzojqoWl5exUn01yKmjr3olTDgypOFfo1D+MyudNWiXM2yBwiBhk
afm3PSn1fHLShQYrnwZ+gFLKbd7BC8ZR2Pby5Xhh6cVS8SFCWeFjjEIMGELzVdWAX9Clz62HPkLy
i+xaE+AgA16LqO9tgnk6mYyfmjnlsa54MhUHit7h2mQvT/6BzifCzXncJ290TWV8Iu67aqVJ1XsO
anPzFrO2U90JhWlx5vmuCtwNR82BVtYU+lPiTbvy+CNYZQg++nLkBRnZFS1qt8CsSgkrlBU5KH9O
n5NZyhUjDLBVBzaDYIqhQsTiDhOWH76z3ycHZg4Krci3s4cJdFEmmUO4ZIB2ugC+fT39FNK4YRSE
odMVyEg5ckA2JBCexby3T10hsssgb9GqiQekXBEExCUY0GM8+XtJkFUZtIL1QV9nG7Bt3qczwQkR
uaAD6/oXJHDBTBk1b7c7Hb1t4LXtDiYja6grgSvtwY/W7diQMEVf7nWREyt+zYDG6QtotJyR6Ct1
jSqpcnVa4A7nCl67G330LA97PEaIZz5GluK2rHLROVcJ4Zuht/BIXd9zoCPL6B/hhMIaLdbrhvGH
xxJbtbXF+15Rp6SB21eiy+xFTAHSuHGXuoaL/MU9ChKD541avTccQXEKlmEH0NkpmGUQe2BwyUC/
2NgzP8cxELC12Zw0dnXxdaCA4/pxPgMskJv7i7XPyebusyKDvnHH5CnLjwiT22Tg715DMypDMFOW
kL/5YLwQZ2pPx+zC4x9qylW2P8VVm9C7imao/TWJbExvojOP7kQUlrx0uKNP5EJd1tNZlX8Pl+F8
Ieq4T2XdvVxC/psEeCO4rFLMOnH6eoAqXQfJCRXVqCr1JpyQ3klM1TVkpNuV0nwzO6/qkyRQf6D5
eE83b5W7n7E1IF6/OvcWaCzARNOB1r23HBbF8qi+6REXfpafCSRgE5cwMi/GY6CaU6al3GqEyAd0
ep+gGFu65or7zicEOhUq2S1Z9+3QqRuSd3DBa95rhMfq3NkhgTI+lXooz0fLu7+pmA7WeURpYoT2
jS4cut7x13eMUY4fFyZndvIVt8lNfXvSIe+ciN34v9xO0cgnGJTHr0gAyWxnI2YGRCBT0I4uH43H
iFNoJC3asleXW70RTidOmApgDsroZVzGxBgKL85eWom5cpm4eFVDlo+d+tzkTajo5kuKHJ7Jg4QZ
mvhQf7uFMgMv6D9Rg2kQ8x3WB7gV8Ffeh8vCSnCc+MRwapXSm/qDw6gLR0Eds4qHhAunS7zll0EJ
O12nBaWnVWkg65O73eu0uavOViw3RVKw7HlYotku/7dj9wOw4egeVEmLP9KvGT+WUWKkM9Q5oJZR
SHHIezxuL2c1GBz9VWpW6KTgBrgIj3Gle9W13Q+fMo7zxbnZlZtg2oV9S8DgcnhMIXGeQRO9IJqQ
SDcYAD5RbkTCaSCayxvV/ecE45qNFD5oDWi0SDXwAG4YQBpofN/JKixDRUg0YubN26Gx6Q0/9v6p
PxETaYglQ1DStkBBLqcLweQwgF4RgEIe7cfXBW6DXBgyfV70K4MY0W6i/6Mb5iiK8BtguadH/hAt
mSNUUyXz1jv93wt9IwbqoQWL0XBjTuT8yqImXke2dlQXy8k3NlQQIjG4UOsnL3MOiQqFvK5QbnKs
df6/TKjYmQ/hYL/nXhacVF+YbgBzHaqG2U9jcZCyXmmDxzk5Xj0X1iVzJj8DFVRJf9Rhuu4NXZKs
SDUzwWGvP+Q2mzFWnedaJRsie5MTImT1YSCzK/P5QZ51IXPjA2i6O6jAAOmog18SIJGtV9Bzsjpq
FlNge+KA22wS7FVlU6sWXegRdEiuTY+yQjvgAgr+2wTiViozUhulL/nlJrVqIeIk/UHbDC3+M72B
HLV+rcv66gmmYGWye+BkYoopAxEzATTMw+UH54NnComUeQIRjfFJup1AGRnahnvTHADNgL7by0ZS
pkAthGpCzZ3MkeerGJKF3kGQqIDF1hgBGv7HBzdNFw54NETOjGJn1wj/HNE4K01fzlWUh8olsIqx
qjKIQOqSF0+gQX956FTbzbH+yC4vqvnpdAt6x3Xp2Xt9NnI5ZtVpD/VPWkMoZy+dr/peO+BFoSOi
Q4y2QS1euEo2qgYZxOjI0ETgAl/jF9toZNlIohlZuOsbXRbEV/C1fJiwQa3eOR/lVgSj2es8vTMt
5buQH58IYHkR1TdOxEoLJcHGbFkBqHrgsXRO6XDC84kKryZpmhBjed8i7nvAuSm5UvapAqdEfPUZ
xYr9Qf/XbQRXDC7uddnl7t4FMaqjmN46ptBva4Vfqy7DzrsfNIijBL36LKmWzWLe7z3A7C6RnHyI
ZtxAKAqtI1uY0986WDK1/iSs5JzIVag/HV/zf6+U6+GCyRX9WdWogLoaMvHfRraqsjkuTPVOIPlU
GUjvVbTj9Ab5TOaofZ4GmVioisk6KOOGOsfQ8CKYmn6Jl1WQYBhaAXYe4LjcXAoCR6ee6OW7ONX9
dFRnKrQytRQ+z4x4yJuFMCgycwdlal6KLSG2/vP+CMHwkE4hizOa3XAPIQE5ZgRe9IWEUj4mpQiL
lD1TE1Bc8nnJqi/sP21WcfWkgR3bEwc+pUH3ZZn4OP/GJa2eNoAympjd5OCi7xCgMYmth6H1/ts8
VSoOjApjK9kG1BHDWUtjfE9L8L7jlUs7d83hPuXyKgTEPuZ98dSKwV4LIEexFGAxxSBKX5AYCR7P
Wg2RH5vbdxcrpVZFzYPRHnGEt1yMbcbx+OiWi9b4e0MzGnYchO9YckmIB1upmwNMjQQ8w9KGnnZB
EyBdXwuG3Cq4z+R2LStq9cYfGXjRQHUuQLB4M6zGRy4dnxBUGAy0osixhmlI8bItepRYTWCKA2WG
jjc9Kj4xg9lY2mcgfvJjh16uUgJLHBrg9W0gp6ha/emFyghdNiUI+0h8hdlF58DXJuIUtxL7qjBJ
il/2ggWW9SjUD47J7kKkeNe0j1Ezf2VDslXnDYOAdRD8phynf7dHcBdSspFFdQpkwPdB8MV5m+ap
p5ay1ZbGHBqWaCEwhbscIUR93msBXxi6U4nGjly1vMMennSefdESsDtCdHIdOeUezT6hoFzkY3Pi
MplwfmP5qZ5YImV5U0FxI9gsjZIBRmuUzr6ZMju0ajCE7BSHQW5PpMlkD4DfbbaEvzjYASWp1NFw
4P3avOpVdFYCJXOt4Pym9NKqxrUcOlFM0b88akgg9q5VPVcSh43xgQ36SrjLpcZ1usBI9HHAYXO4
MmVVBaRfcKHcR1rBRo0LZpRlzuTAPp7nUd5VKNrpDfzL5YInLYP5RN1/woWrBeu1RxHaNBQN3r3p
YD2TuGuk2klSJHPzPOYf/NZWdLg5vntnw8jVZbdm5uym31Ip0SYmt0LjZZK6kbsM+pgZcgU7OFiF
EFMcLxaAHofJmLswZrACP/5+miRzIngoJXUiSr0Q5HwRDjTOwUVM9i+4EFSOCIE5XH5581HVL03M
axJrsqkRJKsTo17cLBdrU6+gLnt0gfufnW+T1KjJIk0xKfmudMIjxjbjZH7/78+ABN8/Y9MbTzdn
Rp5cnfU+mwp+j1p00w668WG7TUw2mkl5+yC7LqVNYSMIbr0agKQtzkVp8vCxDuNC7R30V3N/+aAo
pU/QSn1yHjxEwWrl/sDAgIuX2bPKyKEvNfdmQjND9smRhcnTd6y1VCU48XbSuwlA/8NHM/2S5iFG
nIG4xKN3Jzd5CUTBh5+eLgTcIR8S/wYfHAJ4S3dJer3+qT/rK1oghJkMnofICMlQFJ/i9c1pZ/Zt
ViiWc5YXwimJadgRZv8vOkBW9DE6KHWikhRaCK1Py0Rlv8gfPmzhGpE2/zyDeU9CDsyJRtrOzijK
8sZLoktfRn2gDUt62NAasfRDIR3iKqptpv0Hptb9hEri+2wJfjcEZBEB4wZfwV3cefh85hfaRxtK
MlYlylOzF1QZS0/CD+7MUaKmXwh1elJTs8yRDNwhGN8rkcJp3TKC0KQI8f2QAey9oQk3Bt107ecN
p+k3JIqDADYZ9brYg8ybJfE9HA+dq3gH9z4R1rf6p/X8SGepcWIeFai1HwaCfawD0GYz9sTtXB7l
XJxVtb6C+8H2AjhzcH04w1zlWOhLZE8dxvGLl4KV1cm4vfDsdXHYH6+XptC7rt3wc5OvfIkZYzIk
o+cm7SKNtPzO9wVJn3Gm7qPSPk++qhDPgspwKKcgvk/6F5Jydba+vYIbR/0Uc1xdcoGw2OIF/+pP
dXBNNq4XVdH17tR3nOd5DpQ6mw5OLoyehYXQqncTNANDAVa2QclkEjm1DPolEodtIlqCzxvpko1D
OcthCwQP9kzH9ZXD4z5SmVEOqjwdGAiBHuGh3K+xtG4G8N4g4E6yhdcI8Jk5LmKBJsyYk/7bepcz
3n0ANCyyjDquXFlzaCnnYbgz5NbtHM9HAHzVW86u5MB+7ksoO+OV7NBbQxsQ9FiWD60N67c71pOt
8uIsw1gZrOMblgkvzskjE1YpcJjEYF4ui51Fw2l7Oq7RChe2LTZVC5aX4Rb6+b/2l+BnuvqdqFzy
NbMrceWbLYS2aIgdF8c7hBtX7b6gp0z1zuagKcEuJoLxRmGuq86TDjyL1Ui8kr4i8KxET/wUkgky
sd/bZm7E2YJce/MiT6vRxJtr0rkq6B/RpnwEEf0bicuV/CFjIR9+kOZkcVy8OtZGTKrrxqyAP/K3
KxQOGQR97UCdIaLjrChq1+8vzwFKz+mVPb6UYYSm8/7zEVYJcEgtXfKN9s0Oi1a4XY0uD9mxe9F0
/g5Z2o/Ob7r8rcG04sPzLoTUdex1yVFssH9RmBAdIVQIGsBclISTwoefSpEccXZPvNNDAp38LRTC
CbJC3eiGk6a2guLV53EpzwsvYNVgee1/Pr0BukAfJXCLDFhKVtYQXpgtFMO+HJeyMHKZFIPAcZzz
QoF1kbqdv6vQdIzWBxnZ2TjrKVu02G0xkpRGfLp7vZRs5jTjJ4an/NdMCHwHgpGAAwQHcIivrnN3
OuywKJFNtphAKgfsp5gCrPJWxNwutusWZLVXU28lQLgatnbUWnUSP0QHGZVU+xakqyYNAwt8FMUl
Z2m7T1MPNJ+otiJkKibqJe27XduqM+Hk2G1FBHYBq+RZ8wBrg7SlQYJUjyOdqZl+zDnn5HbL3UOZ
wzFaWZf5xA0sb8DWtQPnzxnI0PO4e86sNxNuDAMiCdQ77K0rQNM1LlKVjkwYloG/SQ9GB7frG3aw
qbcdjh01IUQX7bXtR4jIV/ZNGDDDqGcpsl14O8pUyr2hFVbqqao1aNSSe+SHNHmX0siuE8zYhwzn
NfGLFZr4usfrB/cZ2xP8IXJlzjgmu+ClSoPBft2qaKY2pQ5uNa4THCA5gqargWao9nf//NWR7z4A
QCsbKHAijtiHz80B7NVPP0H+6kIDqp+SQtIhgDL7dDKkVasM1/kd080qtlHidWkMnnPLxlk2q6NX
sNs1imc+OxfNTD8fXSas0/Johd/QXZCtP4h5k3bF16C/EiNjoaKzBN0SAHo65qY0yn3E4d2YJDPg
bE2r6mveTwdjLBnhsXFDiEa22FMBWhqHY0F2XmuIPrgvV1tPgVuzAD7g3JKq1aRsIoaKeFOE5ikQ
MfuzHHdlpik3z3/VsoVc/5OGykK90fYncWlTJJ+R6gd2wBUxsLYlEDsr2jGCRtT8tv9+wz2tlo3d
1u7qPMJK+yKhT93fV0QZ0MSqgaZeFUjeak47WR2Gx6iFSouAmHrPbWhluDoRQN2869UQthVElUKh
YCZXIneMjQkZpfb1tS0jBAdTZdqqw2HnqLWdpkB3VuQhX+/27ANfpHbLLg9namm+ToAA9O6uwn1+
Qjt8xdAu15dlQ2azvVSFKRvx+gACCSFLVuBisq45KvKWjF8lnOeBZONJgczBnPc36vF/q6NZgbKn
0gV5vtX0G0FKYmK2EtK1Eo9+XMrQKWbWqhBagwndGPFFMmVQeQZIp+HNxr8AW4+BKcs/2yM8LtLB
ehQuE6SpuJPIkJVWBv6U5SmFEHmR8aQnO6afg2CR3jToY3u8NMz5Fv9ooH5FgFN5vljlDIThAhzj
r2Z1FrSQinXf6hjH7LkzNL1pBNrg0DzxHwZFxafHr2qRCl13bOqFMI8OUmdj/DD96k/h8htiBKkv
0V1OSuvGUga69b3IUJoeSdqa+FuOAShZk8hitUqXmYIuITue1Au0oqT3I/frJ8Pq/cbfwvw8UFKC
i/ZJDN/jSda4KjXQsKJSvxDeRP+5ULstCdein+rJxbyrA2pF2xKKNa8zr2m76ysD7smTFcxZ6KhC
ggFylaqzFPOntmo8p6nBIpy35ZnUC7hPvvtgTkl3IS6FCeo0S3eV03pgwKWi6nPUv3GkhdBrgC8S
QWyM2PSRAS15u4BB+Q8If7EF/QtzxrhD3IbXKpw+4qvcJ81fS8K7yE4Ju0BCI/aidwCPnOtl5zW4
KcES6XDcc7HfeR2P4b4wTzF8ovo57ezjfBX/wt5ZGtL/5vIXBBa9YegmFIzP51JHD+vmzGUWqHVN
YsuxwCPoGka32OzN7a9Pdoq8BhZlibb5hC+Vk5CJZjDda5THyiN64F29m1TdsNhCHp1Svt3rOctm
qWC7sme8iLXGNHHFwoiMtQ4RHVW8Yvjba4dU/e7+JBArj5he69tKBq8+whv74A9FAj8hr154Irz9
6EIyd5CBlBZzMyS1VveeFHodaOJIBJ3cr/vdzIWRGZv8xtJ9Jl5BsrVUV0G7DPAjYGLuJugEIui/
suJhhptGlOao4SxIqa5S8Is1bLs4i/iuP9L2KiLJIaoylo690biDDGNfF+wnkkekIbs4h+q4vEe1
pK4ZqjIrFeLFGn6LTzd890R+ZK/sWp8Oz/1NVqSjxxghnKLOi1W6HzJ6NPjTynaqC2cX3x5aslER
OnxhiO4UFZgWXZkmCxySKYreTAlzvT0XNpeJdp/bLi8DmHyHmqGWHPDBeB9ahvjhBfp6bMuUIUMf
vxKP8aNuro5cXUTktiPN1pbP9uLqSvN4a+yDVoypjS9bHDmZDwJJvNQu57h9mGblS161WrQQ9uNx
c6S+GDaibYrnMapMnTIq7P1KmQtzMeylfma9MKxqwGdCcHVLcb2wTE04udSNhWJbJWzruk2tDLKl
xR4Gb7YMEiwq3GaLkl3UhZ7xe19Vq4cqp3Kpbgkkv/GGolYMrZ89WeQkVCxl6Pv9026+GdJNEf16
SpyK5fuBqhDQ6814WQe+ZvOviRJtFY0AE6wd8aaT5scFbV0bk6bLnZM4ZkOwO6+W//8K7CxQp+P2
C9wM0Ml8NBAC3LBkJByjJFCYxLQ1E4njXtjSIkDa52cVBbp0ucJTLQGXFb47TgNapfWsdtkCRJzu
FERHgBWVpy13it0uGgkkXmMO63U7/GOKE5lU5qtiXl1qDokPfWBXpF5xTCpRfjSbcrENCyxbtG2j
B9zM9MQJWHryVRpHjmQwC1OXyzdwIYbQpy9U8JObdZawHxvRSUmgsS3hjw9i3ypki2TOvODEFrwg
6JxLWKjxaRNBhw9FdUPaHaj2DZslTTiB9fZ5FBVTs1rSfJt1vPYXqIweXkraccg/uKONqGNzXH8Y
ia/AKJdqh6B0Bz4wvT/bpTfixBQ7SFe+HYtdcFCbnQ30wMYZyxzYRyonUSDDwmldJlLfvLoVOGx5
SDUXKzCWqid5fH3xNl5Fw+YQA51mjT7FZPpzsACK7Nr4f9589FUn2H0gajQfsB8u097BRd7nZ+r4
95+KA5Ih5q3IKY8GDGxJyCKQer6Ne74Ed55NtI+qC3AATP1wh7GXmcqnQU8CgK4Me7pMu1g4hbG2
Ou+8oxe3sJZPJ+cAVgdozritWzNsFXMtWjrac88Qau5RDpNlfUGauLqEmUneWn7saAaD43kejMtB
Pm+gPyhD6/3WFB4bZPN+iAS5DylqJBxGKyv8wOBuPGGU9FmNFDpwnc4d8rxjQJZFAmtD9TtpzsY8
ELIje8EOMaH8Noews7IlnWkAvbyfYRDf+e0nKGtyb5EgOqiNIMiK2BKW/h2qX4hNNI3KhqjlkfqN
qATMHWaA/UC3rNT1BJo+PY9mDGbK0q6C6d5sT6MQB8PvLGWeCigFXY5wTHJDvDp+K1sA+KTUE4IB
9R9SgoE7kdIb+3wieB9H/gIwZ1iGhGbf1LSMEdSk/yrERQazpWUqvb5/qWY8KoFhAGSmjEnOdP6R
29x/2E46tW4SFvPNGKDVu33wfQdiwH3nxOXXfqMDYNImWBYtCkowzUS0LNi0H3iCk0WPqLrPrYVd
xlkBKMajqtgZI5h4agGPTLH+NpMe5N1UJ6UNQgcLrTBJVVfy+trLz4eP/OySahIjwO2Xsc0EasVn
n9rVNjVcDRE3bta4adiytvQTwjPKxJVP2rBnpoDJvB8YoseVsk3Opm9aSTpjm5EYPCZfHjP7BZjU
K8GMXz/iV67aqmvbokX4Hmf1lv0HepTH+DAP+sVhGRP9FiR8Cjigk4EPBF2Er1c3DP0RqZcP+X01
Rfhq1L7Ev6eUFMXxzpmy0xUXh2oFRgZluhhy1B5atdZgjbQ9qJNr3Iyh1VAmPHhROrWBxCIzAcJq
WVCtkcSz113LMJrQs1atUAgpwBLBc9esO8J0iVVE/HnYXZ6DKKIKON+P0XcxngQxWIxxj8uXa4vA
xt9nR8ipvbrFmMLA00cKaAYAYEfZZQURTqR+FklOBrRvKcvlB8LEAzXDEsmosi5/p3HOvM4OQz2K
bcHBwG8AFf6lnxKtp90Y0UyxgKZrgUCMpSQwYpgygFr9rDt/j3CV6Iigpxe1tX7IWvJFzh4grIUj
Y6XsBFC/+UjAf4VI6KcVDZLT2+0faJjCZoVaXlHNyGPzezf3JeUFHglrkRueStisEGVhgL1BzTUm
MyBkzCfyDp1n4BNQTRNZ6rZgS0gGedsjQb76yzwq3RVyvP4GKQ6DzkzZTbwzg9hTPjo5s+Rw05vu
itWPmtES4+zelzSIsSn7Mk2BOhCbEqy98t41XnlqwzUkhp8y2qURb0PY8blHeX/dnP87my7nASoH
tgJobKoU87sK5FZR1u7ndwvbNOUyNU6PfxmpZ5weqI1NbxEG6kK3XeDH28dXJRSYruJ55rct6yWn
ZxrkLDoHLzNj0+Bl6laVxZECM7ojpN+FTx8uvbEyxdHo9L5cHNGFr9ZGddi9/zbKMidsl0aVL1Ks
zLigWOSo6NWfM8WfkP0eoAPkgsFlaDMfmoh1+NO2zeNyl3zSG9ZfsMqTiWsRZGP/0fnFRk8rFNdy
udWBE3w4SHKqFbkA1nSu8QDbPYpzdUzbKB94Kpo8nhvGZfAa5CRqTW4RkhM4gY6ZkGRctkWBp9Gr
/BUGG+xfy5nDBDUyYSczFuH5rSQce9sQqPHwCX2WSuz9N0ogHBX58p8S3LFDOgmbD5e7JnINxbdx
37Yzi3S94O940ERfkv5s4f7YLpaZJht7nZb43t0DzvKGoQslZL2qdbYWw3x80NvsmFAQ1TfVYFa5
APFVUPbbvRgcTWaJaXmJuLyd10wpgusdPOmSkd6/Ay8TXSCkXZ2rIPX35I3q3wG8TkKmb91m8npu
ekJRo0tuze/uZLVpkGxD2UTCIv7PKrejCLGgbd6qsF165QggoF/QDzWV0kynEGEwk5UrL5GBeTlO
pUX+/QYLHaHy3F2BTxQARIL1Lm/9gXr1/wu+GOyfNw6t/+b1flR6hY0fduK8HiwEukjEF0e+dDnI
D9eou836MQqv7sfqrejzv4i63voPPCPLUeYDQLC77MkLGOOZfXbI9hMiY58peko4LW3oha17Ex6w
IorUz0VPYyn1cxkU27wywy6YyXXrhH5xrcYQre0F6RfoZYFJlN9v7CO9/KTN/WTPlbsCirYLjDMq
zud9S+HGzggx5oN8XVUzo9XJlCEV2gRlW2LUPgp6USVTP65LhAQGLcpy5hznOk6whwV56pvrVARt
jC8b8shH8EO9Kiu/Ig6Q7tQVD0vFzf4ca7T1dOavPmzf4gBzVl6leCON2ZTEnOUsSMSqiIBpmsHH
mJhgx7O2AKo4QaYf1ap5AaMTfpmHA2y72rPY7J6AgQN/soevEEvV0Lkat/wrz8AR0jkDlKheLLhu
6fwKHbr7cXNajbxC6beOXAb3Fr4Hi/2kdw1tfAMeMBxnvHnOqvo69lmjtH3vJI/lbsBB9kFGXOKx
rBohTLtTtKRsGb0MPioc0VsoWdstuA4ZdnHbs74L692XtW89ZLzCfM5vHL7DMKbzHw7CU9bZtue1
VB/df8vAiTdbmSSDAfRT6v94lGkQC57h/hBtKufcNrwUEDn3saf1GpE93YHFNdFgIkDeB0y8v8tg
U2H6a4TnLCtj2djQyTh6QKFRNeH49IKpDwY2n69BKsICbvwUqGzMyhWuCPFqJ0lRTGuLGVmUb2NL
QOb/XDNZu+XcnWYPol8HTcFf6dVsIkDzlrukrvcJa+CFg7j6nOZVtcdttgcTCkPUj0RIMLtNyFKo
IpmftI0tS7fhfHD2QlfGA9XJUR42idN9xtI7TlwPpvCK1oTIkxljppUyYKQ/dHdXwvb4Cs0j6Azz
VeKH0BEP0IVXMhPZ6CQmJd/Ss/dNjpl2DSYSheTrSHsOdw8A8H/AsPmU4p1nhXCdk0p+7spFkGR3
QtIJFwz8CcD2TPfBFh67EinX37CdAOmSHgxXaCdyrDPtmBeIpu99eLhC+U4RYb1d8LGGKg/Vt2o2
B8cDOhTHUPCL6QtotyNRFtmlZvqFYT9ve9Xwbp9SxKqqwde3hIbK8cNamSYFWrhkXxMyFFZKEbQR
BMeh/dO8SJ3zlDtRgBmeNcLDK+ttRGH79s8n1cVD9Sjod+WBpG0/Atc3UyoW0XePWzTBCx6NP+CY
CCsvbk/i2uGdk9g2ghsCjme7SJv8gR+Ss0bC94RiVfSjDl4z4ANgvCKKYWNrhg8aQMuUo2/wOulB
H4DisVgXEfbDlnGidO8Vi5+l539yTJxFDAkrZF+QovvAgRfOd5dyDbkg7PeUfhjQPwOtZY+9OlMj
tEf4Xi8X9r4r95YQ+NGlmxz32MoYA7QDS7uiaamTFEzlIeD6VFHB5yrlkET6sYgjj6YGCuMkb90V
rnZMjJMeS3tSAbzfng5x2iJG07uRwrBXVzCIhOL4dms3HkBlf19hsWADBlyDxMxbmXGIbfIgZVty
XVH+FF+jw7UVpbK+EbVAUvzDvxfxNiv1JPCSOqTiRnjnzlqCVng99MMVMXxoiIRAokS6JnOyXGCo
PQr6RtQ2fgPoMiYWlGSe7zKZH34P8pwM/j/M7+oNKMiHl24w1aCurg7NiBM/fyxgFuylrfElvYK6
cr2lCPHkLBNs2eM/6slWniroUo2uN8ULhoWWIWySbovqEBllUhnHMGYydFwfQQaLuwUD49D/DekZ
oULi4hBvxIZesCKkh5fFb2EbVm8y7yuE9WFXD4zt5SamMgNnaZxaPsHkDJvHSSJpXwPbBsOERUC4
RgvD7XvUzWX2dgKL9nueZC3650m5gB9zg66/El9GHuyERGREgQYaCtksP5N4xssfV1/bmhft7x/3
F60ZX7PIpbE2K/X6hyflJ5dndmkTDInTkH3Qv+qVaB65ruO1slJIKKsOkDhmiFEHKx/6LBBH73Gk
0I4SrYIleS+P9efgIsfxvaoqsI6+mPCBVvD4DwUq98OVQ2CvdYwN53Mh2vf9/rq2Yi3UWEu/QaNe
uEIkrk4Bdaxy78gnOJcnRPE4R7owp+wboVFrz5eSipbyW3UB2Te92RXHh/UIXExEbZbAdP4w/r76
lz8jKw5QupfsQ6nc/7HVZljCh31nZxRShx2zD+nNZkmzXg6kgYO8/erJTgoAH8aOZhC1LnV81GUN
k5//3fMCZYtnlcviNUVx30mdNGo5A5ACGJ+DcqlsKeuWZoKsF2e4Cg8zx3opQPzCRVubZme3l3Ao
Qt8gcHTBbGe9WTX4uKYAHUW1tnp69cTK1hOkn8JJhaMQi9zpuglOgIQjmbCevwAYe2aSmIDYkkmE
WAU+TDtQWqffmzeDQRVeEBRFKdknzCDmJlCJ7NjK7TudeK2ApC4seUb6V0vEx2CbzV9cyI4L9v3o
tJ7pHoR58DL+fsAhQD80QxFW27UhWpieYIutRCCmJzGuby+C1fCBPMSGubjgvMi3/66bDIz0H/xJ
HuxOlX+U3up4TDv5mPflBt7kZ6IYGMFqs5QyPRVnlDqFPczfPCSYZG6DIpT5H+zi5kF/3KfyIF54
LrjnE7CJ3k/G7lbthIpiUzLduN2v42ZXvzDfMuCfohWvtTsNaYVWuCFkkLGN5J/5UD4Dd+eUrK+W
24Yl5JiUOR1yKS+ZrCNYvxU9waPxR4Cfe8jx+MX7RBVM3EoTXgtP+SsILgCPIqVnkpDteer+DV21
OotprAwT0GEbPw13cxfXRveKPI04h/b2bSprQiED4zOiKae+Jz6Irdasgexff7PRWG4jIwuzR9D7
maqe5TqwipbbB0FfporC6bJ8ND2SDQoR4d9qkIXnAK2hHLZC2yC/RXUXK1HBYEr6zYHL8lyqs5+i
CetWAmD251OuuUs6FklARkjto3jLP2T/Hyc1Y81Dm1Bu6o+m/f/uAq+VxbU22SOalYyqkGg/6QB5
inT6yp0RIqZV6FLWOMticNxZ2seDfqMpycUrHdi6vwp3gK1Hcy462zqgBsdtXC6PHJNrFcuZXdC/
OI9NTSgLhfeZKYvxNf5Rbaiye3NJVFW0wtjLkEtAI+Ield/GpYPpr39v+CR5RhPYT+Drq1sVqAgQ
OowEE0ZP5apOvt1T4H8atWS3nk5xAiqvINEMhSi2Gsia7C0pxLAz5zR8MRlMXl/Kk4rr7QyGQXt7
DlD9omTgCPT3sPDyvAhtp765Y1yFYjXmbmZPYhMbOqdrUnlxq1bh9KLoNrG4FLb/2q32sIQekatx
OG0QOiyTh2SteEnvBLeKQ4ioLJuI+3eKDB2Aph9c71TyNGK7XAJEFw3SdtU6fozd/nkpJeH2rFRM
bgadHds/QoMT+r9GDM38SGtYnVKqVBBNgjhl93v9fUdq+ro7NTyqGvqIw46q8SQyoxYXmxBCiAH+
AKrdrQcb4avM+ZjAENAn8grZDp/Dvc6xPh0S4ilz7ML4GfR5zx3piOvgrXudWKt+ErjAPm6/ry9j
u2fGeirbQrjgkFNyiePWJm4FYHZ8LMU+ocE7jgkvBL0Wp0yb/vc6WD15J9b03rIndbxa2x5HGKbj
5cknryCJEk05nr98UhX+twlYTaAedOZDEkRFyfQWrKnW5hzsWdnUINPUXde7NzRmYsjj+nWGPM0h
wvx7uarozFAvRj7Ev1VqmTXzXuXglgCQXAZBsiUXmPjGcujZi65nFgeOXLj0RVKAnpCp1/kHY4w+
SXPQ4OOBdo9e1OBVb5C8obM85Qgtn6AQbmHCv9cVvqsqbc323Cb/hSDl7X3HTCC0IarGztlAmdJd
/xObjexQZVSAUoaVcude5oDQoo8eR44hRUT3cj0M32XBR4CkP0dDsip6rbfXrheeaL1VQJmpP1Uc
VFzjKGLwBH1Vb7koYj/xXSbH0nIFkNmx88tw+MZlN0lN0FsZdrY1XBfzi+cPcppk9awEWzPrFvnR
aqbcvQFnrUXivRdNJpugKGTbRUrI5l7E6HRR1TRFbxt/O4FxPu7u7QaaVEqiSznJLLpxnqqZAYyU
LQZ0MbSrpsH9LeH/QIwc/DtTAd/O8/xWg3mIU+ptm5F0Ikq0P1GV+bl5erDJhFfybDlCDsjvjNPl
eOqUZ2HDrah4PKT9gO3EvbgdGEfsTzwjBImf6AnvFbeUMEgFYHtQC+BIHrg+HXXwBrYdwMP4RMvE
VZdP3S9FzWty3Na+lu+2WhaSWR+VwBPlXenKaZpAXlPtRrC3pM+4Kws+56Kcsd5QfHughwMHIGE8
Ny0TaEsBiNbim8WP6CfqlPCw2yLPRxS/oK8nGnA8+3gr4mUd+ajPxQucoqHcMU7lwaekbRO+fyjA
O1bTlRvGtcLJtZerb1izBVBc1TSvzJO5XTly2EhuLPBco11c8BIrF2kOG7lfA4oUIvgGWfhfQe1F
GFNgeqjaKyv/+fargJslzUFIpVtyoVtNOVUtr5TK+73AX1P0PWXJWyGB2tEJZv6NBYUBDlUOnSX2
W18aWdhMs6lq7jKL3LUmlTZi68LgGrwzk+UPNqqacyg+9kpMpC/NYecRWhneIpEMJR1uY6nyQG+D
l9pJ6V6TWMt1m8/chlmf+7DzdZIgNnSyifSVWxf/8DsZDaaSh92z8b4DDtYYH4Yb9BzQbvQvemTB
4UtcU50O0nyqinAZohlRMqyQyAQp2MPEvYYmOotCBSdMx1Tqw/YnAH1iScLTzRYjAz07/lEk6mps
i7W8qwvf64hhE/v+cWE+EjUtV4VfOKD0E7YoyyKARfxG0kQkcnpXRzBpHkkd1IID5eymjOvq5szZ
eLDmkxeGnPFlbnoi07NnGfLw1NcsFUnQ168ozDPdf0xbLO/S2Ebe4QqJBCrIoKiSrO/jfCuy++Be
ZFpYhxunzehi5WynUGue1ib2Cpy8ALhKiH8gs1HGqWh/7XrlDlxYQM5bxDpxNEQHs8PoLvt2SIwF
vV5QkLNthShAyAZr4cyWU3Myf79piLuMxFJNcneZVFqX/XcQiVUGPlKtoNOlsZhPagCKTcFl23SY
VkQsffgpvPWeQFmHoD3egRtz7IBW0OAAz1V1AuawuYhxIIxFLOUSFysR6oIHEXFFPOQuhT9GtSqZ
tkBwpatGL2bCoBycoiY72u9gHtMUA8xpWw+m9PxVXbCiDd5xsIbC4cz7JjD+OQ0a55zI28b39RRd
KkUF7BETJ73L0yBRHjTDQzGPEyKmjg0TXG3yOmFc31a3HmXwLQIezck9D4E7ABUYsL1Zhh5FKnWF
sPv251bnhriBhHs+gwHUXXGF2yxJY8E8inbmwOLCK4FmV0rua+qCSvjmLozbPYwJNIStgAI+zYPj
arCT5ManetRxaGr0t1mcyh9k4ICiFC1xPro/uExTsY1S3L3u1J7/R3iKnZ4jrcRSlP7IFXXcz9sz
bKsMOyK8QuGpJ70eGqA+C5NKLD0YSxkCtyBOs/0UiDIP/4mdVQrMtfXwdsU2vyKASj+pFW/IulRC
kLv8v9wc/bXJDq1L3zLpKpBgjMAYrwdD+jluaY79XN26YgYLHGQovQJXu8LFZwrVQYiDIUFIKQKM
XE1zybuV0mlQgxnZCsIJjUNw3LBFQLsYMdVMvaFpYtHxSkOmUjY5Q+PQdvQRj/PVFNEssxVyLkGb
iwh1aedx6zOSmw2OjKBmgGmS1eZ2WImZ3z+ikowLKA9NFbgJ2+HyVJmypP6uBmSYDzIYvGPT13Uj
t2AFIbrYyiTnA0hTeJ9+r9PdxNQsBPjicwhYU6tHs8Bapf3k4WwJezQ2KtFY41r96MbPBveSW641
MH8rWiAGcdCFXE0894kxVCcRPoavKr/ZpEButuYSzDtf8gJMlBnkc+fsiqQex4Wr5/m2ym/ntEsX
sHeEsWBZhJ8uCNlxskupDzpXnFFJcMDUD98YS00pdsuq8EVQLR1hB5p76TbKXuBBv+C4Z0puotiD
HbQScmJz0K3qJSKt4bpb9pHOgV8OJLfidNfSCWzyTdDYt77zLOojP8e8YKS4/fSHZnsFP/wgqmMt
XRThDy18zoGK9DZ80Aj9OsIb31C0N3y941QSIe7TSemy7p5SHAnAnOj9GFw8qol2zlBoC9o985ZQ
+NKRpsb4pyh7ctRzx4UUd+nw7BuVrwagRKyMa3KsX8TDmGoDW/EW6szg+aGLtVramisKbBwo9qP8
AaZ8eNLCJa+8akAgysxIT8ABc+QEcus+EJRQiyT0xWC2c5HGns4B7e7paHFk4EWJ/SNTiGkF7BGM
cuwumGcVPqHcBtAAAibVCG4Toc4oH056iASA00cdFRNJmqMoSKmven0TUgHF1QhUOuT/s58vhU2r
Wz/7sFnbC0oCnZiHO4aHIHn2I8Gln3cbT1RcNlaXxc3fsDVN0B8QOH/KoWnpzpDBjsbpZZ3RmbU0
GtOuHvgZiwA9rKJxgd2ZJShEibgsbFD14nY9dgLitTdI1h+MhK9D2e1En31wZ0KbUzmqtfw0S9dx
1KWd9PRSeWR5bLnnACLNqk3cxT2ghRC2V4VO5mcW5xB0w0r9O3Czan94G/VdruLtoAEQzFDo79rp
m875H6Ue33+Xdw3q4OsnPB372GXCo2P76qdTkqW2eO2xmzb1c3e8/JQrwF63Sm8rXzi91wc8+6FY
BIeGL8dpyG2/5R+36ynTrE6BaLthkzS7pBFCUitPLryeLAfeDuJM4GPqNfQP5aW4L/kmUPczkG4w
k5fRMcSLnlaSc/dQb+pkAspfz6ekJNvNoxFVRKXJaf9FsANUEOh6/tb4zAewK/GleiK/edqSA9LM
g3KW8VeTXfjyjGir0ImAbFOs/fo7iRIECdnF5lkFDBacNjQzvEBymkJh8f5cxdq2P0+Z8Rb4b1IL
oQNfuTkd0TmsnT7RBZMMXuh+mtelu86nU78rfnBNfYA1Vj+bQyXWj1p/WN9/qDfr+Hmm0zF82cHX
1YQBVaba3Z3vYU4p6n7BW7Iq3drUJr7YPLAohgZG+wrlVnGTf92DQ6qra2qjrhLKXuAARALPCKz3
9ZUaCVsrJrwfBGAQ8V8SjBXhcUD1kY7Cds2gfP1G7Zm1HfUPO4U9fuFIEHxdJw3CCwmgrVfd2RYW
rrrF+0VZks08Aywtkz3w9pFeVz9z6w332LjFEW1ixN6D96KiF6Ag4haL9/2D/cukfwt4R7M96jul
U5Wgcvy/Km+WzGqu6qQ7JZFWQuNYU2Zo6eqANiYzomyBkayBNILC0YAdfbQlspTda/aOcY4dknxJ
rcLKnIfWZqZLl4kha7HtA77t77QHx9jDXk2JQBUCKgPISlHM+qsUepPS8UeeH/GrJ4+hfoH/Xn1D
gTuwXFIWMvVUmL17BiG/npeKSkRVhbmNXOUzytEamd/fpwwYQKCvh+UI93n4gxNJ61x/AVtJPSRr
9aySvHsR9M89c0cWIvmPRPNGqQTV+hFP6SVx9YNDvfP2P3yzGn/8PjDSQLabCSAAGq/Zvvo/DXy2
YGuJqdYf/VZwKPc+NcaQAhGD27rImp3ACCmtNRaF2RfSCnIhYE3ilujcdaZrDAIpo1JXHR7k1vsz
yv2Hed1/Ugzl4Yff16oplxjDlTCVQJuaWnlbvhldYnHr9hmXT01lhAmlpqp68Spd/UdFP67vmVRd
LctOyeuZl5ZDc4s0Bl6+VIt5GXT9x1+b9y7OvTY/Tv1hd/DYgZbbQSJ+sozTFZpG1IX78SBofWRa
WP6V5k/mov/gNnHjRlXPygwyod1XW6FhiUXa0iSUtGhOLQ2TvEM/lJSLJzZTwPbKWzUTRnUYWv7L
+yvI2W+bx0IfiWII8F15qU9sMmyi5Ciy1EMifuSirXJjSRe3TOrJfyzrrtBXWC3YUBjtgYQrOndc
XbNU8GoSohbagKeUihAuNOEBCubcTRnBwEoTiCKrIlLvh1UK0pE0Z5mDGdRzLqPKV4Y0Fdqv9veY
LLRre+270t8kfPHECObuzIoDLF/IOTB48nwtho8Y9wJqjoz8uyhIRxe2zJbSjPd4BqaFtKCfcExE
TSFVSuy9jBGnhVN5A7frd3Kyd8iQb2is5udIVb00L/7oub6hOKurqPfsV38Bs6bVEGR+Du89Vg7T
AL9W+RbJ5zPLEAxkWT8XiSi5GE8DKeU6VnOYab1Yz/f65E5NcRiuZv82tJGrBV1++JhQgnGT018T
NsbgVgLbhV1kvoDBfcoslAbURXCM94NLWhcOiwNgKx/bWDPhPuUH9HqUN3p3WVkQC3viFh6xitPh
MXIsireCLk4eouUXsFTjmqZdZl667q31byuFQ+7cwBpmI3Hk2EeVHMWxPJZh312NMwiUBK78yDEV
2V4yo/Pmaa3JOITa0bNRO9ehzyS/fxuBQ6qEgRz71OEaBZ0KbZMChykrRRv1h/Fzn2MuGygtmUmJ
NZhyHxtEezxc62diM7TGhRnEU9XK0oOnPcmLGrixM6q7fVjbWDgNXuY5OQNE7UvqI7YVs49+deSc
BirUc2V5MPwGtKwb4oxS95XqJQbSFK8ytwYHPf9QTQHiZanFRI6DOVDMuPdxqaE4egdBAkeFnCsh
A6CCed46zKq+mAXvjgcA/Zq2X4fB6rkRJsnOioTkBKQvTJMIHT8+3sM/whNEJlTpxomhgKPXMtlr
xAoNC2mqFuBTD9fzAOOBtRgzh1nscJ7LbhXmDtgqFV/Qqc2g/UZwkWLarm3Yf/JkZUkpLBo+KXTZ
mNW+yL3NdiFF0iGsysYHN1Ma52l2XTrGDzNVtWrSnltqhMLhdzpaA4TI9dTNFh582dfLo8qQvixV
S0/iS4lQt3nCwco1HSa7+tFsH1gDT9fzQtOS8gVu4cABFPJaGWb23pgf4EQAN4sYFJa0868tX6tO
Fc+qVCZQ7Zez2fp+kLAqXo+56VPwFT1eLk3uSN1V7cV1y7KJwjGClagA7ELLvt9wG6filU0MAyub
HiiT82aWyPPOiv/elttqsOmB9ljit0ljNvoPKoyiDi/EvuuSFxYxaqMsc5WK1Q0m3DtM9XufHJQ5
SMQwEdug/IgSfRsHWyHB7GO3N/hvfnUxM1lk1f9VtqVwHqbX69b+VSI1FOpyt9EesYogWTRBJcnM
2SKrcnS6ou1ysOzuAeho4/ZbqdAx/5ZuW5ji4qWqkIn5O+jWuuB5SDfvoZG9CHl4JbhheDCTMr0q
sDscERJAhdSaMq/+ng4dg3nZqiNxVQSgPBcS5tK15avJ1piP2pi5e7qpTdKaXVxDn67Uw0EKHKzD
LTgAyFVpcJn31B0Zf3xW/qP4ZlHRKwjygIGJF8YydScZjY/BUcpP91U94BGdC1G4lZdifZPaW+Xb
ApHp4y3L+O/qHh36tw14YH/jI4PENaK9WGB6Nl23SKbv6HFir4jj51BPjZ02Se7x0k56Qi/4w/CO
FhKI3SgegH0eu9E8es6SkZ6CWI6aIwSAtHQrITn6n1RFyV/HtaI1RFawBAIM1VVfvO7U3ZIEE4VY
rIEwma2UHse91M/DOUbKrmbqciev7RbtmQPj7ejtUekBgsimsw4MRiq6X8Mpz4XitiTyVYQNECIE
MZCLetbgMocbhLAWwanruZFS88nOsMBdfT07tQ1pCgCU0rA7/ha3WN7yCppZCt0hb4HkI7VK5SVV
6UAJlyyeMNDpCohH21/4frE0pSsBdToygxALHEZ3uHwILhEmrNbUqkxmg3H/Gz5fy5MQc20Raq24
wrk0ixm1KSMDB9PqjDy1tbt4sDtZLO31odmg6Q3mL537lHvjDHObybZWOpv46XiLt0yTsUTAOjwE
truEs4KCzkZerIxukGDXuEin6lzdNABGZ0hfN0fi0lg2eVL+xy2mV9/cqCeCyDk7BnLViTAvQp0h
yKkrJdXP799nsorCOfhzmXqNwD1KwvN6tB//fBZb2YFvvICa1WvYGQ7u9l1/ozwSotjd+CumEBBU
p4cp2E3z0HsWbwoeu+qTKUPIyDdXs26DXqUX/xt2HQmeEXkDzFYxVu1M6EC0QsJRSVxsH2lyH3VT
ErEL2Avl9p3l5k1xbFcrXQ99nqvQCLyVMXmd85hi+enkFCu03xCfOmm2MONvdtl4tkxG8OlrMoLO
fx+ieSkJS0dWo4kIgToqY3M8xvFjYSAUQXuGSRczYHAWgfkhacqvRGrzay8mldjjsVClVlZwjKNO
aB4LHXhk5XvnP2ksT7xpPiVnWCUPj6OhTW/4yCtGDNGu8d+FowBKqX98hSu/5KZc8kef9g0MajUw
+rgtZxy6hd+Un5qi0UmPmKJJxaFTLLaG+pJlPvLgy6Afn6cfpbtNfJfEoNU4nncQvej6gxpeebFi
1YLhpKxL8mb32l1728sYxGNnOviFyehQkaBNGAPj5iijfz+RpQIVzqf/25Ao+weI3Px0LRsf41U0
y3jjDxhPDSjpEZGlUDxiOhPHZ7WI5iIMeL1QG3OdzDRyElGwBAw6GaPYVXrhDfG4TiM6lCfY8hbJ
8cY3TC8FuRAndbNEJwSdx6dQzkxaxsbEgn3IoxSHqCg7AzXS0sDQxMlsayNCAmmlGSTjhao+vyJC
yuwyvFK7upW13bA4/f1P+8U7ZSLirIpItk75cLi7+ppgZOZbo5Kcow5+sxZZwwVItICelM6RYWFu
acqh7twnQdm7Weg4wgtjrDdvoM49arYBhxcEqK4BkCkzOsBHfzXEbrEWMuYQ8bsZH3rCthl/bX/2
utZe47lyvkZ5DCfBKXJZTuLpaAfn2FUjIUHpT4mUiFZHTHN+Uf3PUQJ0OiUJqvmhYZMpuq0bOaYv
vLOFNEyGg6lNzAvcVp/FkDniqLYgOImFPvZap/Lfnt7gj7r4kNJOwB1mceof7W7cdeApcHh9pmjJ
HQZPM46M7XJZQw8bnDnJOOJaK864miunumpzbNOcZnnLPGk74wirABi5TihitcnLaOAmizGyqvAw
w022m7FXjiAtwn9/Xrs0jDwKb0ahJr9ePh7RBP9XIEnJuXleCowtdEy4UkMSSy0gJG1Pgt8iPrvL
/2kIgA+Hogmp9btkHkcQ6OHvlx4VRyE/mhVTujoU6/fBDiePob7q5zw+FKbt/c05ea2CpePZaVnV
vTU9x4VEPEAw23ZLZyrG133u4gFS5rvdjVabzk54zA+cprNwZNrLtsqFjljn9B8o3DfiLUKshuxQ
byRgZqDtI4X+eErQWpyEFUa3qNikNVb14Az5ljPR6OIglaAMcQ7EvXbSTZTZctc6i3GSLbpiRElg
tLZJmCe3BQgTAmKJFku4uk5SJbbUds4WCggHEJ+mNGSvmN/5j8n2/qgb8Z2GE9Zb7MUMvvL6VHLj
18LWM+ORcm4woTbqX6/Kkezna6HcwLfaP/Joe29xufPyqMFv8LVfGhs4fwep50+rJNlnuvARLGEq
FeGsprfdUpTQXQVl1PPCK0fv0QWEkMbFKzTHP+8gv//j7TGfSxdWjgQ2d9Ole4Q/hu1yjM9p1Hqa
3RfhfMFeY9dQwlQWO53WeEEQNz0mvolB7A1D2qzzYBS6zMAVbj0KQGYo/HuXt5J75w5LUlRN71w8
pQXsR8tg5rSll7ngkuWylilA4fbw6NN+H5/Mbj3aim46uUMTi81HhuXyRViNln3zdsnUSFFSUd2I
LLhHqtPDH8m2YGTwf41GuwNcJkxiKxXGEyxNTvLMb1D3uUyc5LuTOwr+hj1aHXrLoq7Im0KFicL7
XccAVnaqGiccNVdgQCd58C4jFFC4t4Vp/rl4bh9aPif1ltMgCdwnNrIw+gw75EhBvobzAa8HPFSV
S9cD/57VGV7pSQL4XzRm9tYQzyWuX52tHkgmRGltIMdT4BYs1FbV5iab7d6R8OHXe0UbM8fCTYQj
1O9BPIkjq9pgt7ev/Rh1IlgSzFd/B+KuazuPJKo7tCGFk+4KK1qObVvj0mFTcfP2Gis2bptzto8j
sVvYbV/68q9BZjzOkNbjapHL6pWvIa82Z3atyEbpfN7lPVoTuzH0YijHNR1JMTvIvtYfpXZwFSgG
oTdZ1esMmwjGYGxUfCxR4K2JB9v4G69RYNGoUPzPq93/Pi3IU70Lk5Bkwf+blls4WjhG6OJXcP3+
6YCNJlfFmg3zl3sAplAO8I1xowCoiZJOVlY8YIvYIgiAFpiJBHtjzjyfGAH/tol0wZvi/xJl9tST
6nVzIfL9DYO/mHkdL9YtFAG9IVgoSalg3jaHqJO1bgeRbfIRDuxpa9SesntScIpRgFPCA3JfNo4k
C+IFjG5kuztpfX18ejYazmFtrJ0wQcTTMZd2ZPS1dmlK/XFb1089CLN/4eqRJ9gLp/6UzasyKy6l
5QariGkjGxzerAAbmeqYl7667UufCK+6Ali74Tp/0JOaZCxQMTRt6Wv85sk4OyOViv15yinOCtl5
w/wDXP51DnbroxN/ZXJcE0aRixgdkrjKkjNMqrsZ3cJ+JT5gENASQ34w/+gZdlqbjVDoY4OWPcKV
AQTtNcu+zm8U5MHChsx1uUeGHKPsudG3+Q6Fw6EpWLp/AE0i4ZouzGOTkwqafNk1jwDAIEVjGpoc
bsTDIMaBMvoFrOGWhRfPmC5ch6dYuHUrRLOi6etKyQvXvADulC/XCXC6Drb/NRmL4Dl7yi0hefg8
FXETr8IlairznC86scbk1Pgnr0lUnP8KQaZimHzX8x8PJvrKSBwraMsL2Eww3NbEk5lY/O5SCD2d
XLLqTTfwieAtAboaVkwjSiex6esW9srSVK0Zhvn8ZTBhFADpuRMa9inwr336bF7KyHWNqgYsZKYw
ckR5/I84rnL1EpdoB0N2DBU7FLTwdhqi8INWgDl+lDPY1gGz18k5KdbvMYG7l3DJY2LyS0SQy8gJ
fLtBq3cxZJs1gW2qi8PCORGa6RanD9u/esvTNT45DTb9XYzlm0aiEfEWWq8W4bSXG4US9obxeUkx
lmoOzk5R29LuRx6q1eO2jooHhRYTbcle9jO7sBTm8im0X0neJfpq1YpVXNbKTFhlYHwvIMGhdugO
XUeNVCMF+jaj7JxH8xlsDE298T7h2SLjZA/rjDMvtMWWtKroUqTqpdWEBruTn4MdmJTrWPKViXaf
tCZLF4vmZpWsY92hndyPf/R+AyxI5MHeuBATj9VO3xqZsEMTLW+XmzPLxqy+0sr+L0kH7keemEEz
e6U4Y8tb21Sk14U/1z82acrpTDOTs/9E5Cnix4qW/0QXjTbLOeAWlvTLwMzDwXfVNCMIOmSSP41a
67AcukRXFoC1t482pQy9ymCWNVXByv5ZsUrH+DNJ6icOiaWIStL8yx1Wu54VN7M6qa7t3vaEM8f2
9/DyYVwzY9F5IsyDQNu8Z6tvT3lgC55fOgO/8sMeXVzLtyMx3BrAcjfFF0VM5+hdvhdD0urf85Xw
9f2yeJO8l6lJIQlK4brh1YpCMMWPcuU20yF5QiOkqTVCDcQYs/x6aiX776g8cVCT3lzCbFIVN/2Y
2Vs94y7F9fi3O2Teew0m+zVutNMFrqO5XbA+d9x3QoEDEw97g79qMHIrHrfT1lI4UozjvUUrysOQ
p1NnCI6kjfCUSbFhDtGRtxGXY62F1TU5vRXyxoz9m55qNXB2HQJa1rBd6a8ou9EyPHFY+Zkdd4XC
KB0ewmAXJQYJgXIw06187ZKVyRwyUSNR1eRH9oK9k1bUDwn5UH+hOJL3BX7dOWlbS0ZiyEXdQukt
TU8B4s01ckhEqdX7H2GxGWjSGz7clw+Qb5UEv2gD5AbQrhsDvE/jl5U4qhu9JAWH2M8hiBCJUPDB
stRcw45RNTnfmaXa1nSBhwRGrrdxQX7fMEMDdQQo7AjSydtLpHXdL9xQMMXxc9s5mUfdXpPCNU71
VjiKbH7/tTu+2bKJmLMJ929iLan77gTO4jUOo5i7omWzrjlb2ygkzs3SFUyoR8FVO+MTFjLfgaha
c77h3+pNdBBamR3CEo7+GtNfRe+B4mgrANbtfQ92W++sfvzvkkQsFHxCjAYKLhhJ2CLN+LMmptDf
DII6EtyvPYsn74JzZx+hLVISdBYNB1DtKMKGD+FiqJ4aSlW7gL5RrNo9Ag9qCTLDmS77Mo+WtX9l
8+tPg5q6fUG3SAPCDVskW4yBzV4lasXvYC48d/6wuhNlYEod0cxibavjQuzAhLRRaR+Xqq/lh7Ig
7sFFOiTL/VT5a4OMqD8yhK41r0ts0qJ9sNupBZ7vqvV5XMJdKvOCZd/eEEY3szekXjxCHtW2kWHg
jeHkJw3CT+ALv8sVofiyYLSDHkImIOYDoNtYQDV5WgbknF+tISwe7Ov2c9gYHv8MiAP0qk4FMrhc
uT7MpNQXc9hT2/IakgDqyyw6VXB3ryTSGmF4NLBMEbq0B5QMBGoeDeFFNAa8cJ8hy5vBAdmU1PXw
BLu81xddsoJWtNgXeaQM0p/svoG+pRCM+Ysuv7gIiJrMDg3aQ4azpWhMsPLItyq2tORSzc14ifeT
ajiYnTLzjUYc6DGa0/Dtf0hv7MfP/vKfECW1xFC7itxS+Rwn2iKYdbm7ZMc9tIGrK0t5X+c1NpRz
d0wmzIeoiQmHGNQZtDaCekJMphzXa/+ZPk0qjgUhhXWmEhCUEiiE3l+O1/VRP8J7WcSn4uBsNlYo
aOCLmf31MJBn4tGBXlCxN8uVx91XcoZ6hWYaMgyWqr/1e6ydtHsmmAm7413zIV5MTckwegtYLb1O
ZgKvEtWYbCaGv+71Bp947oLouTj5195c5JXSied/YM4DNKuu0ku7bkXAqvbICnwiY9msI7JTdcyV
XoIadJrzWMUg5DjbhadFGrjNwB5/gBYNcEIhjI1CkvtABBiciUFIRlrVGO/SYleHjJf0YWghxhvd
/ZxgzQktUEHaM1leRZSVzaGDgqfa80oRiyliuWGS2IumrYYNewtEgJYOBISSbE9TCdfLUKY36RRG
SQ639Uy4V5DXGAKzbtSwXW03V0N2+l82vtJn7DC52/cTFBeTLyaiTsm4RljS/csDQCeYDdR4SUsB
yR07XUzX3c+73r9EWxWmKbGdhs0YSj5ZicI5anTCuI7nVXIlUmvMpvFsl2qUMvEs83Aj2/6+IDd4
GRYylqwlNKqPN9i2fL7lffSt2Ih6Ypyxwec7xwuIVr0ecjrIh6C6jE3GJgnwI/hX8RRCYG1vHrMu
P6474Y4SIkZKGrQnTQmuxuu9b8DDqI622dKcb0LWRfAcIZyKkruyImZXHVmkGjE+A0BmGtTp9LP8
ZfZFSguisnjNhjNvwBzarOwo+egTBzxoSceDK1bKvp32bPxumaBA0H2tiHnzCiMSwFIsm1wAZudp
j4OwHKNl/dpPdg7m8+8cPwkr84wA6x/Yle4J2u5hQgbrycprMElXfYjLyG+bdmp1lqCORE2ED9Fv
+Z8sBQ9G1+xLvSfXhc1vK+V4YVex65Y8P54tElakSSX0drflLE9vM42LqBN0hNS9AHGAJrLe0KfH
Sn4buLWuaXg+RX5gytKYVM+kwmioWgU8YGeN7A8qIMJThZd0iFdGkNJBCErByx05hDsibo1U4ve6
SUCB7I6B7Dn2sStg8CR+Kc2H6EJV6hcIuetPiUJKNB2uYyOQmkoFTBNq1oZhl+dVomM0Q4NWBaer
FYnL3ZHkzPhf7xO/C7/2ahz4gaPaKDk61SdwZhPutF44P8Oo7ufGmFtgbMfdHxifxaeMKjfdvebR
w6ZEvnkt6N4TsW4ElYSyCz49x6TDO7w6SkYVdjIkYrk6QVJToT7ixrNGDgkgbi/4V+n/hkRsVNcC
KS8mNsIGI7aabAcNEqlkgptHla+7WvqiI/GdocoINm68S7O91DlvaYdkLv8csvi/bZwebyM6sqBF
z4ronuVsr5T0JwBoI3k+ee6Q3r/tUDUKGiaeW9mclsnxtIt+o5JWPthb3zYmzYZx9tw6owmuE1EP
TeJOMbMpfxQu2hfCm/sVM8srZF+gcRUzUHTgCtiJMLmrIRZypj/xSu5AKwG8wR67GnDwWMi2vIpX
y+KT43tuj2tWPUBXan34ousSzl/H5BnhSDUiIIcAr2p8CxDlKSQXwS4AH9kvs0+mlDUrqcq2odU3
qr9lHFCQ5aIgxV7CG6j7tXWIFrI39/bzaAEwSTefC9S1XrEYoMskv36Gcy2AuQ4SHou38wR4c4GV
kWmuo6wlp35fGjxeUfUj00vrUyyyjiI5Xs1f5QSPkuFkw3SMefURszqu0VJgw56zy9OqUIIMTyV7
X3y2Hpc47Vh1l2OoD0ER0Em8MZw3ejehsV3XBh2SGBl0t7iD4PSA59ryacWFCjAT+HR0hAoCzVX0
dzPNQFsDsVcK0o+ZvW1QMVk0b2jE25Pt3/0fO5Wao+qVeAbgCeFCliPe0Tj1wGnF5TNg9ee0eF4h
ajNfhzzcCmj+qZgF/V6XAD2jYQRZ2J5KVOazdjS8Emezvpk1vTXCaZ3woD1q5EqBPy93CaddT/VB
9f3uHXpKkrEMIBpiAll0qoQYkhnaQCmO+LRRGm4hCj4Q6fPFYeaPWhBX06DE0W65Wlr2fbHLHLkT
GcffXsf51hNbNuK2G5KwqhgaHnOGf6DUCiDfxLoZwjJE+UP0XG4sVqYhfS3PaR+G871UAUwlOf7O
8s/jLjFffXfY6pYbW4aETUehLMEXEEh45jeqZtcCe1Qdx53HIaDFx0lFZCe3elLa3sC/NlZX9TdZ
ZnWxXm01MfU1CLGXDga2Senro4X9HjYwF0pmB6jOtQxW74s928P/Kp3P7FKLsyNgmfy+onLAQMrJ
cgZVDTIYIQUoMO4M0fzKLw6etS5bI3lRir7MxwEJN2L4lJ4RTVYeB/rKkrMCu2BXk9F/Un6nTn8k
IanVgSrMFlSJMn1Nio+dOMI6NsaGIoYRtbB7HrpRpEITqYKev33889CbUkx3YEbrHKSbvhw4u1Kq
1B4A4vSoFpyaqqi/8Nrx5GMd1VagJCZKicjsEoyvCNmDdYY4m4pcquyZLGrCdeuTp1R5AiAyKDA7
uyszN0Wg/yA3NBwQYNrXsw2dHH5Nyl1WVcwXo1dqrsxM/DBwUEWPjHYln0DAVRcgktAIYBHabEll
4pCtdEiJ9GAFhyVWGMOZCKu6Q1VGh12RERdGx0ldHCeA5RbRqDadwiA6qfkwUCQ/gPk0ncMQHaia
q9iP9egyDplNvBmbSSHUd8e4rSAxP3WZVeESlwjRYQtggvlZTYXFuoLokkXuOUPy4paxVno9mj+w
EN7Heyd9CKZkMFaXA667iZoOTXpsJRoJ5zTIxN0S+FMDnGuzZP6tkzH71AQEEye/YAQDKIot39cZ
eSAXKUjq1ZbHQnYT5ZTO+TrEKtrXqljMVmcxpoDd0wXE0SJkQZEQpa3+yNo9JE5sm/lxRdMH82UA
8BrQf/qMantX8VAiZxztjY2p9SrNwn7xcuGNui+RI7et/bPNxKO04m0c/xfEtpHbP9Pk8tvuiU+v
+7m1f4DbwDAnVAFMUr09HvLcY0Lxx4N422RNWUQnTjnO0dRWaRDqqojp66BCcL1B66TyFo0JX5ws
jYbttRNsKSwNx0G86gdPytB9YUt4usRbKbBZGQsoqj8x3nUZXKZr5cluSaoBbNc7xp6oVXgGNbiv
XhkvRRovx4R779OEfiQisu3po75FbYifz/UIstr8eTnSAnW758dWqVI8RburHBZtdEnMx/QztiPe
H4pbzpnVA8dsgBwbiBhcn1AyX5TYVk5xO86Rd+a1m5DtfJEAn9/PPecPMYCluzNED/Yzdo0gr9Wb
bnq+SzeVcU20jWGZ3ZSPbjaGMWdckqfOQp3zF4rEbyudMUe8N18a0Ig0k+EycuRCvfPJXe2BMoG7
HlIM/LslbHh6o7qb+E6FAluYeqECVitULrePdf9k3afE+W6LYvPIRiKW7UM3p66tiw4G44qsYISa
5Cm308HiQiBw1x8rkt74R8AcNyqo7WOL35PFoDYGfH+lW7neY7pt6glyr8HNdTMYxAkAxUDccd2C
Re08w1I4ufpXdPuqJ3r1KzQ64thjyv6Eer4mQe6uME5t9BNs/8DwBKlO2P89OZl9epHl+2looOQS
+xt7Ju3byqfatAohtLlf2fLKk5SRTxy2VKhmJQ6yGTYPpdO0BDg/pSDkdr5DHCpaYTaLc2TnPBUS
7QG7KIoPmK1pKmxlgFDPGJ8exyVegTvDC1EEFiki38N6Rvr4cB+czWTgvFngRFMhCYXeTT3ayulZ
4C4TSZrJr58cAU/CH/S2YpCrtxXH4v5KAYHU1+kvGgNwc35tbnN9V0yib93vUN7PX20l0UorrOLL
gxjKSWt5/JBzHt998q96mX6IEmguLKmOMTLlQ7RJ4tyZR6ZmnL0oxGYY5qa6AylAnnUIO7NTzEYU
yIsKkG+5NsT6Rfdga2l/VNrOi07s4mzZyXp6n5QORv1caIi3YimYJ3IWWGt/letCSZ4gvXqDEiGD
rmHYkyBRwT3xtVeZLcGp380l5txCaxBKv12MOXwwtIiQ0tjstPUlP/JSGIPvqa10l28Etv1FeLJR
fyw4ecKAIO2FjWADd8dPH0/g56kgfJLrpFXLseBhrVB5wnsuX/bEMyaXN0dWb8Rlp2KJvLfjMT53
HvCuImrLmrT6kXSlK/9IRYULNvz94VQHiJqcuiISL2vnOavM1O7x6eCNxOjq5CYCSLGdds012sxa
kdc4NQNCmE11iH7ocAdYxbZBWYMaXPAAkgd0caSobItePXjjFcbxQKHT81NrixupDufFwNWxAJkn
pxFskABnKf1iD0iopADsrSx+RjrbyoVpKif9MA0WftAta6EgGp4NpBo3T/HAw7pkGR7DpaC1GV/w
XsuxPANjzvXO1NYhapoB+mfW8SSErhmGg5u2maYUAEC4DwU6rPjFXdiR6cXib4BKMz0+eysKtqlj
ebRtrYWV4BETnEE4/EH8zShj+fbYR9Zd1xQtk7AAypfgithBPoX3LloQLgq0FBWHUCgI2Llvgdo4
oX8FOrqp1Up5vr5+h9nE6detVkM+Cu0wbNalz9ThtrpWNNzIuRK5ZelvUUe3tEbPEgOkOcaRPTvw
xoqJJUN09LBOUD2kJMUrTeKpWYVLkiUPHXyo+zx2Bu8CWu4BWcAq6ECJFsyJ7vypkPvbMpxZh89m
5/GpehONjQVzSA9Ros8kjkAmwAzQuDL7osAdAHVrfAZtLCp1VB3i3gFuXNVnjL/nEKwbKHbBbs2F
BUEIamqCXPEkdOswCLI6Sj7pKkjfyYHCuho2U/PXWRleFmKrYOOPOq95N3Q5SZdJB955UP25VDGX
4yK+vG/5ho9GEJ/AD26u/iVzvPBx/pPNjAx8qHyYyH24VKkAVQTqggKeYvRfa1+TiAjsB2+qheSZ
0UZ3WXV6MfuY1YIdhDpltZums3Z2/sD8VGmE3ks+lRAy4jJKIuia8dL/WHlKcPeKgSWuM1b/d3M3
8t2U361AclatRXow8BffE5nTDK8E09clYqqtqbId8qah/X4D/0/x15Hokz/QdEbD+cPmzCp/d3af
sgvbYwjMO6IijsMcnRHRmYVslw7Qw8F8BDY9xNEYur+fUw1e5RHOs9mw601Ncdr8Um3FuMb01LhU
Jjlmk0UGirXuaOAWqLNDguOGd0LFgnOzeUFCzNPTpZmSEGuNFfFE2Xk5MKoi3AGWnolMxGrKTnsa
hLVG2ppWjrZLiwRdp7+MPDGESA+6CVcOIKnrqF45CYhR8JKli73LvDio6qB2OACA5/OaUqqwdxs5
Nh0O6616+i/747iol8gBQ2Bkwh6RvLVOdAKnJorTLbQNoQDzPBVeEOgUt/KUwN6nnA3+/Nf2E8Iw
9B7V+LDK8iSFVB9e5DQVgbxiyIoKjsSoEqIH66zLrL+Lo4HQtJlXYDUCGfM6fhUch1BWxAsS/c7m
ByNJq+atxfR9HPm5KkKHGYjmQaVGB771H3prfT4/ODs/eS16+Es31vEmaWM6zG/gm6B0MbGZAp+K
FtRuSNEs7Eafs0EtrTyMshVJ/akg4vpCnA5HxjbbB2exe0HcTmUQNJCb4/tWXryYrmqF1z+/rfT4
+D4OlVBl3iZl2MUmkempED9EtI09F5mAdw/oo0u3Qh1cMoULeOgw4fZp/Ds/zaonNZT31XDsPi/b
spIHQKPVv94m6ufGk8Qn9bOnCs2UoMcDzsmtnWV0gNCPJoq+vHOdeziy48buOyuiP11JYNbQ1w6g
QaFW0IEa3DnGM5tHa3jjG32RT50+fnSWjicZl2C0vGZewKXQobL7T18y9Iyw0xD91aij9+dVE2De
+zeFO+iTD6oJ/x3wa4zAgEj1BMbAT0Q9JhzC+YS36NIdlAPUgZMytX6iMPt7Y8Rx9yytZUZLI3YK
DqlGh+rIi40FVmqusDJMdS/b+X4HXDJsnIdB2u1VB3Uu2uoDTP/0YAQUVeYPsPvgWacy2xjlKoEY
mWVGlWmK27SzA39MZrPdMh7RyyWseevYT4y7dKyQPvobUEYVhM2fx6yvsWRdTOhGezaGHPTNfyj2
EVliUEQivJNqs1aj8LrfA38xOgBPS8IgqOkSWiw9ADCtMthCjJA6bKSJwgd1p4wz58r02IROUciz
DqRbrmqqszywhEVVHbHX21BlDkB27kdgWDUM2gf2/8OkVb95K3Ooli37V0sZZUGvgHzuUKTwmtR6
NTHKYLxuNqbZPZF/BSVXbFwyhMJ+nfRyBydkrXiN3vG7m/AFCrLSwCw1itqQBwhPZbXt4HEu+pKd
M/sqN7i0LkMidooen2qBEiItjGkV7pBhTnwYKPIhMl66JJTSLclkBl9EY0ttUErJH6mur1EXYfZP
8z7dv8rk9ot7EM0Qim67EoDVUs4n5hXhY2NVmfSm4hzcm2uSB680oOupkudmZdltkmbBwFPKgn8t
cQQWjTmkpde/y4bVI2UTDQYgLGlSjELql89RUHPz71Zm7O/ruYqD13vqE/91vXP73JZcLIKORu7N
IDltkQ0tUGyORoFK65mvs0W0lQczLeLzgattqxZ5ErPvlelUw11IokbpVSv89vSyC4sAJnv5V1zd
KdYlF4wstPAqiYH0oNsPz7GJe1d1PJhRUyKr4Iyh3uNfgm0qyl1ZfGbiGFjwARLcw9IihCjsxh/R
2ojiLq80qObDhD+zMshJNEkxgrPXqYBfVVIonVUiW0FDib+2vy3npJgchBQYFeFalP15oQIqwx3D
PAMHuGlgNEZzf7wSfBcoZI1c928eXOoaBmYY9sZqUB0ncroeU2pU+Uf0QnJgglHiLwg86jDWCKiu
qs42S1cOw1qrfxgOqG5sIfnP3dIuiMsWZ20eC1ICckLZ25+TgEzInfKFOK/okqkk1WUPmDT4frDF
hTlD7N+FGKK6DD0sfrPD0BMAJ126dDlrRXRZ+77rC3wvPDEnLeCRXobxrITkCecc8m1fXspWxjeU
LhKzFamdYPoBhf/dzzwKaoDAXtkUFYNr/0bnI4TNQ0qHRuTYAvRM7IP5Qb9/16xmcD6e97Lg/0SY
bgjEseGWnGj1dvn+mPlyBtMSLqnQJr6Esk5qDxjN/9In/mh/lUQ5HfSUc7IF33F19aQtC8YAGZD8
efC4ZqTEQNOTpe00tUSjSAGjS4L9J0dQE+5D0aTE4UtQ5g4lNOBSmsh8CLhjshOt3oT8b3JSZ+mU
glWXDWWYqBdHIDd38+OMQxNOwTD0C0FDkZ9/i0KLcWeadQ7nIVIM5ObksiJ38EAJu+2iqmWsUtgQ
Iheu05dDymWotS1lABflEH/eH8Di7hKojeuztxFss0YRAG4gqigp9WCVb++Wly9/VNidvfMoIqdQ
YEtJ3IcTYhOgiD+sQ6tcJKhQ8eTWgQpatNHwF7gtfKLuIYAWZVr3Cs3bioJtngRuwDiATrlwACso
NctNVBeVFvNSuWUnhvf/GOvZpYYre47a6jhS/OrNgn8mxafcOGc1uR7v2w8zNLm5q+nynd/oYxkc
K9KtAXQ6HxhO+MPyKOJv/+anNkMK6FYZ0v5JoV99eRCVdJ1myob1SAn2HF6GFHt+RIWeJ5Cfn+Ad
vCUNQ4Sz22riYof3tnpo1EHlcwP1/9MC+H9Alw2bbIfBxubpZ2uUDrHK5mlEcfLBs1Veq4LZmITk
jihzWPgfuAwO8f33t8lSoQ22fhbD7kwbopm9H98Ab8LLx8VCY8cM6tnVXbbk0MdjnXMz7Mqa6tjQ
zylX0sefP//FjcWNVQTWg9TBRFlXNZpdDJ9dOkt8eriGw/7H2GvggkYyaD1hr/5krYjAwmyxJF4B
/u9pAwzJ4QWvkZFi7J+GTX9JE7eyCYPxUEGDFh4HhtpexFqduLkOZBrJXXwVdqQBY6n1o/Icg7Yz
cDU0Koyg/taaemJ2ulox4uQp1oZAinAb/A177vFrWZn6VvhOIkXRJaDZQ4ghsBc1fLGFKPp9K+UN
velF3h09gQLVlwrLpHcj5bQIzYLMDuAacIHX+BOpRcfjJ0li8gjNLI0EuCAK/TuJzIxuSLU9n01d
DB1YUr6W6ruH45vOFIWXloX30yWUTCIk6q4SrFq2tuhF/TXtApmzVrKPhfP+7uT+Q+1xMdf+0Yn5
d3+2dFDQpyvKSmOEMqkXK3ByNOLWYwIy8+xIlt/RWzFsiPeti2EtLXVc8SnSXXiTl6438KXCQtIC
RkSAgDbTdrrbwFsFEmTiG43LWDsJAE2fPk0H5h8B71jtMDM/pwxu/MrZxjtIJFtuumxzmQTE5B94
sHJ7H1r/SeQIGqVIxOiRfl+rBzmt9iKGcdL3VFXR+zdyBljXLzUY7iSCPsXh0CmRzuUQGVL+0DPP
lkjDNcgtPeCBin/1p+4Bz/eZuka3DRtGY8Wv7cmBkDOhBGoihIxxcge7U2RPAAcZB+OAp1Ts4JLN
O6NXDyO7W6+TT8F/swFi0qrbLnDHeRxB17+KIOp8zQFEgOGuuVNFZb253jMJ8dUr3Z9g6fb/Qk9l
/xUXxfY7iXDC9ElRD1IQyxRXXO3yB2+TgNStj1tn9Yx0hc5TovXdsLwCjxvyApg/C2XZcTTXdY4A
+DRt1edsKT3AwTzqfyhB2JavPlZe+dUspQYuzXRTngOaCnG7mHw1HJT9i23oVUSZMDx8rHl+x3i3
OAEKvy73AmJ46plZOynNMu6cZmSrWdsWq0ifprFRusdiqu6OggMwAoo4FSV0crWp7afUyCnHObk6
mwCYqRJ6coU0Li9bY+olEfZV+mKVtFqSwfYwMXuZWPfvwMMzaXljSSulC+GKk5oN0wKJQ2CqznIF
DUooW66txXDLquGaujb+gASD06Cvuls2VQI/HHubA6Z4u14gzGv7RhBZSlNsojC3eetZQzP5EmHH
2QdXpYUEErKAwIxTlq6sUUwZN6sM8aagqSr2ltFTIJWylpsl7d2oGchryT5e1xlfbxwDhNGDeRmd
L5cNFW5rEnNNlGuloiEcMx80lQLcZFTwuLC9PaVfLt8Wz1KjzunRj+7qGssHjz96zjYmbtzhzAHR
hd5h2CNhfo+ZKWxN5BzwfpedTWf+3GtFwzsngpJzaBhN0KQNvzVn4APDslL/BtLbvhhpIRh7PDr/
5IAASpkoPuPlW7T0rV1iPhF+Wh0HC90uH13+BHRN92QT4ugSLgWrIAxNhVVKiVRVUBgo3xpooCWD
EIL9E7Qz8iYgJ2VVrwEplPVLJHO+NReEPyUxDtvzkzAJDpwvPm7DdP3VoV2rUz2xlHbpCI/Hz2xT
1qDMi/UQQ+RQtoyQIPDV00btX8z0ssOkrVNDBsOE3c8H4yu7Smu04oLE62d6Ps0m+Pbo3v7TuZAJ
E+skifUGnZzb/2oZ1BOdxhH9TJhKUXZcSR/Yl8WdHT6X9UrFHlqtIK4g813OolrWOoiS2ZH4HA02
GW0oFJ3eomF6NivzIM5s+ZvlDJd9DHhD2ALkbwpLmDrrxWyKOXGSN1HIARn4vNWvsJ9UXBVBnZuD
nrxj7tuX48NMkFMHuL7B6THZhllDg6j9qhLQYXWJ7JFCRb4tw37wYkP5OQ92x74BxM3qQ5A7f/6A
IvT/zHJD/EtteRCwISyGWDD4odj+5h2bQe9Pit8jCjS7MVlPL5RPw3z45MTDsvG4ZbS2Ybt8Gq17
SUChVS556Sf6l+T6Nc2Hu8O8k17oKQ2c5Q4C63J12slPqgFYEhbtcyKR4KXbGcTsz5ZCSbpy8Swf
4kWRd9u2NP+YZ5lh7/8hUOnbcbj2N1qI7Znv3LHUFzypQtJzFoB9hHQWd8SXqmdkzNkRiawoFJu9
4JOA/Qy22fkgZRFv9DVxYaydJtPzNcbRN23KGweu37nKYMCRMGGWQ+dw6Dm98samD1Zd92r9cF0a
Ig6WOIcQcJDoR2OCVNAJahkSywJeHN0aYTGuk+WRWN+sNqcCw7opA/SY4RoXxiYxIKy70lce7e45
Mku+dTZCvrZ5mesy9ZxHiQJxEDmCWFqvHmJcRM35d5SI/+QmxoPYF+Sm/Jeky7bWtJWdOjZ1UI7J
juG4PgMJvgcQ5WNBBLz/xBD3mDI4h/kRYcoOV4zHmZ7rDMkfI/Sy/vBJPintoMxuBBu5YXzVCrEb
vOmB6o/h7M6YPoJQNbnkUgZInCvjNRGQrO/jRmhexXwVQYGUZbMl954ThPqCWFYxRaCgoecn/gHh
WVVgXJTCtylmWLbGhJa6cFgC+giqDZoEMrUdfSe0BJpT4t3G5zWfvX24mE54FfV3v+HWVoalc00a
Z2mnsCmJciAwiiPlYvED9B+QbHjC3EjBx5FInUCxeVd5nk9u/WpG4lTGj+2Sa3PNGB0hQPmIwDAK
XjTypaMq4h45ATa0lLnlgcmHHAsrQyk2C0okYEImYgjlktFenETB2kyiaeLEzODlQXPYgocVR1gr
fxtCJvEfMGqJLg3xX1wHU9rC+l/XQtZwaEOwfN6QqoYHfaxoM/2IzbJCwQPEftHe6aEd+Piz8Ndh
XH40kcmVX7cizk4wuMnr7oSig7WYt+BVw5vD+RWX/AIBhpR8bw8/pnM8diG1wsPiC6mBM3SS9e3d
cxoQZWe90AwVVn5/dfcLsfwba0AgMtuhs2ufMfHd/n74fP63+VytrD8ab+mQup1eQfbk+S84Grne
U37RihVV8lbo42orNobU9GcSAt0GroGT9/1vw1PQmRKPP++466tKwsjnE/Gurv9PjEKKF7quYjDz
xalRNJBNINcpmlllXprs47evJm1EynkjT801Z4VK73a1NUPhGnQYvZveNpuA/YhBfqUDXOK65Nn+
AlfQ/nr4ZjqJVRuVLfyllpJt2z0VqFQzc2IB14i46pPLf7oD6E0WUFPyaUmK1bOiC/xlCQUHphSI
e4dx+b9gj/LI84WjZ06x7o/mfLaui2r3OaQJsJ6m2xdiSe58OK1JTUek59DvxjMCuc2NiY/4Y7/T
/PAexLRDUU0C0tMQj978YdDh9zqzfROCWN2lOc58hAPkZ4zppTEvNbo+QEegcCxguhWpuwxqEmfO
VgEQ1i9KOI70Zl/PLEueuGymvgq6QgtOEZJrgZ+bqswEHgSj/yFlXbi0kqv9NBfw0tTh+j8VuJdT
0PYMVW2K8pxbixhagWelArfymyxgSRiXDBdtdcskNnsjeGykmg+IsTPgQJu9O5Iv/F9iXhSvxCM5
dxMHGb5aBv0D49o82ZjofheQrE9OLnD0wqmxdx+Vm0czP1GmOhv5bdBwHsXymzA8nLdQ7mXh7fC8
gMo70RShBoa+cDbK/r/d4FLRyAg/62ckToXjdCmkmjzwIhgGi7JZAlDXBsmllboqONa+nYbSCv1+
CQqBl0ZxXa87Z13KPRAdfOe1Kw1zmfYkKLkt42zR5DyRj/I2qOiOb4zmKGiY8tVgIsmH+InN9hoF
pDTuBbpMezqa8Mr6T4knDZVmgfpH2ZPgvQAYq/OxsKitxEOxuI9d/i55UtIyd6dCfSTJgTmGuNoV
bOwjbYskmv059Fhd5WlYTXkA66byEQpYtB9UWVrJTO+IxKUjnRP4o+h68nTpNracStV8ZWIEQ6F/
GZgNMFR46XnWaLb0yTogEH/ECxCO94aMxicI8smx/sSpULx1tIgkr60gWtrcvtj7HwU3TzqPexc4
W91cLMQ6Ho4qdfUwwrKHrhLYS7KQJgU71S5DFuAL0maY0sA7TtFDSMndLUCpiIMjJgU3mse+W+B2
kXIB37TQBpLGPX9ZFpCKS5NV9QpF8Y/+1eQJVYgQa0siem4D6X7oS3GBSt359eBgflxeJAj+6hF8
YAJ+PxfbWXahFRuMPKzRsYf8B8ZpNx4QixVLZpNTXtssNUIw2yWB+NE3W4sQfj5fcQQyceuGEVik
yuDNANPiVN3zLFs1uYZvIUeVfDVj/c+j2OUxC+k54SJVcVtVzyv9Y2xv6hqIXyIgkO3eYcAm6Xdc
/WTIBQI2s4ZFWWpeDfqYbpDrGWgG/fUmvfZ+1pYqcBml2LOCN3qz7elT6ej08e5HeQN8fOXZC7jQ
qtMoqD3RRSeIGyEvnm+GLno7mQMDFsDL/c70LP1prKkJzpC2UI2NQ1WiIx7IS1tCYWGGERdr3Bfy
kp7xS6vUHlY5nIz5Qd0fD9BVqTC32QfZReWjByaZFb5hTRtsH0zPk4NIEXSNxvQWpsPj3DaP4DaI
m998kUyl6eFDIUYEHUQ4egwlteOz/lx3zpbO7Ntw0YyG5zo5em4t4c6afmQfy3GZfp3+WrnjF4f8
LCULwLlf2eIRI80SVj1fblX+zQ2JebRqbTnkdEsYEQtg8fezxuBtvHb5PONmEfF4zOYMJBwRaHGA
ab5TY910uffTXfd44RwgZk7FFTcr3QgakvqHl/Reg1TZ70fdd/QWPSL+/aDihTxti3f6McGvYffL
j5wHgG7pyAgKiWIgyVDC1fthL9XAEzGDc6nyzwCKtFFYvGjqerYCAZDbNhYEi1Hi/CZuYe3+A2xG
0ISKZHiOmbExxEhFtMilDaQvE9IDw1sGsjPfe7S4m/pX/9Em5GfaJc0+23hCrye+FgxSPlRmifGv
0J6kipQuQuPdQI7EWwxZXtW5i8KTd0X/fv5s7Uk8YCE9D2BwKvU2qlu43FsvXmoyCeXm3p5uDmOc
/f/t6J+Yicxl3K6BmN0qPq3YtAKHQnsYBW+8L0vE4cE7pRb8K8zqiCrP20w+4GVD/AoNZqz1vUGd
f6UmEAjzyLOHOXlB1LJnVtz9a4HvcmK5O1WGe70139ikT2KMC/AOLZboV9vmK+KMS6j4KVeXogCT
TPNJuDmyKqR7dmGwnI3YDUeTdYEPB+E63hR112OJEd8dvI8pfc+PfDb8Qxz7yCfUOwDXkIenkBcW
4krZ/77ZzqRy7go+3tH63m6tjLaN587EIVrgXriZW6NbZ0sedXPbvlT//X8I7mh4KC7kX+fYQvz9
rhjyGXks+wkAogXP6uAshdCx1yTl/PMappG/aXdxxJwjng9ex26UMhhyqehr/BHeYbcO0HDEADi3
QhOiu7ahlBTdadj+gpPFG0LdXSS2/dU+/wePUuOYxwgP8ADm2nYacHGtqbb66dT7p7Oi/1pqpqb1
2sD04RNhuW5YDADdvD4uaR07vQhBHlUHr71Sfa0AVIOhCZVcKk6V2MTj4c3LhIGKUyQ995nBhXOt
S4U5VUEFl+BXxCif3YMQJdKnW0+kEg37Yiqj1k5Jti0ej+/oslkHzRYaZ2D2HWGipDz0GWGfdECJ
vA2Q4+mSn4FtfcDcJAqbWBUAJ/j0W4fNpz7oNQxEsLHkMN53K13s/okgcSoPSFNwJwH2GQZ/pu38
nIFgnR+Y/Lgat6kFZ5aroA5ReG3EEWjhC15YQesg73K16wtCqxOrIp01K08b6PqEv/DauYFB7FDj
kmWp0gOeM1ceS5ptDqlHCE4Zagp9leXmBmj27MJLmubDFSRhflI8G0/Gb73fktukqVuj5m5bJZX7
27HDCqA7cHvl1niP3LOTbhwFAm/iYSYguYXAGraWnuk8dCCT9JRYecBHKrPnhPmtjsRHX7BsQ9gm
NYyBY30GmFthwYqx4lqJ1IcCPfpvwHXd0dxnvSGXHiloOG6khqj9/iC3vlFlnb6AwRQj30rMm+dP
QQavW39c0NQFsj5QVnyMQIcOiOakn1VrH9InyX6naBaT6+yb5H9Rd51psx6Jnuc/P7E1MwPtf6oS
7U1q4cQVaRmS0wvln4aL8s4LheKSd42ZgyboPS1j3mAMtauY8IDajvQHOO2icwLDYvT6a6jrNSGV
p7ANn7rNwM01cGgnuA3Hh+/z+jJpEfzxraBJOoZcqu2gNXwbJnvikGndOP6Omt1cHdLtpi0MTdt2
p1uhjBw7YulSH9L9joW5buPh6yeN8OGrlmFNcBEX4myMGTM2Tp9IJgvjOKs+jEy6Ef4IobDe6cON
R1DW0iEqEelkWv4/LXXYLJKmjlMwiRZxThkF3zZFJ/vMj4ZbE2FU0nXq8QtkFu6IO/EBRRhWLV7P
24NmkeGGgLVyWpPiERJ2Ivp4irFDIGllEb359sADU+haoiR9cxewIYtBJPXLaFS9qQ8s7KzduCGP
+L2mkpmjLfsKKIzzgf8DZVzUzji6ZUFP71TiLRg7+OJRT7duw5ZIvmVMGZnXA/+1rJ2ZSF69Lqdq
bqYnDOKPGv8JB2xXKqNpEsvojGZAW5gFikbq0qC0LZgh0q86cUqlUeRl62h+7xDPRas/a9hFKfu7
UoDpNKuRQ24JDNDOA7+RDyN8O9cBULqOnyQXbvnIPTr9PvndmtyzI9AgsrtR9RdZ4sPjgjjpTPX0
YMFAXsUwqp0YerAEySZUe1MikHW5vUIAA2190Su1hds20o/teK+XaUcfzrG7TmQP26KOtnkGgUfk
ShT7l8n97YZWp3w0n8lp/GtO3Ncj08f/Gs6q6FLdOCvLUksObin7IgjAK2ZLOugBNbR3vFbeHCYI
ZGDG2GHNjNuDeBLIg2Z91lwNTh8DptehF+T/J5jXU3+Y2443N7WQWaqkDH//4mGsrqIgwu8nP8wA
iA25hVEOyRFEBeJwRyYlzLnDQoiGifJtwyqnKdnx7iJgfYwJDWS7RMXbIrvQGxhkSeBLYtV7uIxV
TP9Tqzs7rLrxXhGStfNKWJgduqbx7U/MGcMgX6LbIu56XEswB1SLJwQokOMNHmf3T3hHVrku5hdP
zDlDK1FkFYWZZSYAiSAiwiryZcvQsmGmRYVPwlURWUD72DZbPTJxlStyG9rhLhq6P3eLK4k8gyOl
9fGjLbgLpOPvGGYnOD5ZfjjSwqCMeGHglnVgtt6TmcI5g1J+G13C/UonpPOYYxcyvlFldiwo4CMw
i0hV80E/MqSW8MTepc+CMR+ixZtMFXyPW9Yl2pRoXupDGqTiLfCL4+rVjXqpqZwM4euXlpQoFgfs
RI1V9lzhyjfKO9W4p7bErgayoWd0/nwsW59JJJw5LDve8ARf5Z9Cb1Qf/BPH9YlEUf2R54PzNw9a
ITA5tt96lBI0LwgHAt3ATe5ZhFcYmMqiJK+HjOBclAle+sGDknvass6MzcmbFDeuo+uBLEm7Qs4K
IpK/E17Ib4xpWf/9uUJGCyuSYum2p6sYree98HopBuOj1JCld8p2azpGrFC9rrNWppdOAspFdzss
3DBKB572dEzDvEG4rleESljdiRI3/pZFg+Um/NIH54lyrTkAy4cxqyxtEejWlRRwP0A9R90ygEn2
y9CUFqkWIgu9sQ+CQx6jzkUoweZDDn+q8pRNdkxjP+wcZE7J/NR+Pd+h8oMSmko+wbe+DTLDr9lE
zFFjCd0hXXDtS94kgDWlTsvnWdLEFp3ljLEf2jKh5Va/t8a6CURJOeUBlcSeToZdEuyX55Nw3H6i
7lD86uIcQQvnxriGYyez1C84v0HjWQGAmfUvrdI4c39YW+HpRkL8uOV4PGQC4gm6zQoc4IaHj7x1
F2G2r3weJnlwS+QBG3aJdrF3SIXOQzYqbQMUp3XDMPFxGdS+jcaXr8hhBS1zKMl8Gvxp3/jaCyBF
lPEWWb3yIuy9Q2KxPfAMmkFnA35xPcHLb/WsUaAz2jXDW7rSXZqE7jweFH0S9R64+BsUnQ7OwkJM
Zd73o57Q8ctAf2DDUtfaSxgwDe1VqYLlJ+y5oi6A3Cys40ZsFICK3XTZRgUgDtfdM5HRgPt8yvkG
q9hp5hdgDEzyYBtwkTlLZjsWfQCFRNDUh3ncGEAa4Fxt4tGtvpZbkyOCueIfvikKw+R5oiIlKZ22
JcD8BVbs+kk8Q6Qyn7QNrBaUCq3Z8350TyjRcVfAh2AiIHskoWWuVvLMNE/CpIItdrqnS+lMPd/x
qN9HhdxmIdoxMIxv8RwUInd33o7qsD8C+msNe2ywa7hFiL9JNRSbQkZ6hUDw33niEso5D+pWPktK
81ZiFGJq00Jse2jeOCAqITd7lRsrb5Ms0BlKhMLUUE4EW/KeyEiPHj7S9cxJoCsRm0f3U0+J3gsb
JpMoPNsZrJ5uyfbnbWS1xwTB/HmQAEzfqGFSVlcEL+q1+2W+F4iN21NM/Jdlhs0BWwBKDgIPeTXa
0v2+h5WeeUVKszduA65ZN4fW1+xqtEH2DRV+ttBQF+2OPSyM4Lza/H1M+y4Wex8tadmqXPbQyFkM
Y8mR6xePXCVrLYDDyIXcUz4JyYtvOS8qv6TPlh/sO+VRGdo9PE30Bsg7TW7PfuS/1JhMU4TlW2cQ
h4xmzgma8OaSOuJBt3TQD3A7w0hndAHuR3q742u9scMUBUpPYyvoCD0wdeALZoSibtYOprBRT40h
Z6d3ktYzPa15qwxnLRLWnuFhUKmB0HrB341xMsFkVjgj7oBUpxO5PFrARIRqJPk0RJpbmLphnzl8
iMLfK14uxAVgokmnmybanRCF54/SwQTZH2mPLUyHukDKrSsKxoPkT85gvlGn2xMMFVP13XMHlNTO
BWUqdrPqXWqVn5ByzILBazV5o8+dl3YTndn6KjNKStbuS49vFmMMq4QLAystDuDEvW9QwLF3zLq5
nKH0bcmxFl5djzB27OIpIpe+E/2SDwb/zXXpvHJ0vkkXDOgfoPFNxr+w0hw0FPl31uyNm4mVNYAK
mb3APysHO0KMWa5egwOycsFw08H8SiJ6M4C+xtrYymohaSjsaIUHivH/vX9xjoPJI8ThcJKxfAAz
2HIzgtuLRx4ptEZBXjOOsMrSedHBmBut0/YUG8/+YtPeledEyERtqOlD2oRw/5feVKy/0POJujLV
B1/2zqb42MzhfD2bxm5ELXA7mzVklmNMMQ+XIXwcKco6rqIPENGW1lqKFgyvgZBkZMOn/gJArHqR
KryDQfWRRimptOwwgNdNjutJq40EW1z7g7U5Wj1WxlKPnoo0TMZ/5p20qUSmhGlISLHw5jGLNLhJ
7JUaeu379CVYlTxPZbaWBH6rcRdSs8VhoMzbDueRVzTDTCSS7I1ImurWJWO8MwGbv+QdjNt+W3Rs
CAxiGwYXS6j9vdpvQq4DD/bO1DNIwQJ+7Uk+9M4HaNZw8wI765BuzQF69NW+Voj1SIsHNC/J1+Zk
jid8r6lh1g/cQPTrICBOYzD2rIrKpkjipupwRKovRejWeNsC122mq/eggJFs8VORWcVm3I1fdaQ9
/IBkgxQieHhhVXDomY5H7JCUdVe5tLhUDHVur+U9qpWkS2wFrAJi8JLL44ppGHb1Nrv2bhBWJXwK
PNaMxo7wyHvP77lpkvLQYkmeSsAq7XY/1sSTI+TtppRlwAQWQMIeJPAScUSnKzvJF7NXSniw3wlz
6buXwojRPejsOnfdpvLNLZ10oSq6LT6Dv0knPKsXmU6pGlRii11fyT0RA9jCLQk9xd02nodq5d0P
+KlxoIrdHoFIp4jT+uV5DrOhe/3Rk5h6d8l4trB+3arTjXjzMrU0qXJb9i1mqX0l8J/xTgNi0tWt
qScioe2F7KzhTQaHRmQQZR+OuA9C7LTyjGZ7QTnblDp8v7vwW8iXCzXVr/2v29dX44d6CSridc3k
5nKs7Kzp/riFeN/OJY7T+ufbGQKqnUugToH4SdejpYIVpfNkDSiQ2kXecVuz3YxZ/CwmrjI6EVh1
FfjXH5Z6Hk4BZnKagOUPvZ8ayLFwRmEPkRr7QDoYd0mZisUN8f/iY9EZc7NWrrKZp0Cs4ZzxtbZh
d4dbufCexOGC/1yX0+/8vhGq0sKBqHfh1T8WAtFLXwMlT0yLPphiwGqR3gWALW4sCCoyDDBaf3pW
nPTG1nPukFYXctXWQYQDE6geb9YKyb/pb3WD2lXmp2uoEW+w2HfiuUentFdLWr7ftH4PWbarUZ/4
+AiUT5TPeAp6Welxb6Rpx8Vz+5J8jYaHtDuZncJ3UatrvdB6aE5mx4gNlhrOtCQLuB0odAo/mSLk
yoIafeN2JN9knM/8OY4dyn5iB0lDdtDnZlhlzzNKa6kAaT2hfO6t+WzzHUi84ftX1gXx/J0bo+V0
Od8TQuePzgx6RVa++qOmxw1J4+RRn4vI2LHcj99V7JHmhOYhx4g+c6/zTSq06I0/PrqGlG4jogfF
EwYecl/pVH5wTdjElGdG+3qKY02j4jtUxp9pPnuJHHSteC37Oex8ZD/oUPMFRnp52A1Zod0WVuyU
9ZSfyn4pw2FMSUVesvrzcOC9fM9P/XDbNt/C4HfAaXRq3weOV1R6NQ0BYf+Vdm3mFWMuUGCz6QHK
bWX/5PdLrZOZMnv0GtwWLBtWOZThYB4kZcHYGXqBkIkeGVgwBcQv2KLUVURFN4WA39+ucVlQpnoU
wBLbCR5d8ElCrLdz5iy+8kTxYfyrVz6eaT21omh9Lhy5ieE1Zbvbi7KPU0/g4HYQL84Hlg+G8HXF
dCWRy5rjzCxogNTVQNNWOP3c1MydRXe2th64Mmk5oIjaJvrR5c9+WNfKXr4B8fDfvqRDjOrl0+Od
GujDQ7PXAx13w2L64nPpwyc5eD2K3M2iJ+eATQh0BThHYM7/S1R0eIuSU2J9BXs4d39AgHmULHWl
nNt/35bUGrzDMXsafpJkhhXX2YHB+7uNgOd3xIC7qnR1bFRyNXr6jt5x0j6y0yfk7UspBWqTNOhn
MJda944b46rT98b/0uYEdgVbdyi9ru1ZBFqipVUH5sXjLSrsFOfiin0wR+a7mu4lRHf0CMtaXeV4
rFwan+5cPd8SdXGR2EVBf/cyHbKUWIlnlbSVwZ12XcoOP6T9pB+2QxD4Pk0/wi+vW700pKTrzbdm
V6mp2rQ7sYEBqB4yv3CxYiDtjzvkqf5mi8WqUNdujFTRRHJaf7raPTTAa7bJjTL6f08KoGGH9bQR
p+o/gvcj2BtKGWBC075gKpwleL9Mk7AQjsxFodNx/0fn3IC8EXZFE+Sr/1KotaaTVa8PFh69d/a3
iOXIue+JkcPegBL4I1laMJpswj4dLptCKeS2i3c1WvR+gyia8HraTXRFrAQ7EJT55kNhThKoySz2
pp2FI9K7ly0xgk6PbgEzJUVD8XuPW+U6bj8qQvMRWi+Lq5hguGfOgUKU9X8+vjUJs/8jh+6Nitfs
dgLXf7EF9qEtSb3yc2ugUR6N6lD2z4eLl4dbVdAMH9UVsLE1D0Q2usMPUiWTIofsx1V1jQ3SprbI
Zjt/9h5YO8oY7NzfaNhS573FjmZ+W81qM1fYMrWWXJZeWmj0JwD8mUmWPrl3CN6ZLIhZriYbLVKm
MqKID/gVlWL1YsswcTMS2W2NG6lkTVARHkhuSwRJhZufouZZCPXqXKj8dCJNb6HyqK+aM1uHZCI4
KhYTD8WYJHEWon0+Car+f1sCrPXh3XN4SXV234ubv5huYyXmjBsO2cBF6xyp3dTY2/h0xKwQ2TU1
ZQtqeS2d54+kvlI1NJJK0Lk14VhcQFHpBPrqn+Sl45+NnXLctnqa8u/wSPPXWovw70EgS7n77UJe
tbjcb8fgBBRfjACWycCGQRlhs9g5r4FkfdeQLCudwOADKt9kv5IgqFQm3DxhGYfOP5J0ec08UTSf
lBti+Pu8OfWbFj5uOC4VWEFH1ddIET/cumxMXRLE9b99qswsAesDddy8Di4QcgQez5P/zTk+RXfZ
kg0sFr/mhtBqBVc0NEGiYjpYsIHWBzEzm3V1bZbTH9Vcp+siz5ATYASF9VTPOJTTyPiVyinFTIIu
fEojAPHqqRngLiSE61td7fGIiinDPDWjpbozsrPBbU8XGXZoGJriV6rjGttekw1IOmOyTi8EH5qx
BpavP45r91mf80/67CovzVzY8yF/KIEkg8vucOGCQcg5nX2J24e4PVwVWQUbGjKpRjJDD3OKw4Sx
HaV5tFIgRfgcG3AQpLg/Tael2TR/LLnoKXGr755g6KrkU1nQqVBq0tsWIXVqYMCe3WQhHwbxuzuo
MtT+VCnkHZZjqJmSPesvK8sq/MVvdrGGKMWu8T8DKes9D/RwMb+qLzw/6Mf2glD2hpOabmKrHnPQ
43y2JOt5CWfMgebkEOq5yf4RwcAXFk3Qvk75UVtUNZHMl/cFu+qCllyR1NlD1XOe2EnEPBcLi6E5
DCMW3av4rL3baRohIZ93jMuqxCclLe8fP5H7VS/IpuCj7eGC8gpqt6vi4sfBLDAwD7BxUlWeigPa
BJkhXzWTzIkP+8mHNOYKEDLoeCeKUSgoB7UZwFbU2gxHphCf9+m0Qwu0TOsMTTrF6N6V3IYcPlBX
2ft5kxGLiCA6qifjqYc/fTpdfyPXzu+to48bZG4+dQSJN3bu+bVWy0VN2H9vdpmaypZ8FzYeJAzK
pOp7nIbBCmDvD5ZPfjEAkOKDCM7m48BpRx2MdAs4zd9XjLPgUjOJS4d2wf5mxCFK/NDnR6h1Qstg
y1R/PJIjUV8sVqopQbXWP0ZzaS1FJHyicOXZ3fPSTtuNrk0ITd3iGJa+gCxxv3Mob15jFtvYNuK7
8bYRJDGd5mEPweu//QjDDs3hnLRMxXRgYWudRXyBw5q0amIWvPoK98kieAsoiBaPg8/5nwXdzLRd
8XIf5GLB/X7pXIYVAMjewW4sonVSiN/j0styHzHO5LP6DAsmJjmvux1ZizW8LGqQ3hCRu5WLfldg
t/+kK8E3x+Asr2Ikx25poVVi13ECk7/IJJoIJbkGi7TVygsPDf+FNvXS1cm2uW8if1JiblJyCdDA
H7ikP9UT9ir+FGZTsSotIC2OvTRisrBE93pmTUcExxsmhA34tx3OzVGVeOHmXM/3ZyeF3RTGo0kH
30ntqbhSuKxPUOLkXOY6IyPOFWNIp4B9perCKBSZ5XvkCVKFSut+iNBv6s1k4XeF6RPULENqpxEG
Shlu7KV8uSZTlxD1iNyg5Zv9H2bnWBsD/Gt3/pQbHYyyAmQvH5GYIOR4Xzqmr23Zq2N252+JaQsy
dLDlCbOyZJHPOJKboCcoAkvSOi6NfvSYnWrUOjyxKKHWjsKXxQv0Uqc/OcnRcrWg6djFZgyPfwal
VtBNqiaMnPASTluG67bb/gHFQ63ZzPaAwLxKKbR+xntwgBMIEoOBwsKZ3zoZr6Hqn8Ut0BscvuLb
uxLix4VqaLEPA2IRMvx6m9faDKjcA5V4oZ4J5ogCrKxbshZ5abyL7V1wo9iGgakzwl79Udg8P3Z2
QIrG3OZkNS32wSd21OKjKahs88dzVZtxbBZNqBJMQxuFCoijpQ2exteFzgYOTon2sSCtWsOiOAhk
mOcvTa7Q2X9ht8lMp1Wukco7jQ+FzWXxInriUwFmVGLosM3TiKYEH7FuloEsfiBr6aZ0WPc6DDOW
8j7OgcLpivZGIKWriJgq8PpMriB0vJe+qUC5WFosE6ixKVkkJO0a/RFWhCJ4497UNj8i/0lgNudc
MrY8b4evLvLfzkWhpJ5bakz6bRAl2Ue9/d8FJas3TRjz9TakIP2/jgCoZiBnVpXq0gsh4Cc4mPvx
7ph93xD4xI4dmmzOncdbCiJ7US2R1TcelsMijJKybFddRNhceM/MsILTMI2nj18OyIyZTl0ChjB7
Qa/nortiUX/Tn0D8KakUci0eDRBvp+CFv8NgF5pGR3issSi9dUb2QanVPhito1lX7PAjgzxw7fgf
6H8eecX+uVu1QKmgrgOeQX3NHSSWLiqzuwkqwdrnXgT5dOBEfQD8Cn5+Nv+Y4jFoU8CZqQDCBt43
JnZTT15yMpzbScRwjw6/yZwaAVZO/pegTdSE1synImxKCWfXi7YPT1bLVf2V66rt++Bc2G9HlovM
mzTSGOiq6uYKheN3TxnrEvovJzVLVTzMrwuagpQXR/pi6EUMQ2iaJaDG2OJYDIAI5kHk5wp51360
ApomPep6PYIfZQGvU5f1ZKEkcjQxTqig33FXb3I4g/1KEXlXG7jwpQOj0kit5RLctBU6IHvMsdQz
rmOgk+CgvT0752yq1fFQfeXGpRtUkuTr/ab1WH/uvM28aYJIhJZS9yE8V2JobqgbEw1wO2IoHAI2
Vw7OddtYaHDkM6QJhb9MF8uLQNV4tp0i1Ngudpt2WVXCJJTsWx4NB3R5IeXYCwXaO9hWumRwICOp
d6IUOvdrxIer+/+/2g7/auYv+PiXBLj31GKknbeO3WtexF42608K6ikauXgP8Szfm0AC01wqyS07
Rpb1KsGdKqHKqGtRhv3W2Vbx8geKebWR5cACucdIWwQ4cpHGIbeFJU+ttQ/s0SKAyigTWTBlWkFu
bcaZmblYnSAqvxcLDgeRfVg/JOhteDzBVJPANPts/J37sscTRcR6/MAO64arOuA+EzLBIBJ46XQw
bJac9hnIpLWm/q2LyFSMrcblGpoyGEFZFDQzzrNnGZawz4XsU4f8nfZfjfSqU83G8SEB9WSX6Tn6
GPKqAz70TxL0IIFXzrz4R2nabyv0twN2cXwPiB/fzHuhiIyJ59jRdcWjBCk4u0ncPLFuUR332yLN
5HE+ZJSNbw4ba/cssBks97Q5gTRoJ+sgZr0wbgSfzZQRTkWWQAN8QXdlgTm9qBojVBRZVmfLxGnJ
TzZGFe5oWP8knER+WYG9Vwa2q47FB19aqOxdwfXjtlSZ9FwhIzNccdwk1g9cHdtwvbvbV9ZFoQRt
uhNtn+vhj9YurjswW8/G1i1+MhorlI9r25WhXFx13u4n1eGhpsZPwzOXhnmKtkaNIROqRFkzXjyi
V5TnQKTlC9fvGxC10ujMcuEg98iD5J1RmwdFT3302TQ3bzSsy7n9TGklz4lv1UdZyFUwwpXPzG7g
YpR/jzAxdSoejIlXSgxGXdKS8+dulkZ8b1n92lWPl9x9N7wOIwrzNjLVe2h6KGbGqihOAkeMs0Ws
U9qp479cXqWZCRVel+hPJxEgCB8BvOcbHY/UZsYq/t2eXPuOnd2GNOYo1tz89CWCLxb9PaOfISQK
uQK48buoccVdYzYb1NKj+nQF4EjcX5OhABXvkLZD8XOSkIFhHo2a8/lV29Imbhu4OBGKl7lFrPeo
vAfhgNsEYSav9qA1QO3kS4QhhL7hYC7Wnso5u3uvjBPBeJ/LZXnix6ntN6Rg1ymNvHP22hoxvbYu
i8Bi+zCqmB7Yld4oMoElxaJyJKu2zrEYqmHLy2eFvMOvmfLnfj5fFHKA8cbSokxSAwq9tobcA4Dx
Mf/KEuJPCh7TwjqwmCvb9TG4X2jspNZwpsYjzq8R7aeeHwNkK7t0+DTLQdDjMRGBtMgnLIVDA5LH
+itllxYyJnINzasGE+6y10Gf4MtawWLCk1of6OPqGfslH9ZwaHJb152Iy8W0YQvZAzW85jBkN7KP
YsBjNhDH8pJFtquemv8L7uINKS350ssKKo0dFEv2Ye66Ew/NYvC5C5uBlyQmmr0OfCKg4LmvXZzz
LakHAYONk6PfSG/VSEEaZNXXTVOTkMrqS3yskjy1yB6aWpdpYWkcb+Fah9oWazdnsn16geYzmuDi
5fyXjYQQv0Qn42UNrZfK8Ph0n8nHfOEkbuMssK11uJTKjbRA8l207ZB43ShTQMv8wPd2aKqL1hJG
d8eh3FdE7ROrCrikolbjRzWt60z47Uau5x1N+add7eIg7YVWfwkgXg2heTHAIQXdUrgNS6J3ZsaT
EJnjMAA5Sp7ickvu88SSrs1reznZ7ekWE9L8xYHYwn62LNcfIJgvf3mnALlji18P0XSwA24ElWJc
LQbz52wUUDmuhGTP9XYC3JlupRybx6dg6yVUcQfHqbQxkt9rwMVCNJV/fP5qGtIRec5Cq0yIiJQm
C+mGEFa7w2fkkoMtqw0h3p3bVF9TVgVlbzYvu7RugDTSeLY4OTgKJS+V/omeIEg28n60G+2TtPwa
k1xN0jEndW9YMDLKA6I6laMRNItgTELsYoh4ye0rNp3aOkpqHN2CzVKbvLbyDMj0FtNaMsK052AT
o5hru9ZgSv6NBTe36u7k4dVTM6MJL7IibopN9pZsq8b6g27OO0pLnwV4LjvhQXJeyv6hgM58KID2
KMyUzBoS8sQZynn3Ogd9GJVcPsAPbKHgJ2cqcX7alfJ9cXF06Pv4JBJENNFmaxcmygvEJMsd2tL7
FfMZ2aKnNkYQ9ZlyqSdgxURy1nGsNaOa9Kcyc5ToTey/M9+gsdOxOISlCuN6zKCPFN1SomZsPrHR
au/rdFM8EKLzYA8A7zN1qlKjNYQX/WxSiHKVaopSnwTsf5GB/tKyDOQ8uH3gjDLqFN/d/j767DZc
uBjpIkgZR24DinPT6IJH181msJCK97fGxvSUJB7DEWi3GoyNWj/jfFFazBJelbtUyBZmLOAe4kVI
6RxpJEYklUxeuTgmQuHPTvbebkg/pn4GUAUBFzQN+zsu3HOt8UJALtHVIrm38LGKCq1Wms08sHIW
IUvPV2slVK4AKX5QGgeg1thHkO3XuxNu5GcjfjB7VprgBmkXpJq5VwecRzQqvIHux9D0Gw62iaFa
7xVKqtY/Naz68QXbs85Rjek21VFFVzpRw5eZT4qrqrTa0lGbzk11y0YSqzPoMeFaHt9Z9KgMHwre
Rag4QMHYVReM73gG5Q3YLNnlC4QDyZHvCBcK+gKIeJfEHhJVztN+37WrwbZre3Wp/Rtm3nEjQ9y/
+Xz5zQzKxsVFu/TP0iFhpZ7r7Zf7aGEI2rY/hvkXjC4VW2CNUj2tpzK5E/L9gFohMK9yhmMDTboV
jJmV3KNzJl9fruIMjX3lh3zNC73dzWVbWc41o826DXmRZzhp6K/VwKVhEPKefDgLe9cc23RmZjJx
6o9k74604qX99TxnPPtxsRxiknSYrcUZ1OISIhYstnrhD2kHUzehYdjxqdLnVY+OloSsXv9GKwbg
IGA6vJ3218sGm63p9nX4tyazCZBZfVT1bDNhomy3otjoVjiQEQ3OPJQzA6yD1FT0qS6LSoTXzgts
AdWGbg41PN6KNvw+v99GxJas0C74yyvFx6SJKEoJwcmRAgH77FRM82qWwRdPGfev5Uei+T/7pOYL
RbaVFZETmxM9YiQg9uxOqztQCsk6TqE+DP9f+msuoXMvpdyeAQlHOFjq0ax7Mdz0Y9sF9L4Qhq37
0oWeK3Kf7ft5pWJ36lDhx+48AkL5nAxFMemJ2UMvnHErBgCx6DlMRbgSPfdnbgVZhbhw2IGruRxo
3XYOhHiHh+q74Hp8jGOdy9EAHL9OmiqDrbZhV9bdGd3PY6Rw3hKpPZviSL4Y6x+Nq8INLf+EeJd9
fvMQ6tdHtmdBEr8f3z0NFebdGbfLqva+0Nr46LRFRa+Gh8o5ceIU0QbmTmC6QW4h2J5y/Oi5jzq/
zcVgw1Hu27PeRW9J47mUUy3BdeIK8MqIMnbcuQQOr+1P14l6f22pGQSjIth4+KaO+KbtGbwGm29Q
3uXRmb6dnJW5uaSiHIVVfh3Q7ESK7ChLS3pq/vrbP5yI9L1X4y7LCh+txZ+fmZ2nxc/soYVmyok3
l3oBLSzVY1UzlZgkNum4mWhty8uGDr7X4I2BY8sWcmF53Sjsx30GQNfpzBEYoxgUeJ82pE7gawt+
KlD2MSJo028dkKTbWsMRkIPgi43kutDGYEhn/zjeJNODK82DmbVgM5uc0oW8GOMOephcepMqOf+a
iPfXxuhSoAU251ZLdnOuJU8kwUuN1BwGNbWZkU/GZ5uMEl3gT+C7FCE7bUjArR8OYewR16i6qVde
SMHPIDU0CWoDx0coCrU4DtEYdkGBzO//ZNma1G1wOA/yE7KrskPodVR/3t/Dr7puYFXsv1696CVw
9p5AlnEEgjrfungohzWmebyomF7EfKwl3B80Vdcv0KhJ90HGd0tvvCwmNaVsYGAtV8kwP79TpZ31
MOXfsijyVkMj1ZjurS4Evl6gEyN5ZU0g9Vi+7erFn3GKWx0AFezTslB2imkseKjm/+/cWpLfkxPe
sm5Gqrq1PDyYjoQTwuUxsCpJ9nCXte8oI/zPn9t6UuOq932uB6s7LmZzjm/prKv0cap2ylWT4IHT
wrYsu3OTp+os0olk5otc7fBOVKwp4IW4D8hxSfE2OjIgsI7pONUe6dnsBOQE71l1SHyTz+itJaQx
VC4TJioPOZZtua/zt+2l7SaxadR/lF9jjmQRx3eQGJZM8MZ6mrNYyxWiSOpRZyPbbwmgaO9DgI6u
JQjXAlrdIGgRzr29gOZqgl8Avogm+p6I1rFF2ddrGCr13pLkKWw7efmZwNZ4AWxKEDbpMweHZ88C
lMX6J5heeroB7iHohfXNv1/L2aI0rHt9Iya5F268hNLMew5WT6E2jfLM7Ngaoqdap9pOrI+0Ext7
3AwG0ol1Fkt4ex0eTiiUOZxeiE3WDT6dxv6H6yYteHTYY61VKVv0l8+arK64+diTzQ5pKWLAs+Qq
6jt1H09wXwQBlmrzQnajsZMdJcOT/W/ZJ/0pD+QO3dc8axHWaG9iwHLLHj/KQ4mvyObjoAyFSCYa
Tc2qoETg4ip/xSQwuyKyxtfjzvb3nMeeL4vv75Tcp1nExEx8i3CZAD7+8n3nOE4OktR+kBMforvQ
QcCcO4rcbgIaqXcJ8P0SVmPd6KeQqMuBOFBzxSWZzYqXlIIOy+vpDEe9F30qPTmGDAjiSN3I94UE
/EuG2sEplgZe+LKTjp772+QSzNCA9n0EKmtK9V+/EDHr0SFzb9mzy2tuo+iLpC5mDYnbH7MgraWO
pQt/vD1h5QTZSdxMhIG5+WwkYmeCTPpfQdL7MTdhVPfL6UODVNmec/ir1f0xk+zaWdo/IhPhYEB9
aybPFViKNfET67bzXf6vMeiTNZRZi7Y6Gwjcv2TBNTP0qT5Cb5NeQcUc4Cx/Pwc2SFCw/hlEkekl
+RtL5nFJR+hpFd/++bnS3vjMZ5SA5wkWb7TgcpccZDPC9f7U4jHrA2+UyG/zy2BCMWbNkKCc/HnV
bNDz+gHxMGYOellvWgR2B7t2xVMcnvs6FlhC6Lf5Xwt5auNKqU6tRqV7od9ZiOCLtInzvVP9gBli
HsP6NZalruKN+L3nmHw0HPe51AAi8+H3Nj3yz63oKDJmQzdgO5aWELaYKq5m3ACqBR3cCIMxxwiI
GO8kDxe02Vlp8YchRQ8e/Eg2A+W3tmcXrMYeKsBhDdnLoy7TaOhObJY/bLsj/kX62z/uZndu19X1
WUE98fZkz5/p4B0abbRUs+aCUtR64IWTSPvCa5Qp45/tgnptzvnC8jnSaeW0qyNZsskTXgNv8gol
qevzmK5u1oZarPv/tHY8ZktW9kX4jsspv+Tw7Aiq9OettF1ex0AuGzN3DWWlHBh/7ncq8rzcpy2n
vXJQ0Hx5c+qFh3t7touN8NCFVqjQwIBJznt2c9lS7y9YLaMmy4n+07tISlxEIgENdEWIwfZp+JxO
uWpkCMKKisjcA0Rbao3fxM9H70DUgZ0AVjwqoLccGyBPPDYbFKQm02/ShhMatLqQTxusAnn6y3ii
30VYCsisKtdfCTAvuAQ7XmE7hHOxsrlwXcq2nBK7xoPlGAsaANd/Bi75uPj68A8aPxolfomkMgd6
Zk0jMAlSkPD9KgnXYTt4unhFYWI4Ep+lfaVoZTdbCUfDKZyP7V2sHBdxaRUDmszXhPGL9rwU3TKM
5sB083LDsLuAENvOJrAL6EmqYFPgYujzVJz0JPxH9u3Uo+YoDUXk7oVyTHTTCKfz/qF/2aD6Cwih
bCx5eGiGtxP99C25NhtYGlULqhlrSZ/f86cQMT+GHM8SUNCVRyoTasxKDdqguqSPeiY77LrUOIBi
CG9lfmmriks5ZJ91R37oCZyxhkLlU93vLhgdGWm33HJoBaaMhiRSr4nts7EI79sPPkxMkWVQ8jCX
ObTbkbpG2uN+cyGCVHZTvJtO9PHyzD411DjQI+VOOEGnmkM1RPT+LfQHlb8Ic3A9p8HTnPeaQDJG
Kete+9xGKpNzzVstvzoUES4Zyb3q8HyBbbI5rO81Sw5gNnpgeQsFypSce1rDRDZ1okuZ/QJDLqqw
rijnok0rk38dvLyaoh4R6HMIaCJrF3T/DvTgzphCLsooV4Bj5xiRbBWN5hNGicfM1ZFQE5yaGbeV
fM4Tyrz4IptjEkkhg0F2ln6D3vVS4f39rR8SoUB7WZlJ2yF8EXe2cgYst0kJx8fRibGag+ZkmyNT
L/VlwJbM9OJuUhmBBjITtL6CjA2yfuBmjw9VKZyiQwuHtfbXqUZgzEQ+JNVodFRsPZ8O91zUjD2V
5ypvgmYbttUNnD12RSNVn9t3RQ7fP2qpMvkAupL1OtsBH9sw3BNZHbCinybTBA4d1jfbN4FW/LcB
fJ3tkqwZbMHsIwXOuA82VF6DUYQlGFqy0SXeysUV1rybti8LsXiMNXUXYY9p5NZAMbUMmXHV5P4V
+Q5DvgfL65qDEqlcwzCLtrH3xJXkiGGAn9GdXqyXNUs5hJSL6wa0/7Tn/XqUcZYINmwNVK1Inje7
NBHUkbi3SPI98i4HpfeBuChrAwwOhF8VcfjUQlGNiRTZCVtQ6ou59GUPAfLKIbjjVTTp6YpR2rR4
UzZKjmRuu+Qk6x9oGko6dFpOaUaXts94vQlmnYRZpM2wUAfjvxEE0Bxxz9+W5sEkGm9S8c9l7DxQ
glJXDExoaHLaaG6YyNw3OXERWA5O6QLMdoTbK/lAvDrwyHBTPhb/EvV+uNCjUHWS3MsSa9IZn0xn
sX1iPKq0QD9VdZ/RN7M1yRTotsIpdab4M0UebfQpxxt/pOhzL+VxadRu+z7vc3/JZpB06Duyqu+K
B+Vsqz6OyqONy/Lh9i9+o9reDXcTJRicGTRER2zVvZ4lLx2E14eMf1CBSryDFSUK7r2KzpnahhD1
WjYFhAY+XHP2/v0ZIpO7lrYS76QKMIlU16Um2Rkw91h8trcmgpE0vXfVghQ04ppw/2l7KvuVemsh
PRx+cqFt+4kzKCNpNWtumUFicE6wN+8v7XcjYjj363WjpaX50DF2OVxx9/qwvuy4wLYOiLYHs259
oTbPCksNhmJS23YbYikjdByDLU68ZHE1sfNTdZ5LE4JVqkGiduzfa/x212aVZQMNFGHy04ugjU1l
MEpod8INCfOSuQ3Z0oFSytJufsLMaVaW5vlZRud8rGu13j5NEXv6csHGrcNZGp8QymEbBziFqKT0
aXmuFODb1FfTT0+p7Fu1g6u5AkFHbjcFLG1E6xq8Zqj6xIoxLjeB9adgkfrzcHmoetWyuVm0JukC
Rp8vXM/D7ruBvZIX/PMol5MpQp0Burrtt4huES4Qiw2nfnOOX3VWo5NMy4F7gF/ofx1YjcEMvx3G
C87/Eha5tji9DMNmbpznptFVKkVyDKJZCIvwJbkIZUbf6UrTjcuC7KtXIT19UZIe69xFwuUPgiWI
BcFC1CuD6f1roRINSG0M8ZF2x9Kf+bqlhT1abqMSBzMug9ebYsf/oxZaSzpaEZVRNNvZeHrhwKfk
GdylZ6Ql4/oxP0EFatCB7DD5K6Y6C8C0Bat72yvVsrn/T1GnhFNL2OWS67jcKEOYqi1KRgcXMJke
xKFLe6NrKe6iyGYKVccuJNii5mYeCNpwveg6Sv43sErBcsJ54sV+5Hq5/YLU9zjiUB62UtbZYHmS
w6APeDAzxsum+pguiwgDij4Jb1f8++OKmePqJXUHMCTt5WctnMQd86300AxuvHf05wsam0NS70QL
GURClO+pZnPivJwyNz0A0BCe+hDGF7Kc+kdFFFwnQWd3vl8jVUUbpNMXs153sSr/BU3OzesSlwbc
Geo9DPTP2tu1u6zouKXdbLs9bb/0H1A8ixblvlLpHgbRZzI6MKBzc3seA6ZQqphJe6dNzPZjvvhw
zpfQjxzi9QKi6qlaZGQzyHxQRzU7jmItgkOGCJoONbV2MwczOMaRKBcqpEXLxc7xCH/08DAuPKL3
gjdm8dvgk4JBA09nPtysoqkIqxzfBeH9puN4+f4XjtB34wv+pJUc17bmBIKUovbHkuXSzcW1sQy8
8I0LOFHjnrXwqamRL0Og3jgbhRUeJ8RpiFColTLtZurm8inKYbA9zTdGowJ0zHQQoLIK/nzOOON3
FcvqsMbcQkMdZdA0lDCcskQqHxPO7L0yCzkqZPRF8v7hdZAVkDVYEs2vr3Lz8qT08fV/ixYERR8n
f8oLwKWgv/tpYbPQsY5g0ED1HbW+xZNcOZ4+5/LL8yLOonXcU8csZ0mYyqH8PI+5G3MyxcOYZTYu
DUOhz8roIKeON+Lz4jQ8IeyX30djYYUF0ywkj9lZXCHpXy/p2LGnup881BL5QTMHnw8UtsOgWy8n
vwk7R+QtpfwuKl/zdSAIrOoVowbyP52D9jfgOtcC+TwP0rQd8WQJVkAFHy51S7HKHVVIn9eeDFtn
Fs5Icc3rrFMJ+6BmKMr1KrC/GvtW2CPq94xEWMa1nHAribtAJREAMjlP4ckeJdDdUpRd8fQKA1II
/Envf6MmgscqBt2gFDSC1ZYdrM7mJUouhpOeD/BFLuppMuS0HBxLfCFcQX5v3HweBvjL3PXpQUCk
S24LuHCMQQ49OXs1WIJS5oDCsSyJ2HxLaBMLPZvKorcDEx6EuELvc6ubCMK5E/7qZFUQ8Texl1so
44NRIvnmieHdnOUTqQyiNcd2xl5U2p/M5GAowERg6lIh7n8CBQYU+1GRfwuKQtyhQJHfUVnlTxMO
PU2fFJGhxm8pG23DK/JE3Ftl7yO4RirdiAPwEkCm7Ub5SMLPyP03qq3tlC0PyFnA2nnvMxmvkmu+
8NFR5rTtZ/HF4fgq1vVn8C1AUHzvdMv8uFKM0BdLkRRHFzewOViAL0+z38DuQBU9E5gjSNnlY+an
WHzCXvWJ7Fhq6jVJN42lsDkGC+k6fA9Sv1KxWk4Muw1Kq23guxJmDJmOkqUmlEcoQFMn5XfLMJmQ
dg4QaIl/ZybwSXLfoqcP3sxzM3Q8VkNU7BuNVqnjcSRj1CH3lCaTJPsy5vh+vfg0co3Ovce7yS89
xlIn4YEZmOoESSyYp03UXTMO+DzjT5tP4yW3Tz8P1v8cga5tHI/ZBxTVlLue4OCEbaiLxSvenMXq
hMEdqgYR8Ki3lfsAnIU2JMgyXHQKP5w337cWXuGWtPdezTv+olcF5xvLnorNwnNr/PtkF8O15sak
358OM56a2KRLUpmGwaKIJGvMM0ZoDuMWgp4IUIpbNDVTvNk7SLdljFH8LKKfS5KCuKwOhmILTQTV
uRXQf335csZZh6euyBPB32noYopgope3sDxkM++O5bt3J3jF9yWv6PITd7lATNK3StFVlJt2jwCN
hmVVMRTT071kQRZhmb0pUQRECK7vXOKUhWR/7fNfkakmJreVdpoR3cXl/ojUl9Gcul9852qo6zgA
EdIcUb5/w+osGuKER6wKd66hBuOvj9TsATonkAVaf1G5/xi+3UfZtibGtCg1/WngIyOu6J3uYZT/
VvLPB46crGiH06r7hUg+fpA/fliLQ+vYPplrW01PRnq/QyoT1NFTj4TA5VakZYg0MKhP2pm70JEb
yP8n7JLzQfHbwkwjVGeVUfTi+KQL4aO63fMDbWexuD3jy5Z2a/ylo6POeqopRpWQFlMLweXs/lhO
+dDpw4Z4+dyQBf1CN6ng5xjos6I91vTFRE27My6/jXArawwAztJFDXIQeHXOJthFFK1NAyLv3Wi4
aD9xBdkGc79HFpMVRFR5OU6OKvf8JFhX1WzsjeTbE3X0GSagCE5WdZL/WxBHyr543bUSiPBDxjCn
18NtyPbMj5ZZphKdSWJpeDe5vJwEBtl/y+L1RLLD0d6ol5AHuiPE71mYVYYaevsYDgDah2Fu8/WL
KGOaelCgs5sZnHpXvDsG3+WTmZN8MrmUdMS8as9WhzzJqXh1aMvW0MpNcoNDOWUZYEuEQEimKaaS
niFJSTU6dvvs2yEc+4clnveABGjMoCjsep5GUJdLjDPqc1gmRQfJsyv8SMGlbQm8rZvsACBavRWQ
zR4BF6CQ9xsmBQ5dD+OACNmobrG2aOzk3guIT8JKSWMbWnmhuMmXZ4uPzGbJLr93a/G3Iq5PhQJm
yPCuAfpBhvO1XG8gLdbpN8SwSs/LvbJV8T3zxq9t33dMM1UIX6tnd4uDtkxspfTBmkCGKOWlQnAz
nTXGKfi1NaZiSQA3o+6V6mFCYYB/JPbU1EsgUpfhG5CnyOOLRYe9fWtUE9rGRfL5PU+JytsJ23a9
ED5QqtnS7VQwhclwyJCu9TJ9HY6WlEkCNV6EXdaF5mukLXrl7e0BoSzhBw20TRmojfEyNNoxVk9I
Y+ywkr0OBB2h/8Fws8U0Jp5gOko+y5TS6xzkWqYhM4EbM0h2SyXY0Ma0zBQXmwj91YBmnbYkG6/N
vmWshPMphCmzYJmHL5/p7xfqRLQx7oNaABTpXRYUsqLyBglLavtpgQPq3dJ3en2tYeVceboJdpZ0
+27I/cHllt3xsmYfL6AV4SqYeU3hARSHHqmO5BGnvjIXgSxqhDNi6d9bW94mcHjwmENKq++5qY7l
xqOAITpcSA1a2hVGYb80X/2dSGne727ln/sUladEiRXKhSxK898S5GBN/gJFsOEshg+nqUQwKPXC
wVwWOUTiT+vvk3EvcHBEsU4quo5YE6KQAfsL/JIxj/ByAA++jeLXXJcTLddur/9Nhsmy4ltAw2U5
6ZFkT7wJiZMK4jHtYl9JoXnct5fwooRFY31l7hsfZL8+oMmlaMXt1DETn5+McK3sqq/hsXsXSkIn
M9MqC9O0TdD/byd6g2dieOVahXO48avElanxX+eyKvBTF7u1CM8uSrEzW+nBJ23nyaYbaBeYuPT0
h3f/jiXuZXgJ1RhUVW8akePK2u5p2kh6OSdD7NhOPUPuEgOW+dqeMY8OtQylukv3tB+Zo5KCqwLk
pusWG//1U8pQlNG151bupMVpDC+ZbH7uo023vSJE9JL/tpv7GaoB8VvrPoazAzinaip8nLwJNbzd
2jjcqrqAgWB3vcCrVbx+2X5taNgqYnVmEE8T581cSKE+LTvkCtEyNdLlW5KNZNh8ZI8sMYu+L1Hh
kNXJUwyaphr6XP3onbx1M3jNe2cfDqGuuE6XzG/pCkpi/lAE5vb+o07fNa2C9TvZW+wiPJtI2I6C
wImZjfM8J80YyZd47/GW2JSGdPHH5LKhsnQeAwgsGTkoOlNdpkUZHsVPP+DfHcAWbBAn8ONn8onO
JTicsUzq57fP36OXZy/U6bbuTtjFaFrL+jtygTMpzlN2jjTb7yYnYqKchH0wj12ZckJ+GcJnt/GS
qVz70kF27X3gaBhH2ASE5R43p7u0KQBsjAAoHY5R9vvqvJKBqYkcS9gl/qiYutH+WS+qvnPaCwJF
jVJFOwnMzzWKRY/FuuLmBMutanhJZeO7yPcWARqUg7SEfW1M/yAjlE9UnC+r5S1ABINem8UgJqL9
C5TdJ8tUZviKUBfrRlTBzS+JbTpsp5/STtno1sO3PHM/03NkqhfMhjC+vEYidCzdZCBFhHgOAXxD
fO/40t5bbaYaOwCCaSlmTJpF3B/+jufds0N5SD+Hw37N2EaZj+gPCn7nfKQwx9rbNErDSfKvK49a
7LNJL1T3GrIOngsq8rf+R4Ge+HF+pWntfxNiUvhdK+/fLFLKUhW3YgtOVEUdRii8ksdzpyTj8sYL
ZV0hTiJkq8z5pJfRSsoY0GGkXKY8CDA2mvJ2iD9VVjRK8PJR29c34IGscwtXiOntyewHp9zLmcTI
S9ASNbbXNPVuBSBLn/Frymsu2GVk3OA5xTHMWlLjfM9MngfNp0kpNX9JMIa+HJanKPkDedvDLoqx
ggs3T1h5hNan6IamQNpnvxp8ZK9SqGvcLp1IBEtNfunLIgMW+BD44GxYfZTMcl6c2KLZTqjEhAkz
GZVnoYdTc83DoyZPN/7CV67zTO0GZ9jJDPLC1BwUgE/jRsqww0d8O8QnA1qQP2zBjXZEj4s328aZ
vIUNp+wpQwJ4qVsgptEYUhkaHxMuW+kYeNcIwVkgBTGCIpQKwY/AWWhSJTCYPK1dbg+VunFj/+YY
meaTKhD6VXRs5ltuJgBaJeRvrGZ2/cUXaPb2BCnJcblRSbRFOipUmyFYZDOuJ1aPJCdMqteJFaAv
eQORrQvB8sD/K353YkD+3Gem+b7B7qB1EbdTlJqe/3/t7mDbkzuo2cRimw4nBPi3nEy9nCMy3DFr
B+ra+JUYl3bMaPw9Y9V5S7cQkf0HI60F43YnqtkfAOsAFXeFDEmXKh4wz3VmuP07vQ1qCl62WRT/
ag3gwusirftOOs/bQIE0NPRYw70s+acs1EpKnksIs9QW4M/7OUDJPcOefCdHyQKghcgSeFRqBzUq
Ys7Wxu6r7vH9AnXc2UhdD/chc1gi88AwJykuZV/PKJOihtcLcrtUaPSLp8M/Te+gmS/U7mAQqSJI
XUz8Em4PFyU5RdHERziqMILZ6iO5GR0kx6yrwMBlyaEmnX172TT/87BQFEHNZ+OS0mDVSp5Vy2/L
0hdUu/UFgZQLcVmK+bAvhSeO2yqLpVStGegMXN97hTo59YFRzqb2/m+sR2bh4aCOE1cb350Ktd07
yfrggLd711KPSI5lTcHD3OHCOPhSOBZiUZj+cX0dimiBlP3h7x6tamKDid3VlKEf4DYX93R7Bgrd
+cUDFpStQM1ynX1osctiLB4e1ylaweK1Gm6nuM9Q/iMy6anNULUi95rx2Hl4wCKavNlxEdFTjHUu
iDjNm+tfavu0Slo0fYinMHhHeYBjv4pg8jkgn65yI46zMz1o4bmjejGrgs/SO+55wmR5P0ioR4Sr
GK4M5ukDYb23pPojIyIMHi1lfmTZ098FOvJjFEoxhKX+vaj81l4gVGgL+NOYV1hwykPXKR1JGcNK
CywoGtUFPnI43vtUeMCfielursavGPknECE7GzVB+2jhSQ95G4N6MZP4aVNEgG+7WAMcXGFqKHHy
waGYv0tPE4ms1wAiRSZbjPdUZ8I/hcNZq0Uw7pSd2WN6tcY25DTnAMswPpymZg18gl89h/A1GzKG
+MfDMB8Jl9HOzATZIfV04wKgj+pjXofYQD1jE80UjPvxcb+l+WMtEIvUggSSqwQRMd4uxuIYNa6N
429CnLMb3UugYCHLvs3lOjCKRcBMHMA8LbVEdR7/w+B2lCcxn3nU/V154xT5jVV0irFM8lX4cSqw
jj5W6vH4LVeFPSe+soz0lNBlMHFLa+hwnLR1bleYivH3bK5XdVhslNpR31RjFA5edT9hYLYWs1F4
qLewFzw64h3u8sqCeULl76wJSdUtGgyKRJwdfSZB9XkpjXfGjQGgxmZmsqSn+uU4e6u60u9oSJVW
XOm8GF9ylG4nm+KSCr8BqY2KR/Cx31HHhGTZmHetxrDEZX7O3OwnRYQxlHFzvlnAz3bgNWAvOKGS
GvPPY8apFTHL3aszRL/KwejKtGQXD1tovX7TQJk7hoBOO4P6TqdhP+uA8TC+oBKk4C76MXkOWD62
cIhP5jbOzosOjLx7NfA1eAWUbcBOQYrjdjK+xp5ko1TfSY9C73JJ8qt21O5jMr0Dl6TwvPOt3lG6
oQc9v+8Ih08Kl8x2pzyynXSmTuKdkg8uWIEqeMhhnwt4errj2L1fde3hzzO0PnvvS8ykyRXod2Om
LUYaE4VCTqM9K0qFA9KkHD0IHuNU2NX05pge7HoztSpIlSZL3QsyRgfRr10YxIKP/dtohAmiulkn
4xxWD9Fwgw+w/GkzVOqeUQ5XeuPQEwNzTyiynW/ZUNMMq5uD1bkSDjpj+FmCucDilAATsg7pXeVm
fDSUWY0pizcjgAtmCPJMe5BasfT0sqZvcXVK+Ek5zf0l6NYM3tDO7HKJ5K9tVgEGuZ4ca4ljkFsG
szJqw86/rVDDWZOg1AqV5Fmrf0V5OdLYroO5Q1fJAJWP6KrxSMx2I8dT0n5AZZXsQk9vzNhkk7bN
OlczOO9lPWCSTHdTDDoI5tiD8+AhJhVZtVpUAFq0WoBVGSam7ZygJvp5B7eSgQPszIIPnCGiq6uC
sRd5tKkVeyo4JCCehpyDsgAZHTojLu/u3ZMWYfU2N35qLKUfmeTVMr1mTvxn/PWw6tHPf1QspQcl
JTaWJ4nn669xoIiw4atcmUNXg2PDy0RZNAu6WI+wmlwuFyWDtet2orARXMm9UBbIoCh5Lq7+AZo0
LeOgsPH2ASfMf++XmXEsDf14ybts/nxtPcvWBXTJp3OmyYftBSYDkoq6ky2GuXN/Xgz+tL5eNInM
MTTptrbUlysbbhtBDpQdWpQVuqIFUQ3Qus/XU8W4JYQ6mSx9mwymUuT+k8GzdGzVUqBIh8w8EU7k
uqi1JKI+c4xpCXUc2FxaaAxqwBjVB16REa7P5Dk4qHbRh2jxOTv8e+OLhTar0sR7zspBxehXm7lb
5pJikhUobVKm/ZYZ02ZzAQcj/5RslMtTBm2IIyD9mkWtKSggmVJpH6mgBrmErkuN+T/EW1VT/EX2
OIEGhW6xz9zaeE5RT92dLi2dYxSTxrTR5nbauPvCsctahoN/BZQD/55txv/5Rio1lh6F39xu8cKH
hRWU++dSzth9hM+2Yjs2vC7CDFScCQQqgLtwwqNo8yQ+m5pMcB9r3ZB7NlXhD/ePCy4Cfp+qcef+
oBVWLO+sM+VvfUDi59qnY+k1zR3OfuE3MTepSM8y8uje3QjJbfDLqaTp3Qun/Yxp5psvmYs4CIzI
IhFlbUNG17NjHaa4WweyHJ0NeA0/b1lsJe4tUO7NTvVGJPiOBnPBi2bYsho94DDuoK6FkT0pQW/7
XEsDmjOmludY6WglPgaHbSFnXemi8emQkpIF9BSkEOwKUGgtJqyMKdnUQr97l5BCniJYWnKfUipk
RnAomYqFoegv2RsVhPwQh0vRzxbhfbLNs860TPQWi/aBWIaNL4+2glhBuvuSQloBra2YZ4GwPW/B
zvXs6BF+I8TGgpvSQkyB+dkpvMFH0ZCQYwXwgrWUgqJxFwvXYE1gCDiSGMrYddag6vGc/xO9Wtc3
wNb7BKTMVes02wZtEoLkap1kEu2ftfepj3bEFlDTTohl8VIw80+DtHjcaKYwnbrNJ64uuXoNQrdb
UuP8xQLwlYwKIIsVKYAc9CAwI1EyCyS8YZAQhntsYEJmY48BxNcc5DO4mELmD/+2veAi8twi+MH0
5mRf1OVHBv1q7EIEYqiRbbsWAH6g97NsfvW2C4+18pNlDbjKpPvvSq2ab1FSXl2jiPjhsE9L9KGs
v0UK5bI9tZYvuuErlZ229tJu2QDCeeJHIl4rAsX/gzM5awAQpeuwqzZwx9gGLNBt7szdTLWlIxFf
j2dxsc+mS3eJeQNYu7EcIadhqsfSQ2FLXd/hFeicqJi7qVGzTo+67K6VtecdVC8Ql7RgSCSCMZxn
fhFzZIlrkQ4bpm4YZ9Hb01GatsNeynCWEsGZssoUja/60kPCKEJ21aqfxihghUsoIH2+2t/RQjWd
7eKSAwJUvhGHtCx078a6bg6qItmoLrjkL3IDAbH7espBZWKnlJ8yfFgwwj2D1GB/TO1npAxtzMmA
rBQk2HOzkzcqvIW7ZL2mvGFUzUdxYhW9c3LS8rDfbTGU+0ue4K5xWnIrhwkpndsPWpCQPSmeMoEb
BwsgDK7xOVZLywKN1vR6P5FTcZDWFjvNZThPt3k0XXsd55JF6w+/ggb9cqLH+Jib94obJMiFO2VK
9pWp5AVs+5uxKGbrk75hZ6rSI0gisVteBVZQwuQUNmDz5emiCjuAl6bDCbgjwELSEn8MA3Vpcykp
m2DVd9nfrBxCIbgN9EB64ESLKhOpZ2uCWHtR4VAjxB1Ftrv5AG7N/SQvUJaskDVF9bi5RDfGPMCO
XDk4YZVSHz+vGMAe+eyPAiNqE4BR6TOTjOvM89NUJMSrVLrwa3j6W/Fg0NJ6s5otPWzyaSd60GQV
+6JBU2N9908LKEe3C2MEZyWNX6VesjAbsI7MnTHGCiPhZF/R2yQoMPWPKArOMX98AktMj6fnboBX
rKkPFBC5TI9ccR4yXbKZuHtMlEbHEuvWJSkCaRx6fbb4OjhFuD2h7va0AN/eZmcank+pIgdR0e/X
hz/JyoMZuk95OD7Gagvf+nRREEUIIYBxt9tl6eUl+MGSY4Ae0Ru5zZnJINb82HR88YMuodr08itl
Xbs7mTSocQrWD0mJHTUGInq56AMq6MnVUBLbK61xXLfqV8JGmfcLTS0Mc8X9sNq+aDuwPae+2m3C
CBObGv8DmErkd4duWU2y0tz3NulGeUGfpU/hXgnAuSlChOezAMuhsy6zW6U1Rr+qdZ8l8MTP9AdT
g6BEdSacCTTMtOCJ8GJevHpS8j3ej7Epv7Fu8VJkuODK9wD33mb7ctk99ASEv1EZTn1915o9yizd
6Pyvq7AOpiZxo3PORCvpUSbTffU/W8j/xpIBSy7r/inAk8nSisRIfRuGXET0TsSIy1py75JZpmex
CpqlY9XnzYKx5kreACug/cXLgxm4EBVj3cC+dIpx7BvLV481huBA56lSR4b68WmI0vLzZT4dIcbK
D8kA6e6IEYTwQNRmJa8jxGgz1X27sUtm/rpwuwnAaexAVWUb1L+cYG6/4wHP6tjJu+hOYcPfujXp
IGDM7K1SsAVDz91ou/g8Iwl/A22halYjuTRTBLMPzrZmou3n+mZR+84F+QC0fPyGM7WionZ52KAb
TUGvvlJ9/asbGyyGLqiOX3EqbU6e3WCLoCC828KMIHGGxln+AMH41mcxQKSMCN1HEv2lALpnnHDS
bvkF2m/o87lRhSKQJlNqqxjivmDlB7nr4XSJp13iovhrB3zCxAbwogePuPiuzHe0Dv3ORq5S/juP
V2q+JfnjCduL8/mOOefLDocumSA2yF8MAj6o8h9N1uxN1GizCDpqZ/jPbbh9CV6GBLs/ko+U8+Q8
XBzrE7JG5R/yVV7MauD5grhFwGkDmG9kqaW1M4XdUD7o/4TjjIzbBfiSDhgPE2nTVC0PHgs8zZU+
Y+m6I5qXaC09xwnEXv96qU7VhleBRfCgbRsEFJjC8+9JYT8RVI7LUCCzE6NU3nR86bVTgUwmnng5
tK+5M6If/uM55e3iBdDUI1cas8T+8qtOPnR9OekwGmeUuxXO7dquitYUUhxF4MLPbB5yP8JLfTrE
NYnCekDEerr5avhPlYd7HjqfizHDwADde6dKfY6fmwSySSAf6wt1QiQalRKMy1686ORkyG2PwDRU
nRqg4pSTLvnWHiRj2/LEhXPEeMiHrYre61+bQV4qLQrJo5kgP7tRW3Odmc9C02Et1G9jROCbA5Wr
7EgirP0Z+v2X4v7XG7GgIp5/9udNUCTYmi3SKhhERp3bkn200GziZibPq+jKnsg0BfMovMNDi3Q3
FvuAu1gsFTyqvHNXpJcIKC32ipnE1t+3xXlqJ31Jmbi5Foq06A4RadUkyouzJRd5G7QanetxPw0B
ysqlxN/vMIhv3f/nC7U1898c+sVLDbAii3HuNIU63UclnmnX+gwuXev2K9wtmi5SmyRZxF73TZBi
FwbPtsfBvKd7enegJwhTdVf81wg+O35uYCZzqxl9wS3AnXDrszzQAGhHt9H1PfcDfpnlLc/dZdvN
aI93mMlnBKtQnHsxJ7wSbGlbMLgSloD0Eg4pO/SS2R6/CKIlsDG6XwyGpiZQp+pMBcXEi0wGoYWQ
B2/GkW2FudeFDvBImzZs1MtEPTc5RKmXT40zXs2qTyCtZITdudGLiJkBgmup67q5nKfy7XEvv7/K
R2S9y1I6cQa9HihQteXQeCqb8FbEorCkLQEnMwRiVLkRdRobcjqP5/VrCvoWdO33d3FBlV+4jWTQ
IAu/deSS/eHeu2ifqCZA42Z2a54PBm1bs7gZQTx2xDrurOAx7ErVc+Um6MltCyUVSwXcDLlptdOl
HorvpNXlhmiuEO9w5NTsuaoLlFTlRCInI9vaygRVBwg9A3BiJdvC9h+x0zW81qq8YeCzOHIj91LI
MYxcOvUq/0ictxnHj/yhpr8V4qlhy501ixgR37rc9O9bRMw2q7DppVIPFAHWNeSnv4a4pjHSMZBd
MmMHMmUioqb+xd19CxydoRbq0h0jXBJDrgxwfGWdEPTA4P2vVSZmY2rBT4EuGZMPIlnj9F6j9KHG
4GPnE4r/4Km0fRsZjisxpviCKVSBpmjMtPkznATt6huiRkxlC8ISl9yulo0x94bxEC8sE1uPbPNk
5aDnpIMbgLqRNJsP7kONmgqIYAlRcLUicvQbJQpTTaOx6AqUFtZd5cWMjq8rk6O3W9bQqh4B4LQv
nkJcDmHvEiTadCOKmaxH+zHZ59L6OrgWvA+Ls4cNjUXPRyM9NT+5qa4b4qawLOCQNw7mycCzKH3v
clqp385NGAqJAACmYUtyzT64dz97h75p4x+LglwQkrL9K/o7W8D98M4DkYsv9GbyzfoeJ+oCiPkM
KpbHOPZdiOuDhv/SKU8eSnH+oX4OgYzRMYa/IW6lM7fAclQiObt7AURe4FrhcuAmArX7F4wxz39C
ScCpVd1jTSQOVAdTvgkYYu0Irm/RRDfAPfqf2QXCW5fTwTly1ekXiCddehPu3CVRPGsz7jAHmtAJ
lVX/563BGzWJtp7gvt06dr0F8A5vhSLKmskDv+VDnQ+mp1JrDeRWBLssKE3e0JdvpHmdoxkfAmR1
UtG3AAsuBUB5Rg8+ReBpEE6cG0yJnSxmUNHDvCzNXXZPLuHKk8VZNKBwZFd6epsRjIa4FoluTNUs
nii1SG5dS+bN4irP9Ve4njo1MWFrCNaUe26SSjCW5GrX5QUIftsAU7OCv51eFqrlyamo/zZhvy2G
x7oIW/jiAU+3McHbAYRohFiOpulRAQrV510+GsPKMLRZX312ul/+2gum2QGjXiCAIAPvJbsT1N5I
tdeLPyVzO+GDnrjnbwjsP7vd4joK8PVITcKmo2+gdE0JCSGjWesOAfIM+XhuwaSecEjguGrVlwIy
N/UGkyM7/MB7v3LCP2phv8Po1mJ830ZDDRqlGGleWR8Tf6VH4+G5elqS0ZCRHHzoRVkAayvyS2IB
S/80P2AqkvXATijeoqTGmZKQ25ViOVZ6xbiFkztckybMUqjb+Ui49ZvoJBXwUNWqXfQi8GhJA7Qj
eaiFKZIlSf5uRtJBJ2ksBw/pjsC2kr1KNmNtj67Rtk0k7l+rbc++eZO48iZhR1yKrUXrIj0a8+B2
zHHE4fyJ4ePlaeMEEtbDEGVbC+YQskCSmx09XOmGLewKrnNGy3zOcu1TjVuICDZm1B6lIbdZphSn
OuAg/eJ+pjO4vHuwUfAYWxrCiAprPSZm1KBx3mFHJmUa/iOD3cXDzqhEt+RDujJ5XIXXFuuSCsIU
NoExXd45BJDA62Yd7RmQGxPGicINRqqae9crvZj6KA+vZDn16dfn5zV/HqDrBTasy0aEyjpL6mFv
pJIFGTwNiT84wt5OO0ESdTMqWpUw8sZKFUqO7gavq+gQJuTyeFj4knG7a1Ll/QFg4FMr2ErIU5m9
425SIGONrLu/a6VlrruiLEY3jMlX6qWE8sxrXmuV95BJ4cxJPWRbjrrGhsLyo9nlxlt71h0St+mp
JP71SsJQFBZfGsfvMUaUKlkIFE1QS9Pwbsi/VOGOQtPyYtYJ+XRKOrJOJKBU4eRfskVgkjloRVLv
E3hnFqLvnv2+jZ6Z0DP+QOR8qf5WkVwtpJCw1zxheEIiFZF3NGgeWgIPUMWKNoSFBC7Vs/Yu3M/o
fwX8wLsy1VXW9+ORSoaB5WbpP7eRs6vIHSe7nJk7p7u008hWBsa0yO8u9pmVpaeQFAp83zR+LMBn
GEHYnJxfVl+8MB3GMWE6mXLwE6giqve9CrJBfxJYWBHrX7IQREBKEpRHO+IqP3fCFfZ3DO/nDQ+t
anpV7ayk9KKgV+8FQPWcPZog8U3K12OPPMQdEVHmZJiFPZxoWzvrReiYLzBfWwnYv/T4figlS9O1
vVZe4NNfq90Pfikypi7Kv0OLuLfGJ4HdCjx32su8z4ZHu/vI0WxHKybHLhmGMKO0RpR2JUkN/Lbg
oIL0WOBH5f4Mg1tU0cVPC3jFWbZuc1mdQsIj9vRCQJvkR40hQielMzkJvqtPja1MxohckrLsnF0j
CZPdjK9AmJ7eYWqywH3PyjcShzf9KVVpSR11Gg1ef1qjYWgDcWf28b1KUzBOWzevlueALZEoTZWQ
OIQvRX0SajdToXGDCbnI/+VTOIxt0DO6fnQYQ5FrpS/o1jp78fyN8gzR4e91ojPR3VnXN6NQoXiv
3idLCeR0pFxnY4Z1Y9pQZpn0b2ygDhxoXV8mYhq8WJE9h4MCeO3ZjXWgHbeKSdBCzV8/X7HlU1Lc
VN4mDJ9jqWjIu0zWHyvcsYxRGSMXSifbvQK21E8Sa4MBonAOgAeJPiNthLV3PPJOKopFMoyMxADS
59dzM6uadKR8xt+zT5QguZgEdbpsd0mva/KeceKJefuPFA1naUOgWqrx9S6tLioXjLot1YeCqYSj
rjdv6vqdi42vDxsOB1u2KuyMTksRkn7WVRUKNJJ6xfeoz2d2o51TIbYNId6X+hdiD7NUNFVWy/cw
x7XvE0YIWdFpkZULZg6jQ36dNwne+lKZn04TDMIx9AV1RAM/iATviUwDs+KFICtqDNlkrTgr/U9C
BYENqZi04XIpjs4A+NLHa1cTUn1W+7wGQ40kHxZe9OQ8jsrIxZ2aKZQyjnm4OxJberjp+bLgSc30
HFdiWf7f7gXGh8pvDurmqH2/i4zT30R3NXHEGUMCqwINfLiyRjAOeQUa2YtvoeNSpUXBB7DXeKf6
W75MxBSdHdGo/erMmh1XbhQ7ptg5CLiCw0ssC1Tjmiak/0+4edEFik4aiq8v3muDoJL/0X3oqp2h
PjCzpV9D7QggY6p67P9wZIKFlLDLtp600IEuHHaqmKJZDiQqVAxddPT8NWoFHXDpBW3s8Oc3RS41
bpaCBWRMweZtZFyrTtoZ8cjsn9UjexoEW44lqkgw2/GWw5fcpPJIVbnQAW9y1VQ4ofrQ0bmWhPQX
TgLr3R6Xuq+FEOUMzV5hmgNE6fBNj5culIBDsG94yprEouEGYXaYnlQETE/JcIy8fCoClNtSeKyI
SF741ij7q7bFyldOfX/gHBKVz4AOhIL5ThXnTyRYJsIOiOVuzaYcMh3TMeVH6Ev8nkZ1gxXx0uKM
Ek97qOZus4To1vWGz3V8Q+n8Nv32Pheasw5wVQGxIqhv+lxgTYuiPfhRNo7zwviEtEsCzuvtI5lT
q+ddcpweI5Dxn9tgB6t0KPecIiLeTPzJ2ox/2osTUgHMUz83G5xhKvYHZE275vlGFWODdTn7MWQh
OeiVr2hf5p/p7r7I2c2HXWqyV5NAe8vvRFm0UKDrCyagNXAnyoh9P0xnZAEp7O6CqPYF/tDueAZN
kxe1UtS7AapW2seBy5dMFylufWnLWpgFKMtOWIgGsi068KWkiRLfZDcXAcpNSABfAdHNLxWg5zok
24d/w9j8EmZFX94NtaVqNPqWEOIQRioTnJZeSYbesTZXfxPKPpxa2p+qQoPSRm+0qU6dPPWo0x9+
Lsfgvfbqk/yP/VqRQPOyO3V1K7sz4EYRLMI9za8FnvtE9B4K9PWkCwceONBxNRB4tA1Mm3npQts9
zDMNPeF5GM04XSvLGDtY9HcO/fqKNAnVna2ExHh4ZRJW113u/XJYVbu5pLJPU4xr+rtQDCL7fywp
QfPmtpYnOkqoNv4bXMHxlE8ozGzF/23s0WmeewIpzsFI42dKUMAu3O3PIy/diAmtyz91P4ZaIcDd
ljhKdKs2MWMleFniHU9LYXe5WDxMBXrVsT52xrwlsSvTUeqIzvBsrH1HSAKQDhm8kBxia2GDUERs
iMzSVQ6S3NRjsCL/C1vPnwyZ2856vCufKC28N+WIezC2lBByloAD1RfolUfCsH7Ho7nriuK9qPCh
D5l8aLZu2GRNvwq19wYQlzSg4HcOUDRlZj15DvbECHgH/3LDqoexSda087cY4b/JowqZRayW26Rv
s01kkfnnrCZPjJIH0ATRy15Jdz2GQMplnOJ/0b33NUCnu99XhCYv07hjVaWaNem8/zziUqz1l38V
p/jYcTSVP7/Z3Bf55WITHI2CTFGK7IHNTyhsfgdvP7agi0tiw0h8EyTElecud7YJbAUorPLTH3Fo
XSUy3Zs9CD3OW5Ooza0zi3Z9B1+74RL+TVYPgzJYmoXq3GjESw+aIBXx5PeylHox9rDtkNb2xlmi
iZbkmQbOwU075YECJGs3h7OOo16dNjPc8QbJuccEIQBNFKi6ACbtOKtyuYZWfDzSq6ivvLmpZds/
tIEVl0pPrXGQk/rjnd6ky909bKKYY+AIRcwUaGd46OGtzCb66cRM3g4DtIosCAf9t8FBjmFBqrOP
ZoCh/n1DTZ1dPAiqvy6HYPco6rWmq14lXQb2DdVZtBgUoy5xN5zUfTJ/MJZwGhPobCzpJaJGOpvP
fCYLZAVYhF/PUGXmLD7AV2Ggj5dQ2s2o+rGSQBpQIgw/frAV01sDeq+sClVMRXP0dQRq1J7wLLfl
jfT6D8/wNIPcrz5g0vvZNajoANzl04XHb4T+fHc34H+9LtHaht75M2vJZkPxTD9rNOUCCd6AgWYZ
MSWkEftrJ9yiV8xmqpSJPC9k6BlrImO+WNYOT8eM7TkG4xyQ+KvUMDK2oGYLrhVTstbKQlUKUR7I
xzgxdhrWvZqN2HzJtqmJXCEaIz3WsoNYrfTleQiNC5AfEzCpa0jkk5dErefA3y0ibhvJqoSstHOX
wbhMcGIOX1qB/J0INRwwYogZSKBG9TBbdaVUlhSpMrFjN4QdoARhcaPYli6tOzW+knpzGv/dCx2R
4ITFmMb2hANq/wO/meMZ+w/+SuYjfqjNHBz0e0BPxrIieLVZslbys747uMs3ePjIRXBR8EBlINOI
F9DGszNwE7BGCbVQTHHRsBtyLpYZ21CJnGckocG+j+BjFZIk7qfpeChDoQEf920+rHSXWmrrTZte
0/uthesB+86SjGADwuAR594c3qVP+CpH3+ezsnZxkDgalqI+cRAFI3bgaOSV6sE0dawd4S2MgaPe
J1GKiemFiXrkqAflphmq/y28/cSg39K6tOyix5Yq725wmuaMuzvVpmtUFolOl1HPmq4Gl2kPm2Nw
HHoiA8JXNUkVoKCi6oksNxrDa46kdzam9O239Vi/CBV5c6/Y/ZUcRSoBk8j2YsxKfFx9AVE7utj3
pEAUuNCjn7vYQgRfkGieSZsxIyrxZPPi8SlIQjV4MdQ4csMwnBrwPIkX0M5n0wkDa4chXkTwIvDd
2wIkKTimk4ctBah4VhGFfavdIlFo3//NGD1INjoqDj4ZKeDG0YTCi0scSHUlkGr5NzwvdemtkoBu
+Xvrd58XLKvfQvzPEhQIvvvbKVWpYoW5z+bMyeF6pnL8DVRhOW6OQKEhSuNx/ua8gllv4lIxE8Vn
kZ6chPI8EL1LjyxWtDTr1kBBIVtih2AVdxbclk4L87zg4EowyJq/ztFwK0eKr83H6+jZJ7YURk0C
BokmBNrzXwfDk5w72CmRWobBXPPVdjzTO0ZcVXyamJDRWDOpvlqRgyeZEZ98Reirk1rNm3Bmghj2
F0Kzjp18scT9o4SUD2h25yXMT+ZshuNY9aGGm9BCintoLWqY6FrW3VCR3vlgggbz5ZFqZGm/fyKT
0r5p23pXOqN58AnKtq40QGRJF1Aa1LWD8jIU93s4TXK2mMsk/Kh4KSaj8Ff8MTeGbSlwZIcDaRa4
D4qbErrSrDYW4dQXdZAPybB0o7WM9m95cO5nAyMS1Z2fOzOqRqa8FWcji+Ilxc6zbUVphet4Vrge
Jdo/EFxqNKmBXXRAm1MpN3idcVOGpvcxq1d7wm9kt4KsfoxvoSEtZ2pz/3oId1JHmQ7rA8oyu1h8
4IkVKD6z8Y+Jnk6LQLYXKTS6Vlk+fLkIOb04VyVpq9BwR8gWXCgF+FIN3/DygrGhhFNUuZIXsyFl
1QVeuWheJR9zRwJg5Co3bWG0s18hQgDDtKMaTqgkDbiqt0epjNdiinXP374yMUaqAdiBD/y/VXRZ
o8k4EGxWgKoGaEAjZYlFelLeHo0s5Yl31S2vGkaxQOND+/9WoAzfMav1CjOs3XPgmbqfAR09oQsm
SqG92RQxlDBFRLE4bk8HtV2xrWDb6lOcp1kc+dGwEPk/kMyrmE/4ITNfV/rY2yCNoMe/copEAv/v
zjzlzhWAgrFO991xZUwhhxTzORJPKd5VqwPUHYaUQGnZLon/ZScfQMLTJH5c0ROY+oIljaHOCS65
Uasv2pG1Ffa0kk8f8kqL3NEmeH2OcyXbZk2fDta6jE4kp9gSPBdBM6sa9a8yAYFFlDx/olvaHx/8
CFXZkUUhnHCHrpnYblBbQ4kqzvs27V5zUANE9i0VSnjYh1w3yYsFRSK2bOQcMJ37ZcjMiJK3Rv8W
c6SAU4n23vLP6M8KxDSxLPk3pY89OKPlq2+uRQTjcJeXpNf8O1KPDfP/alTFdlK+3LR/MMI6knxD
Yvz1O8Oi4X4kFCFPtFZsC/Sb8L1fdxRfz7xvoezWdzgY1UxBEToYpQ6256vuoWzctHt8LDcDaGwN
a2/kzFFMJ4bQnPc+JCPDKEOqst3W2bdUpi1OdO1Yowx+0JOUc+JUF5YSxAD8P+8wRt4z0J0oZw/y
8O400nnOC7Y+thItun86cEnfTH2e1KKwrWfzWmTv+ZD0DrMutF7Wrcj+pkBd/gTT2/TvC/UITomp
7arhqJWIwlvreKTNz0tAVcrXA4QND4IhgjEFTk2foELJCN/SZz3twQR0LNq0rcSjVXpWoe0clKnG
rSZ2x6WgS0yvG2hO9Tr4TuCADrJBZ3BAZcZO7TS6muzpPSaorGS9hXbva5mVpjd9zqBAHIByVdPj
AHn37FQ7E3Z6yzRdAmcJGEsbuVlFa2iJtYQ9y9Fz2JUHWz71xOTbBN/atKsyBqbyjSRozNKROPxe
l2beIBhwd7K64l6uO0vEzn0fJPYpI5jgHOS7DLbSmvz9Wp7y7x6FmD87TsfzSWlXcek2n1y/86xI
jI/gb33s2urwV3CBoq+AQN4MUGvQtAlGJyGBOpTqAa9TEVswMDcI9OEtGVnc89QNM7V+pOxPPxb5
K05ENCGZGMB/1OYlaba8N0F6sTT2c8kYJ7JHQAnUy9f6fV6Zy4/r4ZSuxaSsiG1ygkdriMDfGsdX
L5BVgmH20PlX/X0s4hrpzbaMvkC8jfzC8436JWlFP2tjPJ4Ab7/xh6Ln4b0vqKhsguFdGr7yu6P3
zQKLewOfa+IQVEh3pXSYNlfDRPt6/bk5qpmc9V9cNhrmoHQ+CTmvfzTo0Py12edHsdBut5aF/cED
RtO/WOPaAMvzTlYNVg19SgDZS6a5Dx3Q1O2cbY8f1YJUeofTzrQqP83p3zZXUPVgJP0y5KShuT7x
kSsOLd7Esh8F/mwS5zLNRS7LpBc2xEjcJBi3FVSXCPDFwoofZYRLT+3PLX26XFg4YcmUwgqjp8Sb
cb1VXVwwYAM4CdSXIXPAApPTa/0Kjw+b29dLeaT4a5v7S2/5ZQzvJrGLiLhfI90NpceMP/gtLoK0
mxDUpMwrvaui/HdUWLOG4CLX4FGywQzt5LvsDuGglIv5ojKGfMv7RS3DIXpkjm2gicMpkNZ+lw3j
+tF/KBHhw4GXOLtW52gqGXMLHdXPUI4+ssbLJTsxCNc8ByXtTCo6zXRn2SNCufo0DLil5iYyobzK
nA8r5HixsSng32trI6yhCBBaIDu47lhX2ud55nH/3Qzul7mBDDP/OnlqEddGDTTdC3Od+oBAgTwl
sfbcF785nKefqlxglU+o1nxCFSi7U/8smHOnywomTODR/+GEv2FutFc8h1IuR1Xk1nwXyGbR/x94
0jUWkAtVrl5qj8/xh51FhSTXVOlCyXSuSfCKAOxHUrSX3U10+/gssSAabZLbOkk+5GwXYZKuPO4E
1/onNkaBcPVXcYsjVLFDXimiAA3aC/weflXvcQV/I6JouDL0sXemGCy1mGMh4U5vxB02ZnrNuTGM
m3DdhU0ldE6SoCUWzgJCdoDgBjuuQLNeyyYFt1dRDItNCmjyChAev7sHX2w3f9X2KCFrLAIe5yLM
4UDCqMPKilEgvYO8vM6QsfYFcjWQ3knCDbervOk16hM2IouM+NT2j+gNzXc869wycncpxRKTVr2E
cSwDz/n6VcR4hnof4wW8zdzeg60vaZHCDueKHuALCFO+WPirk7c3ha7M/nNojKzxx6GSUJFoEPWM
Kh1NXJsI+HZcShkSdM5au0bFzPim7pHVE02PfKqdzP/K70/WdJ6/RVTC91CKPe+SSYW0s9lPbWDa
zv01ID7NHWdO07IH8YDt6KTt1c9MQAAp5wj2DwhqklHzEwCIGs3XktbaUScL7yd11eJ9YX6iinsL
WQzA7FrRw0o/2+07s0DC7KS8LYWZiarWbHCoYqq139Rfg4GlxlJbLQq/i6PpqYpd8SaNN9rj6ljD
XMKxL4RIPUzMvql8n3la4nS0Xi+KOYn6XYQc8cSYb2MNG5AnZJlvd9udbe5dicTZVSAZ848+nylx
GS7JhX0V8efivgfUAzimNFHERlljUQt5HsmLIfvc0l+AbST4ERivPOg2HmXBETGxFf5qVTTp/7rE
i3B7iyQUMir8taqoJEXFnAmDcntabxM4UcIfdNN7dUEUkRi0ByGelrG5pkz+ZzeFZ1Am4HCyohJP
GWhLI2gnFbCTcFMoFjcxhF85BFjLPV2A1f4SpHTssP8kMzEM/Aq8GDaBlqZVFUjwqqUV/L79nCqy
S2WkUoAstM4gJOBJqpnIeVw0mPoWLzO7GJNBjmjkDz+fQngBxn/Fh/+TozwVT7bTSiKVUVlZGh5A
GrSXZ3I5q9JE7JEgEiLfOR2VUnO/ZuevI4OkjFwESOZ5i7qiNdj5+aIajzPt2H5qbV/FTDblfo6X
Zt9FzbpfMgMLzyoqpYGbBQ1eYf5OPnEsaQHJvAsGQ/LSMX0KdzNdBYTWuG62wrLuppizBZLOELRk
Ecp3MFnSNHI9bBCYEVXsv05lBSdDa1tG2mA367UPUjRRkwxyy5B6mcdWyOvgKHtp9aVihLwG8FCk
AhdROEpOXKl7PaSbQRHrJLTaiva8VCDO6AbDXod0Rv8mNzArd9SHChF9bIgI7IH8I3igk4TAZdoN
ynwUJ+XTArxtw4XyZdLz/BQhF7eFtadsNaJFBNkwoyzRpZfehiblXmxkmAvWlL+l7X8XehQT7VNP
yfVWgloW4hGHjFU6Wts/u/mEB03K5v9jyzao5eX7emt7KtPQMua9jDLOFhfgXXTWumxBmKnlcn1v
3xxEw6X9fOsCteVCXZ2+PBYJCC14+nC1ymw5Sk50KJx+X7aVA+5v1Nf3o8yG6V69eiz+Yi6O3QtI
Yc+l2WYCAZbi608a5dCxhcHwZqJ/mmZ5RsfDUq1vdu1o+/CSpQPkXZuo9A4wlJIrq7JyxxwmeX8L
FZm2gi3Gv6eyXhSNcooiszDgihRCy15MA3m6i7veyXHhNHwc9J+GHBIzVi8agM2lmo9OpXQSNTeu
aCMtXlsAveYakxCxQkjXlkX8s7YbXxori6QMFJWtqfD0Dy2hpEBiVpC10F6zmYgQao4YafkAfaJI
+LecSTpi38qZeu0sd28Gv9aT7umN9Ihp38N6jKwQs8bWtvTskr9R/XTNu4e5SAMMwK1T0y5yqIWT
MUwqsrajlZcm/md3LeWfbZf/u8tvslBbdnWco5Cf0mpq3NNNtKzZTFskjZ+e9olRhylDP6AGfu/A
LD0y9Th+2bHVZGrDYG0GG5f3ROc0A1HV4b1NEkvi46OJ7wDvGR5AorzD/PLklZMCYNYHv9IjpgVC
0HRYjEdr1BtRbLhZMK4h+/zKWEGb5g4Z7VZv5KY7cgczTHbtc5gWBIlkJ9i6bn5iDwaVEH0u+/7r
JXOk7i6GYEhHQCIq/jnesJtQS/rlpO+xhJ/YCZjZhXA6KRJJSNl/Ux2eyq8mNO8GiwWwOyUUYsAA
ixiywIeSJ4b7O6WRyTQYZZVlotueHOtaL1hUt3cWfws/sgbSeZBZ4/6qUrSKjKXlvY/xgnKtopvw
wieVRms3FHdLIOCCTkwR0G53vg8oCbVjIRZSy+8W/rl5i4qx//II2wF7/Ifj9kZuwH7hcWjo/OQ+
RqkqLAKREi+h+5WPrYTdRiuh8NasMgnJo1vCMEBjCcooTjn4tI243NFviqiV8aJxnCyMagXoq6LA
W08XM25F4ZWXfvJItYOMpyJrSP0GUjX5L+PO7rcenII4TxaByXg/hfQfbUsNiX+HboGwMOX5otcX
lZyE7ppzwkrILR7Tt3SHjVVLH79IUwhUNArbGAt6cFhWxUNtqyiAWUYSzedmthVTHV0KeyjWaRS4
BOmyKTAisZyx/lXd1oyBUTYG6eeguxy1dsthUY5vJUMd4iMI1aMhSoXM7cMPjj4Qgbegv7uQbeyq
itSJXStFzBfUdjWjJQ29EIKxr26DetbT8gATELvlb4QnAgPfSmxEEeR4UgPrhrwfsEZ0EzCYvN+D
W3ETkFYKxJnpwOM9gVfwUxQNb1S1S09i0LfWNyfh1jgHX36EbVIRMlzV04vvAdcsjQ318AZDdIJD
F5PwsPFy+0AB4dEVNp24aWt3G8/bBN9knQlSBQpPLpR22Vuk8rzz4mrBzQG4tqwYITynWLFjm152
wSI/zBOxM8bOz2lw0I9uanFDJJZwWT/Dm95o6uN9sc/0Dj9FPg3Seb5sy4L485KXuAgjoqghhoUX
oEyGNajn6tx8AutuWoxY9oo7Al9xbdSmH0x/sG8MRA77uDXrFINo9YOEBeZC2we9AblUmL5rYnmR
B/gYipxHEsrFv/XLS8nM3aoJj7UHTDJoh5viPMc9VqGeBEtO3HHKSzrqIv1Vz7w1dcsZyUyqetRz
ESt1EHDr/3NJATH7aYmxeVmLGAkw8/rJ6WFRYqG/fP6ryY3pMvNb5VDV4IbuBuqOmwqn/W6+S0Wa
eyLF9lbpN46hEB+3QZcOJ585NWAbyW0L0AwLnSA703E/ep9T9A+kPqg27l8kAIHh4fNrBMQrafPA
qXKpw414r5w8c+doRWEZtVa/vAkZzThfuVw5mHfhpEC7SxK4zMI+zis+tuaACihIr97ZNZYTqO/O
uCb1T8hzauf8VIBPAiDjTRYubfrvHrMi7ZDNT98Gxho8UrQoCXXa4Jru8iAHOdfuoXjKpd2OJzcu
N6zGqI2wpI3NRBYO1rS+/+T2sWzWvctRfugHwk0OvOksQhkvPnWVVN2qEv/yM4+c7jq0Fu50/Ewb
hIx6lIxoG6us4iO8OChCXBqPXXmW0Ln3nk3NpaJI05zhw1Wj/1OEgJWR6iN2KJ1kxD7VRkD/7bxk
QiuTN1a1/9o4hNTpPY+nVz99Q78QZ3AQMPaiwJEvVfEiExRH2gZsm8hF8SSH0en/xmxwLiLWko72
pfiaowe83ZY8wrBO4RazrJOsLfc1wnUzzBfOTsTl2Pi7lfjQhedw9how0IkTLnxwbAVW5CWJgLRx
FBSz8XqJ+ksG87eq4ATiVmU3g61nWxpI4l+kTu3N54bjB+kgcNNgfimZVGUToYbiFdqh6kA0A2rj
02wdVoHDwO6kVkcee8Jfmdos1eErFGq3cUdaz4b0WKS4cBUy6DT4BPZqYwlPm81JrSQ4L+oxFX61
/AjyZPEAlCLzLAmjGqD8qgEmkmZ4L2MQdqqvS6wVUXkNWm8Yha1+ooTokYHjZx8kU1EWA4ghaYRV
Nar//btsYakZm20qjdm4rtqbErKvkhFX7smXWFM+noYYi38+ZoVvHqLF6VstJ8J0RtTB9KUfAXbA
Zx290sZ9+b80RGaE58zsDfCEeJqOLJtK47o9obr2N/d4oChTfqc/vOsIL/3KFyiSxApCvifBGcjJ
gPvuarm4g7iRSSBqDmBjdoUcrH8p8vtUWbjfpNxb+/0dd9D6D2fQgryImfCBk5b4NSTYeR6ZTNIP
65c08rZIMa0ikSjXcHiKxlvkQJnCTxcGoNJMoP7h5nbyAU5oH73g0qfjs0ihpv697Cw6Th4iqND+
taks2pVlsU3p9cITsl9urUEZKHS5MjM3w90+egop8hgaIgT1Jv5EtVYMQKN6eLZinW1wprFDkMo4
ygybQiMaE0bw92lMPmp552s+wgcFE2tOY2Fcw9bgaiIResP+rnZNFkQpNn063rFPEZCVG5flps0M
sgGhXjOlfofPLf0gRlUGVW6wBpnK48epK7MUNcMOh09cdI1FdGisVIa8sRa5p+sC0TaFE8zXzwHK
oEQ8v1/BrFh1LTByUdKrzFfAo0JmRpi5y4D0cTgejBT+/h34y+s13umr0C6nOzfE92wJuPRaQnfQ
cVXmo/6X65gCBAT3iKkjsZh0kksto3jDVbrXFZaySC4hLQ7IXKno4Qae6w572Sd9u5H0Akgs39tW
s5AwdqvCOR0Q2nkh5iF1hriBPRqUf1zjncRYh/p8FRxEMDeD3O7Nr3GUFWBg/xFiNHUhRZq12VNr
VGfSsAWIY/JQSUinofayz6WK660MKo69gsp7LIUhcwnocHQ/+7jzApMvSE4Ds9C7jh3IefXbAh+/
MoTFn5tgL9REk1pswO0S6A9rqaqJOzHRtVEHwZQAcoxCE5gJa01u4Ror9x6De80fV2LymI8YDGBc
mmcEZdqKIm2PKHQwZ/5Tph558yT/j8VqJRVXAEFO04HUEt8bvgtTkrbPxQrIuuXoTr5uKW4cGMPH
vjnZrzwcqq9HRG5fxN23H/mkNSNJcgmWoDftyL1Y6krj2SxAe10HadyOwBQcmQH170w663kvWsD9
EtM/qv46EC+xsiBZQXBcHwV+g/IES0tGXV+BIsRyrr4J/cB/6zhZZeEp9r5B/41DUPshl5WoDabe
a5txyUa2fFs6qV2rX9UL1Zy/pc44xgB9yxY1EDXOK+IUFGKqIIb5RnhmQUBczA5aLhUks4eDV7HD
/9+Qaw3AmaXLTu6MgId47Kz8/WDIym5TTwLm4kLTcH+waMjxiohbVMSC4TY43D7GwtGBuyOTmFps
BfbMkixn4HmxctkABDLbiH6Ic8GMlH6FtBADxcDFoEhN16PSyO1o3ANIcsqoVi0d3Quq2RktAq32
jvplA5JuMxSKPX8dc3A97Nba04pRnFCc0QxpvW2/ozlXzVqYhQDiSCjQuHeQsWM0c8ZIZAl/JVcH
4/kJKIOzFGCXCTF/6CboiBA8DguoI3no0z6jTRha6+fV/NX06yiyuVG6FZt74ZPSlLf22KXwVXM+
sh5Pri8ECUsBhVsXgRJLnuy1e+4fxnU+hfSZOnFMcCRcFse8kTeGri99Pw/dKGsIc2uZpicJyxgc
DFMP/HyeWm95UuXDuV6tcFVh+bGtcRFVpCak9PBjx9ZnVpPrB6WfNsP5GNXsj9AzPyPQ+Cs8vZq7
cyD0JqxHYtHKD0ooV7fBlmXptv8ubSwGgw6gAPTYjE7pcKwHZobp1uuzaq9vagjgc1cEXFQAhdtG
Am84MejzMMvGWNOyWVAhCG0LjA08b9TC4TsdWNF2wgRUWEeY+hREW1B0ph7Ahp/Gus67Gj2NUMel
4pVTaSAh2zT+v9uiHpo2S2AXvoJMP8DfM366G3KQ595tIAz8WUWvJShP+FSIDlyzHlais8PtPkDv
n+6xUAUnuBFvudSLa608zP0SUEM0lgvsM95miAanUeCDc2V3op5V/OYmhq2veABeScNzWqzIo22D
jpCl9yZnxKSLFQAqzBFqlKyUrEgcGknOrmkKaL9k2G9F/DIr9UuCfUar8IMpSlRtQiO+0yIL5lMy
UL9tRZ4/5VMlpBfy0vqjoo9hW/PjiqL4kCwxK5Evi4YGb3it+QKLUVLXKO+qsRcsHK7DxrjKR3Ci
p0bfBz6yXM9W7+f0Wmro8vIIYNbuj0+XY5gPK4AX5m7sH9PdFSGA+yTuqouSD9wFcjU6dcPlfgMk
UYZaM8NzeIuNr1EZvgvGQAp8tALaOyZtk+TIGqQr4VqTymjpkRX/2q9w+skOKbPiOEvpDNgPNsD/
8ISNRv5GOzYOxEuueCtITQk2G6dv1tBobLwh3Qm77K6Es4CgQwf7jELc5Cp7qx7ApjOSNRN2CnjH
tB7urigy6xVwf1t2VatH1UGsivt8xp8+e21BFkurKKrKXyUDvIEUrC2hcmfch89CcoTHBO5xTv1i
snKUtsBiqvwwD+RJgaaKuqM4CmpXodmQoKpMpUTkUrHKrNI+xJa3esHE6z0pnhgwQgKSREF94Lef
DZVwjfBds7rLYWDLHlv8yzivD6t/aLDqRwXn2SKwO+OD2/I7rZ4eGsxQJYEC9sZsoeM1PQfJfPss
Nly3C35IvzKmi6zRDFMLIT/twLACDGVT4kD/ASlOplLarJTRq4jKEq9HzCu5h+cJmMhGsqMk8qhF
zbqcZGJEO7DwiTxKknDFkZWrnDce6t4Omn0dak6178twdQm06++F3sKBfzYjYCWoqk95K+rcSU4U
7OpjzkQaZXkoFxSOjG904j+FHGIWFO+wvnnaaRh69GHK54hWt4sZoi8CYMq4CUnxL48743VIgiaV
asdauaauLJMUkmbdbzI4T+VttzQhTr+63ja5TiBlxE9tR1Ka6a2FQIRkZ2lKma0X4W2PKNEU+eo+
fdOfz5yLxXSualdIQr3yBeVlbQhKfXliyrmriZ5LFtItmfPTM0d5XATX0CWB6cuOpTnkco4bd8jB
hfzIhONa2IEpB+KI//M6Fz3nTbTJEYstk4lw9SpQ8jUKgnpAvAWaiklsSikdDb+2J+Kx9fnEFHDd
T6hq6CjxH0+jfh3w7r1ybkr9/saE+Y7Jk/U37SHwBa1CvIIG9Ea+ZxUt/fKQIVLvMZXUDPgyhvq0
UuX/qb8dU6FOGI6dzl2QDqR0QKoHuY4olEsFc0GHQL6AJzCcevy/4KdgyLdXsBv5bB8xn1A5zEKx
6yDO50YkQFfXRf9e9+3Ly+7SA1kPmlgQG2FDTN9rH0qyLOM9NT/PpcbbNXLufzoavTPWrSGWLWLq
/nsAgqf1NXeXbmMM9pRSk8J/96hFlSxEBg4Rx0zDsZBEiOZYtt7RjeLvxUfmfTkrYyp4bKs3RnOW
BRJH6MwLaDwp9YqskNk/TS0hAG8I3f3if/SColJNeRnPH3YICJF/4MMA0DBv+L2sVVHv9tn3Ig77
/llJcxHIYOhPQ7h2FqBgclvabsFP1vEaJuVcbTtmgTA43voXPEi8/NYpFms63rteHs6qyBPO+YC0
Wt3IheBSETPpyDBMw6gh4qsoCkUn/zuiXz9nbUQLgBLYkzSjLLy47Sgx2U9RD+BJc4L+b66lWFq8
VfqOrbvfabn28NH69uEJ3+xF/ymAToOuXF8eHRoIahX75XdQJFeAIvOZR2NnW9ttDAYAW43QmmBv
xa5Z5eO0alHmgHOp8xUjOOhZEwVbBBYMDpRjroQADvoSfzqt/v3O5H8boLzn8g6aXlV0qUyId+VP
/SIBd05LOA+h+3+B8k8399vak6IGbbh1m4PcpiRqFX+FmdRqgCXBmjwEKb5/eVhkVDO62DjV/G8/
8uX/cyPylFAhVGnUKzY9r3FjsIdiq7kSajLFJqIGvvz5ZQ/hi6kdZDrM5S+0RfyzpeGIZvWMNaWM
sqIfFQHNyozg2JAVzeV+gBkiAifK3EOsfI3iuchyzcuIKSUdajpgH2M22Pumnfx0lbm6mrxS4Rvs
QQYjfiGb40fBt00EqygALDvK206clXaWqWlbNXVJx+/N/eL6PGnWRtY83ZtoslVVTjKfYZcVkT3q
eeEesOf4Gj8uAO/Vpm/rctmlpbSYt69yFSM/19LU5hNmMxSQqS1rvsMvzOD5qKSW7VW0AQXYLL+S
8bjm06LXoIDlISstZieRPNpp8tyLreR3LxAqvTaMS2t0ddVmtUsmcttV5f4pM40lPHFBGubpMZZA
C3mDCBTUrb/LIY5OoAmuTMF8RvQf26/R+beUktkn9SOPf3aFjv1fTFCfyF/xbI1Hh4NH7xGJF/J/
N+7Yaf5z0XzqtMPhist8C+GRkEw7BYqVoAQUPVlw2mfjxUhKe7ffdN1KDx4CwIl8hnxH+KbM+0DA
Dfq1MxjfhrxcXiCvj/x2E/kTsTyxPzhp5rRKfpQqxcuzGAJEjYSFOgvYHos4tV8vW0laEzfzM2VV
Fzb4+88xrb7GF0WV/7HS3mqBfTUl9yrKW9K0SCY6t//QtXN8jA6Nha7OijUV5lBtx9hKybmHQuRX
MI2g2NiHcXWCcfi2+Zxf1op/b7eKCtXa7mVZI4Gs+Nd5C84CM9/w2byR0PGF93tJUijBHFmvImUx
iu/A7b0aNcZFw1sKY5JNmFkgR67/neXXj9y2AJWXUHZ4H2Yq2xlaBDuTu7vl8scyPkJwabysc6Yg
dx/sql86kAKPfYB/VH1+hT+fqzfPI77Nz+5W43QiGJ2OtNVixwK9YsvGONUuEkVAND17OEhB6L6l
dc4iv7slaqzQ2/F9x7Qx5B6GAZa9gU+27KSI6mjmxDIPx9WZkJWVd24zkcWLjygizzFW70tu5lBs
tBaBy/6vMTHlKDuIZ5RIArK/DvEkFwut6Oeghw6YKbGR7agQ45cyOuPaqRYyI1qyklGXK8BOC96Z
EAYdJq5GHS0RcHgK8Sw34Kh6SK7wqGphMXqdQ1tKBOC+ELwdMKKiCmx8h9tUJLiNWqlrHJIUFdFx
dU/SmbjMu0jZRC95oTAcmkdQ0GZTUi7HHg/M5sy7LHwt9HDPBQhNVDsqkXt80TA4cBJjk3NISYcx
PAE3n1YY4BNQH9v+5YzwLANqz7HdS5JOCSwsB6nhjSzKKVKKOksFef1xaFl5ZSTAEXjGNma1K3u/
1zSCa/C4Efbh6+SBK4bAyGaNl/bgf+jdKLJf+u88guACiJk3xDPWVmYBpK2rThju29zpGEAmTSPe
fycr+37nXZibWTyixZi7Tuv1lw58Z7wXBV5blDzoHx9c9OC40x91PLJASUMNr1QIA7uUAujXnXdI
jQ2twdr0I/0/ps1zoCM7KqGjOzoJ+lo19Dh08lLEsbxJEivv4xZwf4i2g9kaOn+CzZOTTMEMWhax
MRDpQd5cY4WQd9no1xWfpzgnvAUmfn6ZxIsBwqiAokg+Hg3PRpYPIkrJGeJhq/hsfslXrV9PTOAA
nTMXOys7MlPW8xktdDl8lp6p12a3SQ+g0dp2rGS3x6oPZ8ktBryeo3xznj6kV1d+1zFkMdUOgC2V
3QOnblGmpFd/SeowRoGuta4+pGLQg0BHWorvpBpYtB9Lvi9DxtRAeflaREtAHHC8dVZ2g2+UQyDD
8gQZZ7l0/UgvpmVODnOxtOKL+jcyEarNsQDsVhWS/WKlrD6/HYHcrZNDEEhhR83d6vWKQRUfQMm3
/AoRx/Bho2LHxIXFwTyZ66ELgChLAZQnSQ7evD26rArLwv4XIQwcp65Ye7nHd3P6+rZ9Hnv8U06Z
WqT8SaLcoBUef7PfAggsgtTgQ4OXokRdoHLici/1QHD3kOneWvKRwgzXDDLn9cPSIeWKGl5DIFPF
6pyplImMaQdL2ck3u7zWfx9CLZ64cCTs1S4dSoJDvVZRmRnGghrl6bpozklGw8dXs/yGb7n1lyj1
jtaMrUoArMr9eleMBEzVhxHH5eDEIsThZbLORLS5mov0IQePDkQ6Za/8HYlR+bta39fXN6sFfRE8
bhPQB6bmtZ4Dc4kxDJvDtdD1WdPvNNf8Wm3S1ap4PZXSBLmw4uX7PQciXsciP4zhHu73Au1gi+kE
rrbrIvpnx6JsFOOvSdOYZn99VNWyaiZyU224XLpJbzFRWLw78fetQ2u+FGx2w2pr0ykvh8Sotr8s
DKLkEx/2Meyc0xD4lm8UH72/rI7sKt+h4Ees6qncl5WjMo6dOI7v/7OneYkK53jxhGHwRxhVzb8a
aEe929cQ0+PDAByKhXbpipF4NQPhOZhMWJTEYggMpUNqgxQqt2tOglqWBq5pBJIicZNiT9/GG+FY
dL6xrIER1DCIbbNyzpznHA7/LQ9NSRh4jUsWpM2zGFOz1GK8DLgm3mrkB5jDAx+357XGYZtm/JNj
t+O9ENEVK/CnaQxcavha4tn4Meax3x17NnjLoEvwIO3xSVGHGsbjRQXyxjNAqPxkWYS235VcVGBq
ur836BnseKQ/WTKNPMQ2nt8bxcWhzWUOO7Oxkssg8tq9vsXPtv1Lm9qGVvEZFGrcDtEUEQOK+NF4
fczKhFmcGiljIRkIeSnDCkJqywGl7caMIW9c48NkWH9BpfBHc18GUgKHKydJfBPqMGTcbQldhQVG
IVtIh4WzxJUz77r+XG5l9t9SgsIkSdCuEE7xkX6GzsuEYGq4zptSEvBsBiVHDI3XDvmaOoTuOjoY
MqZa7cvfAiw7MW53zmHzY4kifZuVp6SvKKEUBhrwoRYxrKvIFPrb/+zf7GqvKlMH/QVGz6HY06kp
m0VhDnofoV8n5WIX5q7XmfApOv+Zcg4Xisdjm/JP5J0vI2tv60qYSbEEBClA5bXjzzBAu5rhAMij
SdRbPYcJt+JdCDlS19bd7P/DY+KYjjOtiExA6kS0rj8S/4wWVczuR8bsvew0COgN9NlD8vS6aJ/i
OQD/rSIblybflYV793e70Pk3NSftJ85VuY+ZE7bGMdh9GgkIeatR397/iAyoPojeDDUQK7vkkASf
PDI7f/G/0AyGQoLhHQJ9LcOoDvvcEUO3AMPOhH5b/sA/Na0NWepHN5VbPJ9kECRKG71npr5aUZb0
GPKH+Cq7sdblY4W2i2FuLbQ5FVMYYbUI+zxbpgoPS3ByhD62ZXPYvstQ87px7mWUGpvFJDzBQIE4
WK5kfbOLea4GcOAVbNMzbSPqVn2+17LEDueLg9pCALJiSXgiNdopebGNsaE6u+vmwrDsiz78VeB1
YiDa+VOg6ZvQn+d0Iw7G566FbqAiUl4J4Gv3iwX6cHKrm74hVt3WRx4aXNld/AWyYuE6vs7Z42Z8
WJ5L2c205JL2sLyAmGJfHNRMHnr6G94v1elHkvyX4TUe41aeWIclwDTGkY2KfvjCvD7f1wiTtNKj
fNUX4ToU7+Qg3b42jAw/xtTQ3+SH6oqK/rJy/EiMckW/h+X9rMwA7rmCzT7dbA9p7cA1ACk1wqEw
KiB/gXwUUEpqu0kHIPB+sKgeZ0j/M7ltWcV6lOYz4lFx5k8LEwQ+xeV5b4urZZof3fa8qRP4jJhk
HIckxQuv5Z2FS1e5awSYZ9Oh27G54+0WOl6uY4BUygV1rue8T2DJVmPPjG/Enx9vOpc9RCKNuA/b
T/zOk2CsylgqteZN4JV3NOxqRZbWiottC7oIS1QWvaavWyJIFj053V6xTvuwi2ip1dSmyr+yvAOi
ma2Ug5F1ZUk2SpwZ600MBrw+sksgA0HF1Dt6bcixShZBWppfp07xGTmKB2t/jmnhj0a79qPhJys5
iPhb9pb6+ucW0fyN6u3gYGdxuVYZNvy4WXiJ+0uzpGbDnnP2a+rkfDlscDLLUSmtYkshFmVF5/TV
579bYgUsL8k31gMu1uqkGkbaWoR0euFYOcVIIQ/ASN0uTSpIAH0J2BlpOqGcMwQJaJzhu1ny+RkX
zQnxXpf+QbavcXf2kGTy6EUcIzf2L0cEKbZ+E1GCwxDWigoEdjARPIY15gna5ig+CuijDtGlVF3s
eWh1jN1FsJUkx3tpSlLYjh6m/B6pQZdQQokH0gvLZa7o6sqydrL4jVsUu5mmd7PyUHQFoO5rS6VO
u8rAvGTF6e13GYOuxeYpz6NUL4/ifzcx99mQbvliAIBaHPdtB/5ISqnDZ3sNR4zr2PAY+piaj0kc
jzX1+EZc8MBPfk3lWTVibRhhLTkK1gAJSMgLnS2uDAmbllyyolfiGllK62nAQYIYud8wTWtvkhgz
id0qKKcWmY1EZmnjs9IjkLxa7UCJhTI5px+a05+/7GZEMWjbosj1gGkACl5rYToXHMFXWLh3c3o3
iJCVvUUn66V9w2lxbCP2dV+KwUYOo736DetGZZ130WRhcVbT+f47Y3buAa++rPTm+kx5+9krW9Xd
kRhIlj3tpkVBTMP6Rg9+I6rIwb0HYkkEW/f6ALD4j4EfmGX4EeTsGVUjgUrkcFKSBuQfeGBd7AWR
u3KhSEnXmkC9kIdmHT/WmQel2O5LWHBlGCdZnZnsQHrXjnfdIuABxRS7kI5849PvK201RyNwttc7
QJoO6FoNcHX1ye8cJWBnheCGthQ0zUs2IaPoZCGPqrg9L8d1Gdn3w4wLeUcRA7AGmkfn9QtxziJ1
m5SJsZCaVK2VSfCViyTKjCA7UGAiUySjSBJAMlE3v5dqQ5Wq+iU9ZlxzowtgFcRfpCJFLuGHAy0C
OWymOMzIxP/qz8kes5dC/ba2JSvk3nBM7wXZkGLrAuOS0DWakMRUOU7rQRG10cy7+jhBo/8EKFkW
p44VQuyzppoI678QVl5m7kUFrJoso3PvzS0IhcgGlqwi+rj75cNlVsGJQmHBiHZHzDaB1GTFAYkv
4I9bOhwfdXr+LxupxQS9/AIWgJDEiBe6tyTzs9AHeVxyjF760VkxUpZ5rMDh3n+Zyvbdn/MuCnn5
bAFJ4CBVtkvIqGxbPRkftUAtQwbkNSPNj1LMe0Z1R5If6IJ9uOJkjmvRrhfRuGieZ6QmBOqvgry0
2UIN2Et9EflZQxnzTxVpfQMfwisbb7wrOAFkznb6WcPtF/ywXWEbYoRN6f6yrzMgHclWKe7Wdq+n
x0b7YT58RMLWHzGM0EsgkGprlNQe7R2OF5IH4FwpsLdbZVpys5rtbR19YdzjDlRJz+ls+7hPA3Xb
kGF7vfIa4MDiYVJFi7fq79VKK2wzuQQibmK625BSvEGUbbppmi/CjWPwO3xVyYDkWtavEyz6bfwN
ID/a0UGUUojmqvXF5W/hk/w0AscLwiV8cstMvVXja5i2r2VGnqK4LGJ7adf3C16adlV/I5Z2Ad9N
QTjFw/2pTLrX0YcL3MPeO03PZVM+84XMpsjMjDPd6EhYMp6YrkFeNeO/LvE0fUd8jUpa/oDXKku7
5kv9HG2w9NBg77g9b1M+3wFWTcP3/+G5dEwdAaAZmoIPtKA6LSq7XAz9L9LwPlelU0O9EhiBgeLa
Qr+byTvGjrEyTNCJh0nMf13+5BAD65FbNITSORmYjNYPMiSLgVn9HUU8B6wYluKTypOMB8YGsREP
lXzxl7ekk3iVh30u3PMv8+OiTDic5NYhMcj0IUACz/TjZUDuPUnbxJUb7WxkBw0AGcJmAxupqzzr
nWPWSQVlzdY4FJjnio2hbQqCOFCE4evCMJOOQtWHmU638p7Yqvo0LEFa95KkczNyY7HmI2i1XJ00
R6w4dJfUYmX1jrg8vbKpt8pZg9ys22qWqWTK1qj0neYslnQwnSYYLLCH8QHV2XQshXy2cPL2lrB1
L2TJbzuljM7TnXpX5Fn24YRU1JLZF2CnK9GlHlGIGUXjRVlnrSNWA/um2KtmeGJW19M2R/1PG+aG
g4+qqei9D0FglXFJhyh9rG9oYGctmANwPHovhZ2PNegqKD/ZpgZkIw3PBCC9vmgjf7nFpVxPaKzz
BITRxQyI942NNRIyxWPcdAsNmzpDC53dqOWYx4GOFryijE2gAv00xEwjgQovAsBgb1ewz945lBec
s263KsXjEK4s9mqcYUnKd7rP7uxSqvKhGR8LxikAdPP3EAII+RJcqUGLs9aopGgJlGGEarKQ+iqS
zUuvDAYyevSAKeptrsjkTHJerSXlZSacwzpKD4quqFDelFSaGRm3LwSKI4EI2XroKOlHSHd7Ma6l
dWoJ2NpzDaBkrzk/Q5ygMlSu4FRG64w9sVRoiYCXpR9kxhTuY8jRdG56jCwSofuWHD5/ekv+VJ8M
Xzq8e9AhW8v82XgcC3STCfrFcS4geLba49SlthjJRLNSRz017uallALLSm6Gnp5OhJfH8C/ag6LZ
rIVNFuH1l4LNI9MqYb84GnMJNipXiKJnWbYrQ12re+T6AZFhY9aimTnVEVWDa0Kr8r8+vP60nX4i
V4ntG1s/mMsoTw979UkMMYlXt4tPkJmRj0UAxatZZlwspydRH54LSoD47l2Uz6xqmMsFH59wX4dh
qKMijW5WDdLky3SoDAjQLQqwjm9xpmE/7zUOCUoZlQ3iMaFHzGTaq4gYZxVFXOc17B7MKh/yo5Fo
9HLlwwYMJPPVFbNFbWxQzJZBRYLpblkmU5ETcZYNyUFl3VWtMNjAY7uWlH/M/7cI6D+GyDQYxFXi
nB8bi5E6MXkLgOTrN0izVaUR1IHhM7XpH42waINrin3bijxv8DU+b8EjfxbFT7/of6LOYOvz9p+2
3XND+KymHZINXnBeKn3EPWuBaV7hs1vHgVYbCXzaMYW7d2Wo+coXssauTfU23kzay8fsielOO9co
ylaO2tAJJuZze0mxGFjfQHIpUxpjJ8tTvIU1oLC30u/pDIfQHv1Xnk1y2Uoc5lwE7pODc+jtuEFz
Tk6BrsGZPsbCgCHa4htW2dhJ8wo+Zk2Rx4/wtw+FFbRCOWWr4IbnopeGPaamj6o1RmNgraam2uE8
zcFqlck4MqfL98Gq27cgr7QocIcZ5vM7P5pqFvFC0Yyin96L6oe+3FllgJRFq/cL8IWdPcbgvf2u
ZfqAQ+jux5AD2UilG6WMt8up9vcWVlhbqMoD7XAtbAUWO4VZqInWYH69c5MiHJ171xnPs3P+IcK2
TrunsH1rjWRl8XxkXB/fkWbd8fYVPEWyRFop8ltwHTmeddID+nq4mD+REU1xlzPxtcUJnz3fya3T
1lYibzwumUw4kirBOx68LZQ/4ZpCdbwdYNXztt7qWrmnmXXw0CBP05SWcfyjbGrjXGC/0kuHGp3Q
LWhL5daX4g/t4FfhdunYwcqsHgJl0ZshRRuk3TFOdADieNfsBmp6M4YYwGstruGutVz8+T2LdTXj
hB+0QAsNyg+7mq3O1M0ZAnW2lnMbqc6FXSGhL1UwW+UwFrYzh2vzchfKRe0kTLXgMVUl16TB9QIn
8FJ2W7KqSVE3kt/sOPLDQqO0UnQmPhDZfdBi47OWe2d8F19nhgQfWtnM+cBt6n8a0rhFz3PDyunK
THH7aws/GySwMn9q8VlcimgeCIe9Ssn3+WmdPZTIcv0s/yUmGwDJODObER8ORskginbVGKIBvLBJ
inhOENye9bmoVdEzhPXqPB1SGrzq08H4HxqnXvUroWEwQpC9LFmZZcedJwwQRt1MAJLBMWBA+9uL
oqFBaoE+ksClnnFyGoPVvJ3n03M4WYRFwHo/DZQlV1hq1uE4L917tZm5GAXoyjACSNwqDXteYjsn
CiP6npdz/KpU0fra6L2akwwijlJqDdfYvwdvrvm7vX5o2+nOfHRoW6Y7iBe+XDL5optGs5JC32hU
saUH/uzx6TTe0NRMOb7Tz9ftU2gea00RDk8LsJv98c0pwY99CGDjrDOB/OOMIjVgB9KT6WYzjc47
C9zB/SfHTn+qjZopUWpmAkMCkBkt2UDFhLZGcQGkGDL78X+qc5ea/IFWl1xnofUohjeO+TakkQ+7
bYjShWzHHnk9z4U6MT3MOxyk877IcUqSsAleHZ4d3SzKfYM9xoSDnlq/B7Spbs+mJwjxhDIoXAf9
NK2W39Qs0+I3jvjpkkJW5QqflbDtlGdJC3i38x3uFSduXFJBfdsKDrK/8skFzeDuWLcqS5mG/8PV
1qj5Y4BsQ+sYj9wk5fLbLuGEIEkL7NPgbEN50EZ8BnzVcexG5Rh+f8j8hHBJO2D8+toEnhKzWz+8
YhZYHuAT78yzQtOCfdrBy/n98YhllQf4FWzdvsX7nt0MICCz/Z6py/+b0gSsWPYzMlrF4LRVubzX
ec6o4pQyr2sFRrIUSHyGt52DWDFlr4627OM9v3pmd16dWX+4+VK5dhfzfzxHYa2ICUBF1+rw59TD
HztVEAJpZ5bXBRFqI7KpgxW41oDKon70VZnfPnhejAZUzhQtZVeIt/qNUd+WPXAs+u6fgxjGdJRb
ChB7+WM5tFjpQ2yMbZ9p4LT32PoudEr/YiGy1gefAwJAw+OItaH8onkFHLsLijcuGcmjO0W109Ej
AQqKfUC+Bi11p2h9AtkpbX0peIMVHmzvDKQwxWgBVXrqMdprk2SRI/Ubz6rvWRejHvnxUy3E3NKQ
er3OtbQ+fGYvLZ2o8n44mGkLQP8d+iPYZ3eLQ0nqAvVfCVvRkbH5Sdm3cvYEI+vBEqRtrNXpoanB
vmvyQaS22q/ZP3DDdZxxzSva2UH7P1NvlVU26F3cTTkCDHvjR3hZxnlEPDrAuQ/bZaJ/MMvyetDa
YADCk9GlLv4NFqzHXUo5sTYRX+8vWQQ1zj+CpLbwXfkkJhRN2JtX/tPAkWIZHSsX+JAfRTgubE/L
k7yT07jW+lMdRXhMg0t+fAguVcQiLr6YMvH4WPWIiIsY2bS2uN/RkioOQCo075HaugjFjKzqHYpH
7m/MtFmhtgiDKSitMdOq1p3EW8vs6EPMVPwrLjGnHAyOOCiHdtjK0iHm5MYYKhuSr0wsEO4GiVTM
Zmg1/gNOKgoBVns4xol49TvgVAYLGAMB/L+3zSROLFDIW/a5NHUnOAy6Lfm7hJMPNkVJgGbUeb/O
LSZFJ27+wPCnn4LRkOZw8hDtkBk7OqECdixPXAQbO2hZgRHHQOc/6Scsca1cxR84YiG/p5KWv57O
uaFHDXelMaHYbL4VCKBhChPLSA56Sm8JWlk/kHiBRi0uG94OkMLZ3yIWKKBWrHOSKFnLOLDHRccO
gieY/m7gVN0wWZ2fgusktYO00KohvZzdbB+S/sKaT4yoRi1FgV7ItgsyuDPxTH2WNlpnKzivVsHs
N/g2s5C0mTaXwv8Pdi8ZOqqO+AVm5YgkWnNvJgV71KEZRa+cjruLRvoEVlqAQq73tUBphSPQja5a
I5rKSY7jNw2l5Ca7sSz5DDWysZOuoM2pGO4Em25bu9DsoFhdjQtLJh3uuSkfIEHsYgeFE1p6M9iT
WJ+nfYUVCnMq8BT44Uh/Kt396MtDQ34j948BAivbjSm+jUxiquN1lMJAuuANhrWLCCHK7vxDRB/2
aKtWx4ub8OKMXGsOE9oZgI8vZc+3fhvib8CFvENBwZWFx8tNL/m2ZA/MPz2+SbH3fz5b9uLDUwW/
ZJvMWU/2RHnW57fxSOcUYr6R/tWn94OdzPCTKwnK8Z6cjDFQFlSWoNKH+NXHlN/etVPDGpobgu7W
vCkbZD79Ez1wyrmtL8b/4gdO2SJKupHMOPKDuDPeJjkzlO6YVWC3ZfUvxxjzjLaSLXg86qAhcAQb
ugzCYzOdLx/M47eO6s36gSxTlZ0+vWYLNH9vYyRbY4jrnqzfnOyD8bwk6+mRoBzzFMXxN9yqjpCV
0Emsi6tbePY1F1WLgXsRMG85KNnctt3hba7HxiXQierkMD2MXFytj8aOyLttxEyyzSr+W9+rsmn/
De3CSZ7ZM9urhu8B+S0kBLNLfgEeFlGP3WaNT731MudmsQ392MtCCtTTFpILnYc8KTfgBZ9jpAfi
wvZf3Nf6c+pYDS65URXKDY8Hl+87GbNyMt2UxOk+vLhDj2gdD9fSimEwUS/OOGOdgD9ET16iPRxd
i6Clgxe2tDD+mU7oB6USYv79bYoCL+ous0xG3+q8S7FYhAh5BACleOuBfMQsjNOSJrIGVmaLsWoF
Dp/5a0hWe3O00+nOvzn0qbWhyZ//X0WSuX5lNhE2gKO9UPQ5wucXuPaEtMivsk8HkJLa9BY4yRq+
VyXknVrGHB9j+zkAL6qdkKR7U964yKHO+Vn6zRH2qw8gPnpImPmfJFW5ilCXAkkMupcM4IzhDZ3+
JVEijI3c14CO/gWN5N5wDM4ijpA5FwLeuv5hc5wYkRNXYN4imqONa9gP26xKQ0avMFNtntlArxPT
VoLJ3GyAx6yU5czKb+5OPM20QsMrkNL+8nkq+kSUEux/h7nSNdbid55q29opJqQip5ZS/RsNo/Sq
nrmFPbdeXTGBFMX/KWa4JfqaVvNSsGwVZBTszj66J2E8lOJVaBoz1CzyHtGimWzZ3TH8GIV02meE
MhKsGKFbi9yHBq2f3srjrM3qBa03qk4PmVuXJZdmO0ecq8G0K+R41VU7SB5boL4asp10KDSwcym7
bwGr+txr719cyp25dmWd55t0IBwp8Fz3TZZs9swJORggtQG8Ouquq+9CXcZPQAmiakO9eOlhWQZZ
rLZ90QHH/kSNZobnVh+Tgo5wNjHzbm7EkKWsomMTCf2150SDyw9xdCj7VqIV8NSHcOd7twXx08fY
mBAYL1yGHJNdebbeZ52us3SSK32THhLzBBoyHN+xYjmTmYmzejf63vIGePNvltftadta8mTtHABb
HZqazOyoZRaqQ7dKnc+c1eEa8iUlY9WeTiFAStHBLCTQRFcoSz5jjiNDYmnlK0+Zr1lzmn3A1dLA
cV63bwCSE8vkuWe52Utok1BTw88tV4no1QMMeD5Sq3JdBNzjqU2BUeZVT9Pibdhd1PisFhEGFqRu
NkfT+55WFSbSQ6pZiND13DR9v2cU5xZr9B68QvyzIuHERsAj9z0pSxkvhELQdzXMU9bwVD5CFiat
hvNM4kmNkduH7od+toBIxHQc7s6YjnKiBR58J8JGD360arR/W2LHfbjlOMg3BzFbaNNwB6zMvDd0
cwHv1iTrTPmwTbMmsMVrEqnGUxLULCSKqXLcYkn3yqv5rEXhw2eF4YPHNAZVyuEj+FpQ89Krjmky
0aAnIOmh3li3C0cME46s4OTKQ/FW6FncPMl7/81g0hpHvs+80KE186P6yAVCtTq3+LU66rcGluOx
lHlYAf7IFF+klRaTe74ob2H21Gs4WVJJMXOE90uvXqfzaaBE45d7JalIdtdZGO/i8K6yrmMpi2Gj
EuEYrbaP6JoDYEcX2br2+/3HIXsJ//3kOtlJXNXAZa1+jIT71rUJ7i454YxlKRDdSb/inJP4WLni
cIu4WTcjCK+5HlxC00dbWUFuVkmWMJoW3nA/KZo4kom11ZnJxOFCJ1K5xZk8OsrCs7lvfmD4GhiS
Ka7BHdn6VTl+p5wW5HX0YNi0LGAwuJytB5NqAy+JcTuFhk28OzLt2ToCj5druFXRgv2PhThF33hZ
cIL7SoOwTgKJBzIk8QEKvops6k2vFHxgL0kvVNm4nKCIRNTNvM36JmdahryuHrnTz4KdqSfpP0yG
/EH/kh/s9ZbppnqVrSVv4Ho+o0VcGdW1m0cEVI3ghg/+NwEjbkSZuU6GkSnNqK1261AZpqpcd0OX
YJlN0rEyhlHUsIHAqXxA2CKcym8qmis9/ijiG6Ds+BuBgjmX/YdhjStcsHkJmZLiqWzEe/OByM/C
s+vBOOrmtH76sSJkdTiRiYVwjruGILswuCZ6Q/4Z1I8vihNAtPPB7shwJTbdtltA2iZLrlqXd86L
6ZwGXSVgaF05K+AnTyuvmaVm+nhyvBdX4Y/MMJ9FS9hZ/WcgGoArcEf3pPCSAD1VKZTVAZE6PW9R
ZzBr4iU3i8l3xoRevlCErVW4azCJc9zzBl5iT6tusIoGCbt0q8gcZZW7KrneeH6ztgl+7bARWmWN
4WeY5qQc+EW1nXX/3XIzr3N0WiKuogPVJ5uHOqT/xVy3N8qCXeL37pKEg5Kae4K9gmpl4SnF4AH7
d40NMAmeINmN0/8vgaT+6XvXc82QUlx8zwmovlu11XlrCvmuUZU1JBmOcxbWdP/DQp7U7DAOdRTh
++T5gkIhYH2hb94vCZqGMaqRianekmb+AigzOc+SMv2/WkeZ9myraOTIGkxKZ3nRauOr6qIUW+b/
NwTNJ31tmEAsqGnbpdQp8V7DbTsqpHFxfbIQi+ZNV8l/u7JwuIf50zHLd4eHFsMFWKK9iLEMAqz5
C7O1sZeu9rhZNo+oH8o3eFCY++jXhTyFhWF735rMV81XlzG7vfbCjffI+YsFODWvrBOenff6NwQG
/sD1oCsXhYnRZJDoBs0JZDlnxZ2wXHye1EGWZ3kt+thl1MnaiXxx1vwyYvqqaJDcZ6NgJIH62FCc
MDc9b4nfL0GPVGXPedmN8YP5xeQYL27gnb10BVyH5Dng91OQgv3QzyzE8IeoRzemoXS6tipam4UB
cL7weyM01nCjPWSZjI2Rtu6u2I2k5WomHARscPzHGlj5PkilXSG/1pri2RpUtMSyKMGy1Y3kX7rN
2zn4FDtQiP8Gh7EULDhwMRM9oSVt0Ne2rTWyhylazpmmFeJNgkxjUJMZBuZuqVxcOZuSZ89DVHTl
HUshwHAbmVo/+lw0qQVHczb9XLSwKZ1O2fRRY4e19doLRI0BGnsLt17Tc0Nxgipz+qorJ9HNsJFN
Vy3lHRraibyVqs78Rj+uJLOCykJZDRZlu/jA6oxpJyKlevP6F4slAE2TXFVAZG3CHvfGDyWmzxPs
zW4MBfu5di+Dk5PfJlnMDk97rdVkznKFGhEuLpc1vtbPMaVqhk/rfK/AQ8FPr3FaqiSkYtCB4Pm6
/Y6ISwj17ccpnUANuN+UDFV+yVDTc63w4I7bpNrhcjq1NZnUmWyPRdxpH05YhU1OmniTM95K6ybE
Uds9iT2fswZc0TRj6mMA6qUhogSbxHJt2IL5/fSJI6m59PKO+muW6YCGYm9g65to6+nB/URAbSyW
xEf3dHdxs6i0fNYTgEDs18gI00BHPclT0KNSi6aeMBZymDaDF4SyXd7P7AWyWGw6Pr6mvp1EMlnO
o/PxcWDDfC9tNsVdWuqShCryI6tyo58zpTvoFut6zvvTjdU4H08PV5zPj8ntpRrDzs3t2e19AXGK
34uAJnBjkCzElUtRoSFbowXAXiL2ine30AgUwi5Wj/SyEELPCHv1lgljLlV77Uyt/Qn34jZ74AkC
UUrycp6JIsS5XTsXO3GHbaENzu/8lhf6S4MklH7HcIMKQEtE9QjjGuvqFQeZIinckqoR2unWkFj9
BOmE5R8NqOrtbfVSMyZmXR/Zs+JC05kcE5C142vK9kNjR6dTNPMxxuWKUisqyLxUFPVlH5JDErLF
XxDfC7gwavzTaNKIzu7lXJnSwEBXUR46Q+q65Mxxkh5hsUgxCvFxI+2ANCNsqhioKXGPBGzZw+xI
for/5/tQ3nBUTY8uIg2LUCDMFeOxDBKznW1cs9r3e6aYxCN7u8WUkM+2+03M5jE3IpaZe/4HzdH0
aicRUMT9Ltf5Tt4KmgWCnRNqmuKql4qOmhVOXFPFVkDqGbT/ev58tPfbNml7VIbKMDGpyh3JDt2x
RlNTsXQ8aeW3Ya1VAgs0qurobW/+pPDF8De0rRYFxahwiDLTqGXfyeCs5pDvTY6UUVdYHRxS9PC9
2W6Ce/ARRBBXdfkV8LQ8kX9CtN1yG12yX3dboL2yy54yMZTyFgBwTOASlgz9z6B+Y/6+heNEX1iM
ngUxmMFmWblAvFDPOSc9nTCTyjuuC04aJ2Ecl05uC2VIG0234dz5xYjcvTzyMTZ8G4+FrIJ/lq/+
RJQOwDA5q8Yp68+ITVT4H91xI7sEvXR81mlqn7gI4OH5FKpBF72XcoGrR3agkv1iEQHkRmnotNfD
eI5JDoR1MdkgHEVDx3gokmoAG1RG0a80dGdHaNpyvGt4VqH3eBdmhC+T7CrCvhMB1oiMW4VjLBhF
6HueKy2pHXZZjdk8GqZ54LOE0QMqjeAhDTUgBkfcbpfjTG4t0TdS6EncAy4giAA8LoYPasFeEHed
saGG5gqwgl5bOo5u4xag3Tv8sTN/2POFNStIllCk5GAO0CU20J8rMBMT4pmZBHTUwCSTNeAJJXCY
zy3bleHL6B64dPUiv9o9/fTlajMyeu+OLm3QQVRrUilTtScmjUfUipXSiFTZUj3721zk0w2qlTQq
K4p4dPITIOPUzfkrm8UFMIREiv7StbYunv+bf38I0ZwX1O8P3cP6KTkANNJmEo4A29BcjjcV+pWJ
m1bEXtj5ZdPeFSM3kAn0PMahXLPMX8nouapia7XlUSd3cCl5w+7CY7OjsSO2o1wwRMPg8CAUaaUQ
Gb/WqbF8StFS3nmdzZflQZZRfXYIStGzRvx0hQhnsHTbkbsUUJla8kEndIcJ3faD3ovp1/eg1nmj
ALh9aVqcXJbbFXBHZglWbrF1aj/SLEsn6MLN5NahYEFsKk9i6bnVuiBKso9yUpQ+yEq9qf0WdyMV
/uTVm5fZHCObcC+EKN5c9ZQVZOYVgXxZqEluj8UMz2VYNOXXcVZM0nl3xFSNmhkZzJDlIOsn5yEX
ovOA7PAmL1YhGvervgalCDBaoUm1wj4UubpiLwcQjbi+AtAINnjeWsSzC3ykURsO0bE+FkMaIhNQ
VdPh7hukyiFF313fwbBXc7BRnXYS0YfVLvrqxfPuHTEe8zbgB9+czN91H5spQKxELqh7dm0ZdDpr
tvPAU5mVWt/egcRsZSkl+31pGpV/O0K20NnQ02IqED/fs3iojzsSbhPxCFxp2JJzsZL4WnwSSV9P
EbECON+xQhAILT2aixJfnw6sNk2u/og3R6in93K5gB6RoU0p2EYJj9dXlo2zdYUGLiW/2ozq69Jq
OrLw0JoOG1x39ewkjXODRwBMDMmiwRQEMqX9I6lBqZKZ6mve2xQ8qiG41I0rLKwEMxHClx4yItS0
lOGhAFuD/+kUZBrTE+ZCRtzfzCUKTXq1Iz8/j37mtSZAYwc+4sJ1TEKpIpBOdYKYgEeQiNPXZ21a
fclDJZq51WD/aDdmO65EVbNCON56/5uO8VPAnDUhHQpQgB6rJ+oOTvpaDcJJbphHcljBb3W8UTjI
dOrIPTb0GIA09hdNp+xenTB+cJ1UsH1jIOdjwvn8f3226j/dbYNG0B9raCp1953wZsRpZWZR0ctm
M4cYLflp5yN9ZvG8j0bpBlWu8SY07hmy9Ud2Xg/5r0uOdj+a8E0o4jDa+NrijXjg856W50NJFb6E
/IpuAyYS1ECWS+cwsq17AuMOg/1zkns1VqahZXh1KQIZB8TltQoDPxygoOVz02GYMIH6S0SWmMWv
tpva98WpxYBPjPacsAWV7cyaGYyo7Q6JWl6G4hvWYPpJ9k51UnOET8uBoOZGXXGpI7yMBy6qhRPM
2lAoEQIuS3OD3DzaNuMFryZtplhkgQc2cI50dOZjUWfzZI0w1/LYkW9x1cngQVkdPthIi/FqWPaq
EAsnbUHNsp2OeCFJgI/OzXlId4FxEQeepCm0PIyPQtMNKSO88SCiUX0mjsC1zEZ0+idF435avClE
0Sa0F+IL9KrvDopczEJRyASb+Rp1UY/bW3O6sz1FTIxVBMPJlgJtc2vbRUZayf0gawf+hwzcGX4g
FhewBnnAh6V7OeVn+vSKQHFDRJGOS2n9t8ihZpkoSAodJyT0Nj4jimRFBZbtxZBxSo97NciCQ4Z/
0odJvMkB4ICSRhSSEdKqeE5zLNw32ZdFckMLFhjnnaZGbcWUmsgtAvxz3JCHo1CA0cqOJxF/4bRs
IF/MhIWsUBtvWHmBWpFmqlkxSXpL7BSL+Rw6w/iDGjoYtQb52GYPZFkpD8PC305efJxorgOrw+s9
OmMAFHgWLju06WhtLDAjMqlWp0h7sdIgPgiMQaEE6hPoDeUKg0g3CVSUMIP116vNgc6iQmZgkaIF
yRlsN0NbGU1XneBn/h3hgjTKIvxLA+IK/z6G4q+0Z+j65p7fVc49+bLOw/1thmfjhNqxHeH4pKJn
UdTSYgJXrCzorD3l/1uF1AacpPd1/jY+TrW5/ZtYroIw9+9WD5YDPgaALm1jCXvgiOmtUaoAPdY+
+HNJd3WndOS2nfh00+8JitNaHTzB7yVGOtUxU4MX3KLpxNYLtDn7r21aJ4fASb49/k3bI/A9GZ/d
P5f/Kl0588bDSpWwUsoctLPrY52A/jAA+s1Z/nl4OPvDCdSIRnbc28z3LMDCmXdLQ/uyE2+52dk+
MZ0l0imet9FExBtH1JBgMyNhyD8QHNty43Sv0r5fq81Msc4RyAsrB4DDbJn5rRKO90dDlkyhl8mt
6jsaJijlZ8kLqVKAfpJlqOSVS1bguvqpzWo6iO76TJBexBh6O+74dAs4zp4EnKqKN7wTbBklSg8i
gf+1ltnlAkhZii+qmqCpGXePJb2FdyixmnE76AZa/2sVmVRrwwJK3P7UsJkmN/WIngnRumX1tqOk
mGeLeMmSDayUMBVItL4CdvhIoDq4w+XhjSd2DUfmn+s3+icARLCvUztTsdtXjnCaocXEM88cP9gp
mPKw8UXit8NkJWxvAN0yPF4L5JO3jhlLfb+au2oZJZbdYVVXSsU9p572MsaZmWfZlJGWNrci0Mi1
MQgxlFkqxsoVX9N9C4w9ggwihqtao4YhUi6aetmPNJaFhDpPF2vUO+9dnXGCdWzoo0eCQgiLWgw3
1izpslxPPBAlzbbGqIhu4WDl+++Zl3w8+Wtfl+l/jYX4KD8NkqWiMa2N/2R1V2ZlPuWdg+/8YHJr
je0JAvvPochSh7iyifZ9ldKfPE1vw9gRf6c8GkFlD6ruJxQOsJnw1oghXG9MfHa+codUUCa6jk1R
WryLpJu5SalReEkkjH1Fc6OTMVRuMLbqFA8jg/GC/kdWVLE5l2vDy2J7nblZK4r5tc9kaE+ko4E3
gtqAjS7zCAezq3XmK8lXkGC1xakaFV8JV3OcVl7KGcg6dmPGGP98j7HpXd49wUM6EbPxOgp4zXcv
nJAfK6S4Fhks7VxGwklv19e9UGdqhjZUdekWtZk1luzSqSRwHeAzl7DxcaRYBgBccU0YEf0eXFTV
SjA5uM7C6x/94yIJnLeY8U84TV/RMlq5DH3/FiAU6e4XeABy8/NcnEu17+DFGzoWpc8LUinRg3Oc
KdBsDMe/M2STCYkblTCCPefAHzk7vqIcQ1J6D/6Zk8kQHp22phsH6cA242kruvJ2piS3xC66I+WD
VXtqbk1RRJ9IpNRhNjQBihQe5Duu0DqxOJr07oJnZ8LPgOo/jY5hl8wbuK0QyxQmDbfD3NJDp07K
TAvSfRbFlBW/G3iqxdm1eexo5yNQXCANW0kz+GAOQYcosjlxCA7I0OK8btwbO8y8N9ZUs8vPvCQb
255qR91UCPW7i39Qq1og3pm5yHGUpdJPANCsxYLzskcROPMQ8x/qb68zBIJGI3p6mQaRXC7dsf+u
us00q1+f7rZytbh1k+/jjuV+23RZWlvU4UJ2Qk2+NsfQsMxIbBlkLziN1Z7niDZEsK92DT2C6rfK
2Ry8TgOM54ccpXRj7MIl0gtmJjdApsrehdPI1D6zUgewgmLuzk9RwoEtwV19+fffcMfG3lx87XDC
HM7N37DUgOnf+QtQMgxS5l4DZsivDOqpTT5DaoRX36gUDtWUgokULEXaAoSuVaC7QUrCa5zjEk4C
FH0MQVeTf0/6x9e2WrFEhSxrC9gxP72VUssj2+WeJ3v5yYfqvxKtSDiv1qLVS8R+K0R0xUsSzKDe
GhAZuTCRqsRA5yrDiui8ZTpBDkkFviWxHSVq4hk9NMxsLAFj8g70twiXwhKM760x55cp/fwB94T8
rqEaCED79PU5TVvspptuFqQbiubkV+o/CQ1lygDPtx7hUEpRmkwAVHVDafBzMT++wceAnJgV3LvM
hSX9fo6gpmWEVlDy0q3i7Khc3Rs/OtP8mQ8xmqx7kYCJXlf6sQi38c3IQHJwlvPxER+kf4iNGP1T
h5oSbcT5QRR7PNK5qmYxiyOx7JKHBwP06uLLx/m+M2fUD4HugvAvyBIdUbeOzD0O6rq+XsRu/lu8
QHFOy12oU+jspf8Rwj9VMmzevDCGnws4uW3ZNAn9vjUxsF7F1pZalOG5DCJ2Z4bxmqbmaRqnyR0b
13p9W1VizVxQZWE94pITiV3gP+vpapV9m1pnD35YXRGwXuF19tlGcn9xksVToLiDvHyXflS1rT1E
HrIcCu/PgG/An4V9v0SP9u9k/iCYczbHk9FirtUx/wHHSVZoPom1xkpcKKN8s9wL7EMZilG8uEmP
KpPi46s/7cZC97Zg0QI0NhIm0fW8fUGECK6WGAw6X4Kz0N9QyD/fYru/A+TJG3WXxy5Wtobd+7rD
hOmwf938BeDcpGOl3/xLVcthOHiTfNOQyt0j0m1k1Vu3Mh4vLqOzYgxl4CDxdFTcSyl9/0G/IV99
pGfa5R4Sz0R84HUpLa/YskCjpnwLJTxUcaPbDIFyTx3pfqawj+8M4Xwbn3asbwCCFM/dTgNKOHtW
/c1/hgZBWO0lPNFu4mbwoCiIceMInKa2GQJsMg4n3BeHCLjcjW9+GS1tu+ndPcinfGz0uxWiH3J2
M8Mgou6E9lqYjBKkxwKVAWYV91yQge3SkPDvjJMgzktYUiu6+mFEQnTKkEp/3/oLhFqxokplhy6/
cZ0A6RmAt0osaXuT11wgpSrHLjKm+LBhdE59Z0jbyGgWd8mRywXQ0d9TKNfWwO1ldIjGeLJBV1Z2
OEYiyIUhB/iAF7mknVB/ljufsQVgKOpZRrYwHL3D9p+y5iu6fq4dZOOoGCbRuEL0i9yoouzMD/MV
85LUP1R8HAUloduZDCB6fvSxwB9ZetLJvH4UZqO6nM3BhxxJE65OdPEOHgyd5Cm+Wt5bBzZ+TqZV
UlP33FsAaN/NlYA15RJ4DGoTWLwJpKY3AIaurLHwLMYzgZehhDyExewO/rsw4eRmIw8iWrUjDEWw
aW+n2/mLjH3Ya0szNyb7bah41IumFdEBwo7lICc/sWxRwg0OZgIopPSGMfv6+4Zp/W/mRlTjpO3W
yBGLUdrpMAkT/WFma5lbomXbKQzlrSqr9X/bWUuWtxs5RHhgD9HU+AOUhMZhUSrxZCIseWcewdbz
bvHlUfAAzCyM7UO/OPrlmPvvEqvnSF0eERZ9rW3PgXEq/aVjniuNOvtnTQZXFP/bboSGBsb0CnHe
aw8jItqCt9IkP9SrRenDpvmQOj37CKtK30nOyMw3zzzL81kEORZcEUIrb+Nb8QJ6rEhIt9o8aCCh
j4FwoENzJqvpJxifiZFySqjR4LzlKWLdjZh+7EZPev0O6c74rTd81lRuP7nWktHs1BNhs2ttAhNq
t5U/jN+TwycrP82+40b9nJzmi9NlmVBFZ+GWZ357GB1o3x16slsFWZTqQb0VR1nxSR8kwv/j09DN
pFgLW8Q/Y4/H2NdWLTIFh30GsnqtjkF+K4cjkHqrW6Pt8yp4jXGwNwLBFNPlVihZ2zLy8UVHW+BO
SM/4u1msdGyhZ9XO25QJZMOd2TEULMPo3PvhRMvHD2u8YlRzkSCyq87RNbxTomDbLqryWZrxq4XM
9sV66w2/+f6IKvoOzifx3AS2RKZyRVq9vA5PFycPsbmioj7tL7lBtHUfnSqRmzY/wT9EOmoBeeSN
E8tJkKdjltAbGP40DuQeKOYxv02I4XO4QTtJahfyIjsu3Gs413v3gb4m5Ryy/wb+XbhY/UHCsN4a
T/l5F3mnoYm34M0SpMNWdruNkVHVpy7bporrFUMnpWMIcGI+skUjnhloNm7XQVhoe0g+Rsx4h1XU
PzILtGKT+mw0kS6qH+Nu6YldsPLhsm/+9/PCYxEyuAwUWl++YvrzFmOMO4ZYriLzmNiKab5kCq1D
7apBhcjD4QWNTGTtvCYoEDk+G1NhN/6gHHvF4e5ynaRcWVnO+L726azE32ODQHuYCIsW7a6Wf8RP
LEaa5REv3twl7y/UXZtKVpDOLqP7C6EOm5Qwy7aMdZzb8pBNd+4H5fonIC4Qsx10oJR4CkqOj+pL
zRMhLeCloFmygMUKaw31rZPuICEvTz1K+ezrYbDxK/zQ+KnDWHsx2LA0OtEQbIyOP+Is8AopUC1w
R+VkRnd7wHJYu6yn14R9aKr437LSzPa/ygPxHMtdrOkAKukU8jwK60jkJ9WTDnO59XlU69WFPRi8
YIqccwDDsR99npgwoCdB9uIDMTH7BEAcbyDgYZFah15TETzzdtlKyUfzTNcDjP1BNCjaSxJxPaxG
vusr44TZfw6xr8NjwXhoZ38gG2pz3T8f1nnvCtAxy/UHPJemUJH+zMU5xbw02ixGfRSHuT7adBK8
/eYmkIyCDuivP4PgU4kN7pVxGvLIhAeKVoCvIV8ERPRq02hRMYC658nwiSapjuVVeHnhUrd9c5KW
yX9EhRP6+xqIJnv0dvmyymi0rhKDUsL/inmVSVnyN8zncDfH/NMVMeZo1aAjYMjd3eKqKK0sG8Ou
aZaw8UszeGX3guW/VX9JaEocZtMO1yq5e56WCGDiDhOZQk6pATvyAybYQ0kPJyGsRcj0VDPwvT6N
VrryJt7UsNq9+ObEgIW94rVtFJRqcTKvry8MNplkHh1zKygJUJUCCYvmbd7yLUOkrKyfVOFwKi/n
k5RIGkTGv3yYrn1wS/oNRpIh0+2WtZC5f41IXJwi4KPfMnMGsj7C7i2QMWIOVX+2AUifb9y/j8+4
GppICRhZggV6yappgyVL4INNpfkWyr9Ytx+snJhjYDxFd5ZLFhihGYkwxRyvc9hvPB/tq+pXaUeA
AH8Fc1WZYOfxBo1oQ0E123VJrah7mZzEXGihHwnmnxy4lPLGpg+NtK2gYFY4m439ezGNJr3DOXUI
ZNUW2zsCUSNta7iGVzr8RvpnNbKF7Fted5C5CCCxw6ICXQ/NAwCy4M5A9jNFtHNpQnxgJv9gwrn3
Ltx2fRky/2SaT1qqjVWfWz/DLhI8aDqf/TdAF3yUi9AIw0MG2RWRMQ9OWbUFY1R8JLjxL6DzxRJt
v2lKxJiTob9mL0VxrdGcmN+siUH3oB62eNkj08bIhBkeuY+FGIj4vb1++uFh3TKa6DgPlV/57g8o
MI2bDrV2Zney66YO6gXlGA4Xe6t4bKkQK1hllHFKcQuVF8RG4yGmLJMZKQn/0jobs2x6u9kRCb+e
UNAszNOJRTsLZZWFZEK1hqghjoJyL5hMNmAYwREjysK+98OIZ+apJCB+acGYbJIGbv+jxJQq3659
Wo93b1AiBBbDq1vkO11/92hOAvGC2QaZiUytER1CZ7pgks1UWKY6qBXQzR12nwaootQRlD4ZTjSq
Knc2H6eFniVt4eJ4TJ9h4dMHvhXkRz1/+2V9T/y3i17M6+R6ADKW/7F/Z5f4VjXkgh1tfXqOulrc
gykln/cDd8VtYSLFtULy44sZP6JgMHLJz8PzJpU734MoHWXG3usg/XluFpsFowmheIG5uQyiSpzl
K61oalE33YwsV408kTSfr2FdU0zvW9dwodR77f4aj1lEFY6/HxoxKUajS/UxxVFURe5OD7lZ2N4O
9tj6zuhoMCob/5L+jfAtvwq6jrlpagTGyC5tzxeOV9TbwsW1EpPcx+CUKxt0wUR25ipAYj7DSqIY
bG6BfS/Hi+V94awfF42S2A4MlhDswPGPPV/yVgk4Zxi/x2Rd5VBFEcjWdvXVf2h/JAgN+fmrewtT
bpAI45HELRPDyOlb6mrbe/nkSEidD87MjyI67nNiiJDvNEKIaqFkKDtmMVi6AaBGQjCRD5+YvGlf
FckuK8xqmgdaE21qqoFKEb4JR1+hin6gPv6ADgw26GGiZ5KPdhPw4kTAv5v+3Qf5pELIiKVKdZIN
2lXHVT7W8U7179d276q3Iunv6rpBUJab5EXAXQYHiYMesnNX6z1hJCoe1qWrqzJNWBBz4TDOjc0l
nVFrLhQE5/1gfrBupJpTSFijKJdDBSla10QFAfkqP0b+Zch1I9+sXXxSb3KXfjFgMfbwgkL9dVzo
DwLc5zzPKPttR/Q8MqfYYLsObVdiadWMpdAUy08nc1AhJSAl4NPEKWq3EFiEomAVDe+m2GwGOYFI
2RuNSUX9H1TR0W01VscUmu4KQZDyx00E3UPburcXBC4XrloboJ2ZpCycgB4CMA1v+8HUn4yne2zK
oN9O8rNe8B67lgVy673pHCS0W1iW76zI/KT837ui8KKDuJTv2Yni3ljanIxrAtehOCvg8ZZ4dWSA
YfGSPw9jfLGlVLo2R5ZtC07EiBzlqlJftwIA+gPEHuCvWNlAhAefuBpjZtTsdq1GJ2usRER5F84g
bI1aqNxK9GUPlHhd3SiHAuBUxu5jns++CcLGI1kVhXgSPASjKwCcLxS2KwlgtMh+kW7lRz84Plka
8CNBz+YgU+ce3AoXjkB93OUSwdRzsu/ltEzG6iCUzrYh5NDeR/uC+FrPLFymUvxfs95kUgObJNfS
cz9wXDLvY+Oq3wR797WtUd6/wgRUydcJPEhCWWw+NWjFyqO9EYdniJ4PjC0YYe1R8IVAa/9QLYJx
BXkt3avLt4mpMln8aShL+dXElzbWxDFSz7NuJ0/kryX9FccZuYWl5daMeAFSSgm1AXPj9RpjN5no
tPOeMSNjTTKaNtw2FUrlNeCDJFIBE1coccDNdnXVO8HoXwjZ5fV44f0UQLVtHAxKcEYEYOcYg5gs
G6SNBFNWgtV0jqTIWwjKsClDSt178bpk0Ht3r4ksUVDt/fcbTscUnmxR24ma5SURmoiu8nE3KTgw
AYjIHR1PYUwgxn8hnn5OaIxl5cZxhGgM3yNvUqR9dUiXvh77dPAUmjSDJ/btgTjA2sm2aX2hdDNp
SAuALu9lTKQ28GPNCk+i6BBrzfQ2zQhF320UWD5ZlLm2JFwnh9+9rTK7NPFkVoKLFGZERKrlbOBI
l6CsM7evxUvlgV+j5HrsHMcvRFHE7r0rTvXAkc4r9fm973FA0q2FjYYdAwmB+VqDtAwKHj86Ptr6
0C3dGopox8xTQjZg8TDaj1rguLLDmOUEOpj7QS22Q0+Md1clt3UCufRydIbKPmSK1wmV4FoSZ89f
86Y8tXaxORAVlxEvtuqca4XpACejS3i4Xkhc5thVCArTzUc8/dIWUh4E4r+6YZPn3uOtyb54sNA5
TRAH2Kf1ap6JUFIvsWo0Ku3ZOMLib1yxSVog7XRpMYv1Ecb5myw48u5hjpsUO9FT0F+LAp9asDqA
gswHOP9CxD3oBa2/cV1JVCDJDTCx+vpA7P9Rs//AUmfg2IwTA73o79c9WPvsoIsBPZblz4jGlcGn
liLLoWZgTVdezN3qmYuyTIL175Qh1Dl5wmP21o6d6Txq+H7jd3CU61ZlL4gdfMJTqsRNFfnvFoXy
ZhSkB2ewcnVrGNdzluPKUcAlCaaod77rpGYHbRsgrGgKbSrdCNh2tAZjgGS7jXBaDbLe40Dh3sgo
MZ56nlX4D47pjnUMhNS/wa0MijP3wUan0Q4a5rlc8jITGrXrmcLLG6xMF+rm099uOvRCfHXL9IyP
fkDVrruhL+rlZWHAScPV+1hOYssMWomwMYjd74r+uCvJJX638MroU3a7robIyhShZ3iGRWYZm2by
+byNc0MQpu9HeO1nPaqMJvprHaOqR0c93xFinEcKUROGXhHZ3hSETsWhg6brjzk1j/D8msoyftHb
swgmvZ3KSMgu30xNhQM+ujJMFV6Umr94oT2+YWCHMsFnIJWIscKR+CLvnnPEA5qLNMNbLUmrqXa2
ylMEJtx4WREbzNygT8IkHiEpBvj+2CeqKstggIL/AjlqNytE7eA6phEPIslFHXd5A0yaor+9fggU
0iwMLgmuUY5q+PcfrLfSr4Em+ihZHPtj6FVmTARwCFw8JFl92v5ZFn+dHthdi8ChZAkGJNp0V+x3
jzL+PDAguICRPjeFVZXnogyHxKVpwXKkfb64OTpc3MVhvfi3T0x1I4MHpj1tT8OuYhFFJ06fIg6l
Nj/2g5Yu6V3kLO8qcQ5yi63c9J+NSNET7GLDprK3X29c9wL/IUn6ej5IOQC+YBGeHRwepEsYYFnZ
XOsOxl+P1ZZ2nHxkHCJiAwWpFL4DVMlbLNZqN40sTU3MhoFvYhmsKTr0hp2nMzm9zK16YYLzn1XW
3fMttIdkpGoOsAotPSbiSOjIDOqduweKMDoIkGiXHJPeQ3BcT09AgcmdQ2MR65Buuc5V/m6X15ms
yur/OOaYXnE4cofTr+BQT5tDX3fJWx4bZXsWgg0PGMqERhKH5aidOrYQSEKHYza6rl+igb0ZaEdm
ZDTBveqiuuPUx4NVOqHd98KjvVWoO1XflW93l+xoVdJq3gPSmuhFScdk8p/Vivmtf/ys4l7C2Ed8
Ss6FzJ8EJ3FWjJ2gF3+OiqipA+u45v7e5kQBbll2ID6wfOCtPV37kyyx+mlfzGVPd1NS/WCL6QjW
jd1BWR+EDYpPUdnBJSv1KOvESpxJUFEae2fCUxQMP9wd02YGk5MYvstbsfevl/9tnRJ4MRt6r7Zk
a0CXfbdtUndzAh+FxVq3vR0QuZ2Nal+nb8j/+Yhni15z42FhGuSwyI5wRFARRzQhOlycRYYq5jeo
JccjgaKqr4qvMFGG6dl8fIQ8yBI24FnoNSnW0fBCx92f18p+QuCuGIg6DeRdEMnZFtdYHO4eL1l4
RXGkGp5ZFRul3xGPJ4I7bfWKosazWA0p+IB5TRYLrzH2lAcYq6N1KTyfX05GlUA2gY0qtLySNAPQ
xG3iyVkGY4gRwTLemrDymma/YMOrys/UnynqqTwAMnyF6GHJuCVHZoh15lZIaHCv1Bf0oo5F3iJZ
R6Zw8+DVrv+Uve+btuoV/L/Lz2CgUZ2NaIoVxMKLkgeHywMxQBdAogVtdHWyfU+g6Ah+VBfX3kam
gwYawT+Qvb0SZdRxvI76nNvuKGRvkSfa8GvcRpSMthQYJnsix9ATggQUL8XbahV5QPJtPtJx/Pnr
ZS1Qz6ceZmCunQrafIhbi/N0uqiFQTrxuE8oS1SlL9ZJVQhChuzkQS73vVocLk0sRZM5qhQG7RjH
JIpUCg6HkJyqXo88kV6QF6+jrEwkSfigkVVjcPTxZmkp6ZQxltaxZOAbNJOtDlQIffGkPg7UFBOm
ZA7x4e9oLciZEI/7jazl7jtishJL0syjX4Er2tOAOPA0xsKViJWiPYxN3/+4mSGZ0mjyrjqIMlUp
cvbYXJZw+4O8SErQIMgV3IVDLEmyLqt6GCP/48WmRdW3Ye4vX+wwLuigUdPkYM41NAxOoZ4u+Hom
eG7TEOnzJdNyd0np6/ol2ZhNSiSkr4FVnbzvvBoJwZeA4iPNj8MU7Xk5lxVnxk377qo08PJRrkaM
a8y4UbjYR2fhvIL37nwJ4H25g2KAWl3RgToJcn6w/3uLnWeSpiJ7nL7asSKALhysRDe3y9DOGOOT
5xWcoiwSap2rh5TGE1sxNXZsaplW0TN/NViZjIwhtjqHWMLWpSwW6FuJ3BaUjPePoelsAkX5BXkb
XJRQNCKSfDGMYsU5kzCCD/fdZXmt0jSnTWzI+H9htEFIhekKeYM6JkNIt5EZRDVRE3ou6zRRZMHJ
YqQ0G5/sXoytsl7rQ5MTjv9Lpc8n9M0Z0s41Zv/Do0PbVp0GUyQNGr5N7RQhFq1WeH+7k/7ZT4yg
3xiSI77bmNezuYV9PXqpwjaSoHbN304SRi844/6m1NGcwaMowLApaOaKQJ1grKGx+TavyW6qMZMq
gu1D7YJ8gf59e51tLyqonsMBYNLqcw9ifHhtiUb95KyaWNqe+AkWGGa6/0QsYBow6fmt8UmCm519
gmP6j8+DHNWzSmkOAQuuIG8tinqXVwhCmc8FG7w53deHRg4lO5jljYkMc8j21KbJT/rH+v4u58IP
ieQPdBzCIPkifHLIRa6U+1iEa0bvjM0iJ4welvZ4m3MyfZ4y6N7R8wQllRmV8tNKTB9lEXxGBEjN
O/MDa+L640FP/9j45fJfDrx++Xl4kD1A1aJUdaHyrAsWjvELjzMpLwAu5IX03Dqu0JcENLiD9Kg2
AXEyZgOL8oy24oF+Uda53MC5xcDzSL5ELo9Cq8snOy4Y6scR1nMB1nnTqM+ZsDNdC1gfVVDnPqsu
tFpoz21v3F8f9G7TjMXnMDevJOZFdWrPUuxlZgIXlfmyXI32oDeCaqU0Hr0rqjT3GRMpniU8fgKh
NEcm2DKPEKw135QG0jOzwzDKMEllRO4VKIRmG+OcEyznbjp0saFvMRd5246HDh3yqkcBL+7kT4Jl
s+i0IhBxs3KhoL9Lw8Y2XaCFotYpven007MP05P0DCvwoulm63grF0jhBboJQOdPHeCt2HDateCb
JO7WCGJ9XeyEXOBbFMHYQmvxIqVFmE2bxyBT39RRM9rYTsVZPOvu7jCrZn7A1BMAcSGgKQclXQcL
tXTn1tyNmIvXEZXs5iIKUC/Xzj1B1hImXAECe0N/V46muOrs5sZO3glZ74HeLySY25yOwVWbHLf4
S4qMuSPtsxonV4pchE1d6Fkib++Wh2NQqRoSOjufTZzj/K0fxB5rprAGjkdZzxq4D7IL4tg4CJZN
efCDIyGpbUzPiL6aGrN2e9H3svCfKQamyGnGZlNVbUaRs/3XSvbcMGF04dUyvjfRExYGVKRNFU1m
3pvUFuW/v60LJCoF92J/JAAIIO+Qa06g6xjh0Fnj6rGUNDPpVXP15VczOksQ55/8rVBAbmcdL++7
P6O1shPNySMKHc53ldxVU6FDWgwf9RnVe6tejloWszOOC8qCzuhPriTWAEX0VYyV3sjeKHWW30uh
FEn23iaVnCGorMfEvnhT5XWVuBkFXuwzYmKt89GWkUDStlWadV/odiq/0AEW2m5tNDr662KGLl/B
DIib8A/JhhPidLhcxZ9HZYm4fDl7gvOvIhCNW3HPGfFv4rlRvjvC50FzzYhLJs9WBkVCK8I6QcHX
rx5EHZzmyizn1HR/yHxq1K2E8LlnW7iq5dxYfIViQ5sGgX6EuVzeMV+lfJeB2jGumwiKqENhrp7x
ftP7+prWkljcp7mp7Fzw1NqMBvfqSySgOlCW0OTI2Br4aUQ/W1yLGxho55kQZP93nzrb/4LZ2EUJ
VAsY8HBsNs7jbsxN8ErHa5XNzKk9BgKgZiCGAhhZycL4MvBS30Kth305OGAWvod5uetI8+oj3cTK
EJl80/BVt5CTYykHqXiEUVFYi1OeFD7TFG8AuKDvoMDnHEZ5w/D8C+V/H/OQnPHnglbE6yGp1ZLs
Gd0X5BviewC3B0OfT0esFTNcb56Q9/6qq2x6Owg53H8Nv+Yt4PwLQf+ELQjT7eGGGoOP2I4PvISh
NTMoxwLGTN50sjJwn4AlvPfMOF6CCsraT9JkyAd/nVIdB9tPF//QEC+TaXyjgUWkbxTUoKL9dEIz
vkdLE4RAnImbj0euZWiQ3aglbOH3sGM95vv50+2TJG1slDFYpYrzVsb1kY60iorwaNXf2xfHVA8I
TNMwtQGkJ/ZAQhYSwrIH3+0hekFbJuurXgFq4hMk5akWZrZvbBVttve5kTU6kugiWMrFPFS5Udbm
efjWzIqI3CkWLk925EnQ/2vXFXxGEW8OWLB/W7VDyc8bud9w2n/rhjDJTvErfQHZC/Onuy/8lCok
z0bvN7YrPt4RX9OEuA1uvTdvBAGxYes8waBo3/BfIHs73IMjDkTVa4YtYWvWZs0o2ocxp+L+dU2A
nwCsY8RjLV/LFbIOrsZ++A6RHaD7UUCTd4LbYUzimkYp7ZG8euB+xPIPBzpvXYKOA/in6swDOLRw
83vDFknyAGPTSm92Haq1i6DoW+24QQT1tMCaokYRz5IIDyCECY7cFOA0AXCjTLgnvtSLn0bF9p5U
+b1/477Pv3+PU88kt0XQYoSmGCPBbiShFMFHtn7SFWe4PqKkCUlRWYomMDcN0p7a2Aaz//MHzxoQ
w7Uaw+/ZW5/QaGC3vkPTVlAcYtIb6DhHZ4klctgyjxpMvIzZfycO7YXkbZw3JoLB3mtaq9IpD7+P
G8k3mVbPWYumFTRau17YrR7/XrvIfiXvJP40vJaqZdFznkp5RpDCiKX9cdrcDBU/yTTh6CR3oOLZ
asXU3ohxw02k8pbd3gHX8GTZhgkVIfZVDEHGbTKWsafvmxXO0GfX+wPzMZiUw8zzbsxmvUGsewEO
dWH9LPsuUs+gvSscNHgGRk+SWFTTj3+GIVd/Uasbw6cMAnmk2ElaxSpniNXmIvYk5U1pF9H1xWh1
ksnodeDNnWeJs4Lakb8weXefRVB56/XBOWEOCWN7l/LkwVubxeuAyrd0kPRPg8NsHc1enBClSL8k
lyNPu4RYRymfCFtpDKecRdRlFsyqAIcWMokpV7AuDoj96E/oqTQVE+tV4CIvWUpV/H8hMgKOnObu
VJHJaDfr0dl6ksS7wZIjsc2BHW94lGtJXPjEDMGOY6bEVTeiTN6CLbOVw5w4sYrhtdM7LYXdf5R7
LN6T6pgZsG1BcHkL8kT0TK4v1SrTNtWuZSUIiVJBFWfl+Jobbgtz6W17HXv+ONPgiTIy9gKMmDOb
ItTCuCfvfPkYrg1U4ZIneFL1dmShim+NgLwcPle885ES8ZdOTiISLM4d6U38oCohO1bdQAuCYZeo
kEs0cDZSOPCdI0to4SJARPipx9MJHQUiYvlLRM/vtmRD8BFR7DMCr43qmPMAo/d8FTBac7r8Za2c
u8/gaNJPlSxQn2IDaLox0HPNqG9iNVg1+nLYzUtjkJlu6wgyr7F/8vj3OTthuhi0JFXSlFS5HB0C
S3GFmyxATsxc+Y5LmO9Oa5lG1SZVHbLC7hDLpcMGOUan1D9GJFUSvyhAhamsW3q8MC41q4acupYf
buIATPuke5QcfXhOsKIoIHripf+0bMNUJr9kCc65nS7qMD4a3aq9I5pkEt0sn+MzmfyPp+med75a
wuLVeuE1AZEgfaezvg19gNpa+u/cuTzYgi6yCpCI9oEuLrS5wtb0xVLsaDGHqsvrcmPP6FdajPFi
95Qcn8s32soTh3i3UEX77gcTog8/oLF6m6yX/yWTF4WxtwnFIMHtUIngNT4B4mGVj5DZDWV0Qi+L
2lQbH22Xst05YsNmqWdQnQ3oHhG7y6Uqgzj5DY51vaVNLj7fDM0AWYnLQgy0RO8tL/xx9pmqikKA
eXvAje/JdhRB8rhQF3Ev0XWQT88BwPq734SDN66gC9qMGJ3DpdHkJ9d+GI5DekeUKGGCSBh2ST/K
kPtvAUi8r45aFMGYTq08o4+TfApdbLZx6TKaqXHK3oYF8yuwlg218zLdPjbaAT8t7CjAAJ7iQv6f
Sqmx9UYeXu6NoRYWeXTO8RMmdkMONpnZo9e6nVnxV3DEd3xiuumnA7LEIZHUOnpLOmnYR+9Sz2AN
Mq80uzXuW53NEzpYBgGh/5Srhyp6XGJyAkluY+36Y/P9m2Eyh0iA9lllTkBs35ImzTCFAJ3HSBft
bpjbE+X8UXwNdatyS05FEeZw2HsqJ9JQ4Oq7WPBDg6SwD+kiGvWiIk53TYCm9QtjupEK8lgfWGsi
B59SZDyKvFgq6YX3WqLgKM8GkQUI0e3Yyj+WZ1tO5gqY7alJz7zmep3uXhr11vHI9ZfKppP6ukSN
BPWzNYIrDvbpfmBcxVsiy7emmSs+3g2kpOEmGlMlhGZ7L4BhD0RZOhADLND3asu7nbKYdbVswrak
FiPPHlohzjdybyMx9/KmibkpqSSY/q7SVQr8kQMRAItTd0A9amNcc3er7FfPW+jxRX0RtOYZKOct
y1Kc+g6wZFP93JFbaqB+vu7AbzF+49ludLCoT6R/buAJLiT5isXWxeAJs/3xt7UcH7OiI9sp8WwW
7Y6+7oKA1DBTPeC92LTOIwZp0hdxL8Em7fVXOz26ksc8WK/BUklOFJmE/UpZqnADygEz7IGEGU83
PIUeT9XPoqDc6PxFmwYQPdUmiK+12HZ+PzXkXYzQjgoHUtMeB8ohGZ16GjLditGZs6Cy6pIyg7yL
1jCkyE3HiS3e6uiVw4SoLzq3ErRzFWSYlJijeaDhMRwbJ4Pln/xEt8EpB5VFYWTo176ioPQI8lHf
o472k7PHMxmseA36jf7LmLYFMxF2ff9X4ftu4idvQQdndnuj14JH5EDja+CfdQ69rrmxRNXh6Nyd
z7NovH0pvC8u3rJ4qmJud1fj2gwHA2aqVvAG3hAioxWuuVVFurjAobt9jV3/y9dY+ZTQKTUhd3DW
OeA9jWBMoxeiRtJ6kTbw+FlxjBwTE4YpUYFv6OEr92NavN0X4wEdSmUolD3NJxRxkhyMrPFFJbdF
CgxrCnYjh3d6fw1v0IXT6ghdFcGgiJVaUJddqAsEPXeAVajrLh8Y9XAK8UL8+364Mk7gLdFrPt9A
RWalXtuBTP3evo4rxvmq1XuYkeyxRXrtfYrLcWc4P7jfvEHBwuswP9aHdPiBbz/kQHAuoPNUeZ45
uW64Z0/LGXzMGq15WMm/UPVQrJIr4pghFjCJiFXAb2wyCfeXBfbk34NgbE2su44W15afNat/wUl7
QvOC1Y6qJM7TxoQJHTCVZvL8ser+74QjEYl9X27hp8wGFvX5wpmMuzJAuQoNUeo5CIIAEH+z+/VZ
KJBrrJLpC7T5lWEmW9AiQO3koBglFMzpHmkzTQDpkIg7foLnrRqViasR69kOFCsMJrFjGrRKmEMG
PDFtTeYdGqtVetdajofDmMlcYe5GNX5V4yG/xGcgRIWRJe/xs3vdmNjsmjNzaqBaKTHAEJgTnmGs
ViKTvJzvonGqsjTrvxKjGYxVbd5PTvFh3vsP1AWIErJIP3u1T1bi+OY8xublzMn1UXQG1YoytjVq
X7xsUrL80P+3R2KldPPYCM55/Ys3icWHfEENpfzKrHDsESP/C7flLsDYn8olobLuzbYfsplraeOz
A0EswoX8T+urWwCzUgR5HO6TBg9QXa/bk9xX/9SRERYlS1hRQiA+MS+kAivAbI4AufBC7H6vymRp
XCamxcEscvKM04SRGM+ltKzOkahRQemb7cJpkJNf+PUBOsNGNjS5+Fi+VdezDBCG75PYqxxTv/bn
qQlUjlgQibd8LGtgFfEGEui2dzxTsEh3HA5G/ji94XOSiCDKGyKwkfIPbLqLiGlpDgqBgRf2elKg
f3AFplADw8gUhL6x7fEEA/xKjODrvfU4wGavdWgSTHP01EPt4IfbS+JT1uBTxlLc4mZrT4qsyskH
B1uRXo9TdBndG1Qxkww1AU8UIWrw15WK99dVeSc8ChmesNTr9HvmjKfgsVvoj1hMn6GRwsM32NIm
bWjapvDIZgM3YE8URqVRC7Ya1gue5qWe3eI1XMa5pRYFMT5/spOJA5ptYuoRk/N40o35KNx5dZOX
dfeEhwWRHIpYrmeUiyGwce+TmOx+l0Fv89hK+rwsQUlGLe768qdMrehuXum8qj3rcpwYyYhD+1+n
m85aNMM4wO4aKCAk6vt0FHCtIE1a9qNBooJkVxDrH34IlvvP543dm08ST9oftX676+u5lO6qRY62
ZM1g6LFh7gP9R4lclWnoSRdEkIpkWVlgMldUGQDYnsrADbqFbSktVZIWsFTNHovZ7JK2DN8QsVb7
yeQl+fcAfQoe4i3JftIXs3iqmgQkULacAlydxMbpbUGO1IiD/RxDu9IdoEErqXgc0urWcBs7kYao
7pQDQFK8vkRReSimKvONNBMXpwKqcieWkTtdY157msZTxx/YgcWa/SAACyrIHF7/IwRzSusdtmBA
M7Wuq69ayNTlwVW2NnSfJfZoJFAdSnZloUsd0CFtPPHz5JNLay2QW4CIezLXy027b838OpcxPSYy
N23vgyCHcmhusqcmo9VC3CoznnCTXhaqRZF64nr6euFg1kHFKondikAWy5o5hol61jcPittJU1Nw
fEg2ikzN6kl8B+88cuNpIcuBSsOA6BqCg5Ym1TPSs1S6lEdempjU36GnznbApqG+8n3mQfexPzvu
ZNXWPDkMylLQHJ6ZW1fabX3zpldyQYpK4O/HyZ6qtmJb6tqh/D2BMwn4L9+oPjvMKDDIYEpV1/5j
FrZrvA07l4Q4fzLag69nS67apbls1JwCdc+gHPZgvDL8S7ieyUQWVSooXddfbbOAtQKaibQqwgNe
z3fWFhKRnp2++eTxT8lyx7zyfmGrteVb0/QrHp2lmg9rQ9xISl8D4vCf+p9MpCc1iyLV4nlkDWKR
emSI6sTcukqvePbP5/UhQX/825Zuz8zcmUkhAaOWOS/HFRpBdvstAeWPYnIhk/VKrcnPSViFzrQv
ConQMVK6vDDi11ZLBUbFZCkSlWnCy/sVJmjNnvg0hLbbFjBMUEZg+5iseW4zSBOmsNTK8cUdYN1A
VtZYyVs1j61fdgtql3FyjwJQvu7a/FuWxMYQL4OxyEyZzYYsP8GZJXZYkYAyhrjDmngm5/qLHdTG
DQ61YgaDnQSxGjw1IKoZvjWSFHUrF5v6r5MwVLyOLS05zQnKA0EJbDtFhxbAfYiI3BUOdtOI7z/J
41HP0zO08xg11kMGbd/cK/kcJX4nGWn9Zyu/DvtznS/fvFeBiTMeiZ47R+6C3oevzXkTcwUBxTmF
9zwy9oVR0qV46c44eVS/QLCJz8y9hzx4rd0zfON02cdoYpd3eKehx4+SGxs+EkNP9DdOxYZ0baXt
tKOVXvUmpSda0XJIgXjjC/TAvNI3NfMzGZXkzZd6V23cvxNofGezQ5BZjgQIWHks2mIelNctjUOB
6H6JCkGo/X+lR7e56iC/capCDTZhRe/V/IDAflT26r3pot5rgH4eVy4tiQxmWXbaCbmekulk8vp1
rYh9y26YGEjp/+53cgHVJzOd4Dg42dzPodMV3ZpT+h7qNUCZfEsEpdQ30TszwXGCZBwFCXcWPdce
FyEXQNahbelVg3SKR/eRLk0J9Sje0F6fbpMB6+aS9duOvF+T4XOBvUsgnXB4dxQN0Xq9Ke+3tuza
eFYOx00JOFQANzFNDhqxx6CG4N/OlJplt0EG2KxKO5EIpAi/UYpPNrKbq3StjWZVbb9wHNCgyGVA
zxM/Rq09jujNtz0i5T3TatmCAu6D8wMH8LPQ4+Tk1+H7gYBbHae4sElvQLryZ32kwbZ3b87bcxuV
/Zb38nO3O26SOrH0+hLmIOdBT5V1qY+VfnLHA2UcUslvbU1RvXm7lqXUc8TymnhjtzGfAO3XP1kA
tHYjEe8Ak/4dSo20DYEUYMk7S7PzNHlgXGv5ln3qE+HgaOGpLNZcIVnhRKw9dlLY3u/2uaJpT35V
P8p0V1XpyFgz5F9bi6PFnOVWdcGunQgoHkcZUIiRR3a7jXzskkgcKxzLtdaZHiNXmxgTPiqpcD2B
7UC1FgvqFt5BBdvxYeSDuiymAjDP4ntIK1hORmjnT+fPNdc0m/Jr7y9wRXO8jo4pw4KyAkrouLMQ
lo2CXAFiAnIymRZRpk1kCwJEQupLom0i/WMBL14uy7YtP5AFrWGJ42tjXGtiZTEl/9WSspJZeVUx
dJIa7dGNwka3Qlwiqr/nwJKwvctuImC43S3C0e2c/ZfLLUkBtO27J3TGEcH5gD29h1meop0fLojM
ae2sw8Okc1VlLHGYmcKg1AVeZ/Bh37S+i7l4z2WeDNFn9p2en7isKowByHFpHCb10WyQbBBI8jXT
KtQ1JunPp/FyoUZq/rU85SeapDMTbKcuGNRCbNfHhfEp3gyVf+TWIL8qUa/oXHivaaulJR8LPEW/
aMpdXRH0rnM2TrIzVeJSCRAfp+/yt44wEdqv9Tiz/u5kth0j8mSERxRp8amqqoo8zIVUq8Ldaiw8
iG332ApjreIJ16u71JyoS/82ijTrfv6BQKKF2mtp/M3e2OcsGiX9U4+390g9KcVijpOSMf3BVn5u
OME5oNghwZqMx+55CY2zYsZk7kF+loqkvPT2PzDl5YVFhra9mj4rrn3z946lCose2Rmr5z0kHMEH
gDwkwiL9B3G16vE4LhLXpxvkhE5FWsUCiQuGDQeKY2Km3HCoM1y+DluPPf4lDCWvisoUdx5HgWWc
Z9vGzQ9hst9LrdXR/YRSKm6hcOIrihnFs0O1iU65VTondr34UOsVQKdCcIaPg2iFQvD5vV6wvMyO
iZ16iKJRJixv02I73Lx6T9/1MFpmhBikTKVxlRWxbb+8Wrh/fmDEGu6KeRVyUh7h9f34RWDAJLCR
CA83YY6hLh2blVDVtcrpYBl8YfHhGQXp4xYrbe6iAYubCZUJeKCS8wsHEpheaNdY5xE8G2jG4KcU
iOdceT7QDkEikoEKX+BsYG71CGgc8bRqTiE9573K7DIuccjVBDPEsOXlYJvL5B8uHzBofd+BYPS2
5ejtuPmbC03OWaCHUBLqi7td7YrNd0LgT8qF2kfvR+2V4vnRjzLfvnBTs/6pwSi81MaKp/lHjj/D
bnzGjmdAhAusV7UC1PvWaBorBZB050ViVcnY6v4/2kjXZZzfZarUUqF3W1De+NnIIuzbuvpBRMLL
nJJOtrB6mkPI/Bx/qSUMrCb8c/05QxXvWek4XkWzFz1nN19DM4+tcYnx8dVhNrJYqQvFoShMIY4s
gs8KYW5hRTNYi/1b64lbzAD6+EessgSGZCRQR7cmblFO50EcDU4su73kF+KIeFtx6jStOx7fP1ak
lHYF6T0sIvxZdX0JzqHhuBHWOIq4qnomSxuueTwSOE8U5taIdJrPfI5ocL30b9GFzK+wUh3GhDYl
edtes4R3awRVuIpyXriqofmBiYs07TmadsZ8+bpWdx6N2K8AQzHVlHq2qv9nQ1qfMR2Gh72e4MkN
SsxVQm6TBm55WDnxquAVO6rFfDplDNixTfwR3aG1Puo4FgKI0P/SuGnnL0mpoNOQnbgfuSnv1sAg
JGZlggXVUojPxs9/jvbi9jst7S/k4G2Ne73muuZp0lgZgsDNEN3ojyECZavfb5jwxztF1P1RF4Nx
NodzjQQJ6p69ZFw20A9SkQc02RU1yKyl6NODvTL3H33bbnDMNzudPN7AT/JZcFJ0RyZDBd6cDksi
sER0yAeUP2tBs9hsRZEWRQGC77+6r2aFdTf5AHc9DOOHLNxxo6nk5lETaNEcjfvtTVU0OXQ2R87f
QfLfUFKLC57hnIw/1QfBD0xNrirplPgexGfZiAVVUl+HtqCDYb0q1gtVHDdZZllVqUqbJPI9S3Mv
ITD/9009r8ppeKaAxKRAfGRhd9NurxzqnmMvNZjF5UkI8MSoeczylX5ItDHKwSrdDdKYePL05B6O
817OsmztF5H2GGv/TROoGhf++S4q8EdhvqQEPMRLnbB63thVTXKlSDu4UgcTavCkmBqqR9uZt8Aw
08j5k/ae7Xf1jJEStm0qju1OOkZ/GD0cbaG6pS1eLsjkxyj+XGQN0qFQMEQcr5DPWQzURbOi2UOQ
pSkMz2FhXjs96cjgzIQnwp7YdGAdrpn4F8dDFz4CMZWiF8PXffb0p+ibwyQT7+8RDk9C/W16l/QN
wMJya6IZUZd7hY2ytaqW8MI20LU3tsOgfwkPhZGSz3+6NvLQBfuTMyAPxf2a6FydgNsNTcE8XeSR
FYxZRLbYWrt188XkMM/mczhMkZ9zlbLcKc0i13g2i14JRsy9E+trahhvWIWhdoY/Wa/BoPL62stR
+m+IQ3iiCjr483LXst493TZhYFp8vFf2vkmWqteUUSjUuT+4HFslmVCoESajdI8nKHdr/p+HcVcD
zOD1i6YeS5JcTsg9Bp7ARHEyYYsb6Q2WtODaTYw9dIdmBa8u8pbrGRC+M8496Hn2BQ8kMJoB/Wrk
kUe6tyrkHrFPzzkLjKJBVfnKvWl27W1EEV1fRJ88BlUCByd3Kyqr773Whdm1hYZjNCUYvfwzc/LP
Wv8Hg52b7+baC8KdFK1dPC5iebs05REOY7xWkntyNHEhBsDI1WpXo24PjxqJCuAM2iDWCg7BWCKg
A7IjQIEAjs3CTBI+fLUH0NZCM+x+YOGtBlth2FMK10Hb3JZ0fSatNn7WE2NVKEe03x5Xz3Zu50Xh
9MFT5YtYgLMScHrUBVSrdN+TnYMn99WpCYX9heQJrg4nm++5ddXT13TgZ06l9SY4Y+x1DpDv2lay
qciSKZ5kejzr7OSgbPniiaKXjGPqaIb0U8fK6+ySzdIJ058PNfOOH4vOxqUn/7TbeXQFU5zYCRFT
LEuxoJqJJ5TlGeO6aUJabN119s3Y0hGqpY114Gpkm6sDQHZgchy8YrpapKXvrO6cirJXI+d8mkyI
C94oCbruDmNEncOZo4XpyyGADOOAUoXXWhAzF9TaVEch8dgF2U3MK5lSs+XM2DdnDZVN9GGWIKTA
tFpuUQki6nFHRYUdYqvsL+lIgc6kbpGL7pvyA6ZZwRXIBNZvQSHliIROvZwHWUzF3GmLFBqQSz3s
ibC+JTxG47WDCQ7Bxq8mbWEHfIfJBqxANuvLhYPjQkosWQKucbJqgvRTalOJqbm0Mq2RoPF7uuSY
Xzq/2f6af9uFy72S6t8tc2e6WVo7meD2MBQDzpdmRdyZjSej045PxSuR102k8RTHpfOeKz11yylF
Q3QmSY2n7Bqq/J8txyqVYw0PuontpmOEbMyABYSNOfBxW1tknNZwLYKDKAFWkcTASxtzegScmWE/
ERa72wVNrOVdzF+Ces6AbOyPhuy+tyOGCS59PPTf6iRbBMDce1pKSVhf05Z+1Wao9Z128p1FnBRz
bGSOzBfDQJN7Q8dVkSIhJ3HRzpw6kgUTpH3kD6w9vJnM71xAYhwPg5dGhQC/UHMMXXBA64mJmBdI
CLwRHkVWtsxP5D+ZQP/5GJuiNgGsKZwtJ8B3VcYsz+TI5iER9UPjZGF75kWPtFK5EIi3JBR2Tpae
d3B9bJKAVLt0pigZzJ4LekJ2duaiH2KZXyXhHHWDYGP1qcFgcgH8e3PfeT34T7N/Z4V9fXBB4weF
4darAhfza978uE5KULQHsyn3Nq/76MvXQzt9v/EJoI87SZnViFNltPJTJcUcQEJSQAVarKR/kk7o
behxUOj5FyKN+bycS75YMk8pqi2B3CuEliZHi3P99iWMELwLBqwZxevp3YYm/MC91fDzhlJF1y93
CrFjCcYLGOPyyTxn+8LHwBTsWMbxNm7yYLrBF6N+zwl+9JTI5wfuicsTcQP3ZMIIKnLaCacrICYM
dHFU4x0p2MoZfSbkNYzb3eI1rhbifGYNzkih6iCvQ+NMyyEMYxUUrIsRlo57fyW3xad8EDz1C8S/
oqe+9rgnKgwO6mgc+kJzcAH57PcQgzsKxkrD6Euh4cC/vflOqGvWqz5o0oTdw40tKDje5mQa9SEg
x6j3KkgVQQ3YQdriL9Yf8Qywj66yRzJ6popuRFUTYZgNU85Z7VlAGqxcNHvaNCyIqPD4E9J/YiBj
gk+JEzwSqmOeZBmVeugAQ2WOh3wVULAXNIzAI/fwOBIvhT9hQs7Gspy+gtEzabobyFg1/768Hv2H
+HyZKjdAM1G4C4F1j9wP9tI+VbspnURDqZk5y0SVjx35BehcFBr2rvsNjf9RvdNyW/osclUscH4b
4QK/wZotuY5ky0bunQ5yv9kgO/5QTclZhVDsOnPI9hdLDzAwTojnOnGLICl3P8jw+0PC9tjc698d
ozf8idv3msa2nfppINHyPNYA2W0HW7Q77Co4PDBDJVaB3Ku60hErM0/1hK3Qjv1bZKZ5Qyk8jOB6
FpVSZF++xyskHGvgWmI1DNYEeQu+IlYR7dU6mF+58r2+eRz5j2d1mh5OErkbd/rinGxxxfrEs8Gs
QZFSM+7IhLg1ZihSy8buz8EYqi4DA+nq1REXfRkR4jpWZvbZdIUnlhLtXfYO1CyqPn8Sk1ILSlMp
RJFviJfreA8giQQTYZib+Ovd0CZHHGxMEKTT5zJyPVgzmLfhgBk9RVNvJnKq//Ddtti43gXaIliC
YC55VvWDXMD3J4lSu7rD68gjmZYHoUVsw+17MLYpYk+OXq6WMUDIaIdZFukicSzCmS70PFnQMVyi
ykFbx4JB7tyb5s8N2zy25FZpSTBJUS1yzXzo7+0wOvcdHtUBgujWpAtkyBBdustDixGNY6PWPLYA
VmR+c9jYgwCaNyneK+MUOUUlHIWf8zY9TXcgCirGz/yKPocnl9wYa9fJeGitMGm4hOyvVMwfNfda
LXdtoAacBg19ur55G5OYdhwwZk+4+Y3zPQ4g2L6ZPaDVKWhKprrYVzYkPUXL6IoW1J97jkCsS7nF
8vCaYJ4+2ON5SQHI1qGu8F2LRHZtFFwIj6oFIYKyVzgvn5FMppYHRx/sk+hJrDQtAfBA97gLPVTZ
bBSZrGoEKjiZuAJq+6+84MKVZgNucV0MbgbdOQ2eLN4nDmyj4zH+na/NGeFaWmGM4lhRixK6rWXo
jDklZ4V0J1PeTKq878RUF6qitL4jRmtMxYF95VCcMDiLHeZZTFhYX2zw7ien5JMoEiaYZPugRgzq
n2sARtg8EsauBnoQnPrK7MINHuskpSBjHw0mZxwUROdNdCmJ+532FEBceuiDjJ3Ohu/wl0t1CxHv
N9F0JPO4WI7gBuUNUyiu2hSjaVUaiiFZfE+v7atTSL+cFfYg0slJaTkNL+R9LS5Tjs5kHcMUFKkB
QniU4i6/t29o77xQY1l/Jom4mnHxGneAdA65iv7TG20TdgzbbAnm1Uh38ZhhWbDslLiB11gRI4qQ
1kQqiM21Pu4+LI3RXR8LEgVHmMNk+dK2OYN0mXFsQ4VYV5cUy/qVcLGf5ZytjKz7rxLatlEbOrTG
lyDP9j4BdR8Qp6sbCf3PklTqz3l/98pUmuA42w4BTaGpgJt2l0VIPVKnaI3J/ZnWCWsEog9IwXM7
SUDbo+U8a4dGsIwyPPu6xE38NyMBZezXD2StqQuC8IFnOA7f5+FvNGHYjgVp9mB8sKPVjgpMTz9o
uBdB4fGoAHxj6/e52oS2cELj38OJVgtuvyfLP7Az1Kg9bGzeYu7kbLa6POAf178pWIC4+ahrBfYv
iDulEP0iBMXCwxbG5PX4k22RTSEhWMPiwU9dGbh2ie/XFde0BuG6sz+rq3eA69Ek83xRhK+xE/F2
jkvuKYf6Bqg7DIovNQoTHRVCWWs3gs2fesOxsWM/YlVI6n2AjzOx3A2XE27dLN9Ncbo/8MaME/uJ
9b96maHehTtdTu3a+7mtbVl5FJRsklH9j65KUN6pfFqxI+J8vcEnt96rupPJvBW8NT8hbpWhLWsR
N7lywlqZxRIHOZiOwaW1A78HMsYZwJDdHxkHxPlFCcuaYUpdPkVH/qIEjZoLGqQkaFypHOuGNhFB
vFBlFlC6O4u+gq7q+RIRU9jZ0tKYifVCtEpvb58g3wzzZpFlte65SmoLUh6YY+hEoTSyJkl8wV/8
DUoeJyZdCC4yzf6SHJu3uXjxccjE0js4s95+7VEt+cKcL3/KGAZAL2EtGfZcqkUujYIef3SX0YPX
RVWrCXnHMvoLaLKOOEOH0yjIoiqiKsOXw92L6ak0oCWk4+VphgTuoYDyuhcgJObi4fQM1FSDr6XM
8tsvROQhaJ+lLZgwFOK8N+EKxuzHYw5LW+kjCRtMRtrp+5sDNnT8aslKr1NP3Lqn8qgm+6A3ZyMh
P8BkBs0XNdR1U+SGA2EZYoqBFL9oivVlqqY0ogVgENJvy91qSCFM7zUzIsEG/kL3o4XF+XibfbIF
IICIsAzN92Djw2nTKSrM7y26VCYuy9FuZmH55p8tq0Q5os2RvLMxayJLB2uCRlrzU88jJJNCuxwt
0c80Mh/q4p2+uY0ZsmAStdNtEC+hDgkwzSijj/u5gIb7RTr1JTgvODMaQJ66S62aS/ffG8sEHLOL
l3xfw/MosMLLSFDayZQgsFRXsivAKUG5QlMwXUFKzJC7qlPb9vCWbSrlIQ89JYVGBLg1nFG8GUsn
EkHpeQWcA5VJbMDI9gfa1I3w2pMMfo9QcmWqSKizwbtsXL/WYRONjD0vInn7UONONsq6DucQFBWM
8wVknluqzmtHOE8scNQacsb0XUjNRM8iOaA7ZRshgFAjfZCDncujLzzCi2ncBTonAFlMdwwtPOZP
1r1x0/YBTNoNGVbifjfj077QOFxmMzLLf+Y+De3wZ1IAb/JqjEAjHE1GQ73j6wiln34Ft+prLR1r
mdvopmIx9W9pLiKCX4FRBb92krpvJ6jfdndkuQx0DHNkHX+NFltviHTBVdYFYw8u4FRbGZTTgQ3O
BLv8CdgtKTqg7grXimUdBrZa5NI4vo56RKCSwB7IXRJNi+fm3h91cDfjqYoVaGq2XKHpH5LfWZZY
kopTAWMZT9YPzHaaDSWUncL6crFuileyZATSE64tPRWdd1yJcrXFeYKJzbMmo7bcYBYfW4GH6d/l
+FtfjUXW+OZ7r5awEee3YIjR6CtsL6UrXCDg5lX91ZQSIhzFclt8oRFHdlfJPcr0roqgPP0jAffe
8rqXpry98ZQHF1z2tMwXQYIYZNi5yP7iDgI+DVpy1QrJzDdDxRotcqlAxesZdnkyPHQNtF39FHD1
xzb+hwoQXsaK4QzE6u4sICu+I7zXXrJpcc9rrfmqiow4HhqQYqXw7/tRUlIgeUisWYbPGT1iKkO9
WqmBsaB3g1yGhm3biRLcyfyN57qE8DQjSiCfWZY41JD5mhbW8YwwGsh0Y5tde3ACsXyD6Z4ZxobY
k6UM4stZBbRdCfwCdWsoacGYsJgKqnWCfNR1T/5uyrBrFonUmXUwU9mLfOi9QeXqVouR9kKsoQp7
2RkX/HUGpEh8188MOHYuOgJonC7BgyLDWR6l4rpyH3vaIMYmerV1ztyDw7aliqUDpVKo+WobsOzO
UxyxNuc9Aj1Ow4hyhK4sTTaUyQLjRArOHmlhPNT2cPXNp4WkSzQVTDAj9CLV7jqnIqJlscsLyN+W
PcGX5s1y08afAJrKCzVKXq04Mp6Wfl5gvDxAMjRsyK70Rblryk3hAj8Lh87zUnSbwyx8WsuM6Uhn
x2Fh3kqsRtj1K2VoN59WZn9CrJowMvdFrZn1ijUZ+x9cNUCYLQ11g1q8A3oB5GFqC3yIM8c6qU5j
gAXjqfQw9h3rjOQduLzt3g78VZ/pd4WW0LYUWQg9yGXtTdlO4JyY4eK9dzCpOJy/9D5JaU5h2hyM
S4r0GfwqeL/bnJT5CjmDjXtaKHy5LoROPYo999HrrMQy7W0zwuGYBZdpEUAfUHZ21MnmXGWXOEWI
TpZVTom+igsi2DarAmvRgr1g/qb6hkRr7iiUM0nYqTaOCxpJfx9WOAgEq+ciK7IQNgZIagex4aQg
s245awLsarH1ELDRa73zG6hk4iA4OL/Z9s5uho55eB/A6su69mUJm0bol86h/H8GCfNppxaUkshM
76nB94uCAUgNnmzZn5OOe1Ls0Sn1vwlo4eUUCcN1uqPl6/5wo2fqFD1kSNw088WbwxtHa3oLUp1l
Xv6u79joOyzFWbBwl2i+/Xwfey6dT/Pvf8nFx112IAo6JG/IqkxRe/b1DsuF9cSSbTFU/IUfmG/Z
fptD5h57oqr10rrmnOtOTvn/UKuTBvK43A4/yyJxzEWO9FgnRrztNTSmY5ppoQu0WO2+B4U08WWS
McUQ+8ivdnjAzvn/TDdsjf+Fr+G513fO+fq48VoJV1cXYrjyeCjoD/pcAAczjh/91RDIYrcE8fSu
5pxr8frQCIttlmfOU4vXKIV2Fr8R1cmWZjny6AMmdY0Gev0cY6MSo10ldnfZG0WLbuyqdjwqtgJy
Wt2hz37FKuijxBlYcib8dphI4fqhJdVeHAB+8hR+N5yz8e7b3h59ZG1Fvw7tV4649WY5LTdKvM15
Sq9mvcyD9p7XzWIUOHpuabkMBdBUAg0gpAYNnu81Gg/7aQ46FokkM87MAXhgpqb17fg1YvjVYYRt
jROquMhOLOJTLberqapwcNKKzLXJekVBrUbFtsY3os6RAXL/mGF6hF7EGhvQHz5CEixKrrS2Ygcy
uUwlr6lESkGsQBDQW+Jk3OuQUK0JAaBfg6nnWkNPTcbSJyZC/BQpDRGXBGqrG2luCRBlD2Z4M2cW
cbjYiGNeERLiYGgzMK8A0tfJh/ouIcJp3t9s4nBRwU+sMETb9WOSpkEqYbnpmVf7zPaDpzgHZrs4
kd86e7+TdUPwkedx+//5oh/KxieFbjEI/2OvLPe1QZpl7sbPP1q4VTNaSiZlhOVKuBqqUxCJQQar
0MtRJvxRRujwhcYrjqwLjXbXqPtDCIang/ljNxfv+QNzPmbqGShZcMCS0j0CimWhW0xso5cL9Ws/
tOJJkSV3k7Ybg/8jrTqU7FfDVZh93PJZDqyHdhePCC75kOQOmGGzUMwAsqhg8/0KzHXZuCPMajyM
oPdsXt9xFJ+7cfMaTwnuHDkX7gpgvSFNY4D6yhjR8xE91QMR6LR4xeUZLoCt0z+wnBdJiuVGXyQJ
QSf7jEGiuSTZrQSBOkmuYGnEaFbYCdZzdf92OIreWzrhMFJ8pl0acgmh0rGYzD50zl8eMLMxEXuu
R/DTgEEE3pSSmVb1v9Rr9Yt/oh3Zlk4kMP4Mo1Vh+qBnb7Lku9r+jSSMS9Ei7Q68cPjAJ7wMEUr8
ZFkirbxFWxQNiX/UHfpOfcXfs/ijnI2SRBmxQICConSOXwYz1C2YUVjbg4nFQBFN45u+U89Pv+NS
rDn+BMZPoDoIdixEvy0jydvAkqsjpQzBu08+ldFrXy31UrGQnJspdsdlc+n9cs+t4nNXHaYi5iHk
ZT09H+wRV6fBKpAF7cIVZ4LMJ3dPbCyhlE0nPG9KxMPNieFuSImJqh2OID3xY3RZm+vqe/9UBlzC
tpjIYK2AdxZjEfpWeuvPxI+lJKHTLe635ksCWxnL60iWu6VIlb6KPAUWTuA/C31kPXgF+QkXIzky
L+jsRyFx6M/Kav1gPMl9QrpB4rbYWpQP/cvxfp19yfupQAHKZZ2AlWN1AIYlMEzz/TF5vr/l94mM
8ZETZVTt4+U866zxvdzy+Awos3Np4iVrD3VJgcAD5vWDnv5561S9CkuQejvOW/abyJuRRHleOcl+
cK4g+NwV2vYBZyHErC2RS0NzAk4KPovrR5dJ/SLOWq8dFAUiaIiXqCurcvqMKrsRrN7VcrsFnwuf
Qq0qcOWh5hZf9rdM3yNtniS1LeRNMcAMqx82+X26aFxvOWZJ7iARsot629XPvgmfZo8cmMWgycHa
2khwJeIISZ1pzczjIKLo6OBShGp2Vgs50D+Wk1fXVtCcPZ901LtUUKhSb+OiQZ6zIq3iTJtGHY0+
YI5mbKv7co9FPEDleH++Fxa0spaLu0BxFn2hC8I7Jkt3EteLfUhfpkDwbrfuLfJEN5EjCty+Hppg
QmGvrwRruUrasjFVuWlqMovAKsTvbzg1uN4ZScPLFsx8Nz94pyb1u2lFJB9DtbEmDrwYNBD6aQIw
3t1AsxcsHw9qk3sBIyDChJ4Po26iLkJ/OWbTy/OZPqY7arpHfQLYr9vceQ7PsOXLSG0Ql1impNee
ghlLf45mByhP2akLCLwf7icoZJ3YgqwysmD9y4rejj/6WOmk9ErQayHVVJm+anRSZHhiUOiqnmhI
iFAwrcwMiENvKQC8I1aQ1jVIm+x6tMMOVT0rKCT8LbwB6S5XMCSrTSqIP+Y4bhltQ146etx19ilJ
Wr8onNm+04PkM/ybRr2GIgz19SCLYUS5V5j82hd+FesWV9AF6bnl8dRDY32rFZAJN7cTJzxBx3n6
WzirReN2uTqEJimo19Eple1oSCJm9GgNxb0R6P2K4/ywIdLu8v3IQZ4EAb9/vTadP5bVSOSRFyMr
HuxEsjyMudlk84zXUih4Nm58QfgAYKsL/858yXOY1vjPENelVm1pEwOO/1Eo4XYG2/ZQMYqaKBbg
RD5Y4RbE8hQwUSe7VKXc0mHr0c3wLWbms+Ej/7XnFayblc4L0VXoWxMDjJsBq5lwhhp+mSy9Okqu
meb1xmac/hDA8cCCpipkre0ej2rAxzYpc3zqe3wL+AtyzP81nYZfINzeCRI4p/cIYUMuhau3/eNc
BrOFvOxZMo36lsDX/qBPLw/nmhJv9r5TsQ+iP1pj43Zr1+zGjUMUVmAU9QgXFZV0tE/OoV4RqOTN
1WFmmEGvqu1uVJPBGnix+5HL8C4+oJ2NofXVZnwl1JwgXW5Ze1APDUJgjKQlLYACKPrGiK/VOMgE
bKBd1DoOTg0dszZC7OtNxeoWcGVXOnlZJ9J1SaQrUW0v/s+mkSnmrmJ9Jn0zuJRWpib/usr43FUZ
0IvYNF9eYyGlG4jxV8uNUZIMhJT2i6F8w+O0g2rd7+jRJdRDLKLwNi/2eyXbLDF71Ts4xFSIYqH5
boNTJAKjUmnKOoWfmiCVod6dAZPTVQjx25Uht6sq1PFGGTnIJpTwQA1c5a2yExoToOhDyZTiIkWt
nc9hE0jTs0JpjOWOHBC88H2hPaBY+fmst+nlZvc1J+zM/scW2FHpOhS8CRnIzN079C7UVXVHWKYk
vPUQaYRK5cpYGN97zPW3lhLnNllyGGEedcLtw/MxM4yO4iLJGHRjhYJPpWy9sBOHnRnIkWBl7O7Y
xkkENFqpv/79OAgHW9PInCFAM99exYCo0cfU0EvKVrzJaxcVmBE6q4yxtpxFr8sSydarrCIBC7KC
H6J+LpBDmPAY8eYUlBzyuHTf9comXmHMt4hUgk1Uo+jUwv5BBKa8Us2cQZ5N7gJOc+M0iKSo8IXt
I5Nj+wXKNE9dpCz1HJwYzQG1PSssT1ta1CKiCfFEe0yIIuMz7No8r5eENjcKx6row3X+sNrWwcAk
0pyZzZ16lqgiNm34Ear3P86sOhzbR5WcYAO+Ec9NbNrX4UX+Xm2ulWprQ7zAQoZV3YmKoz2fL7Yc
pDtMATrwgA7YRWxrK4zeQuAcy2MR/x8VuaWIYsYMGXr+YNOIijiwP06OVK7e6ytJ1sjUK01f0LuI
9Ny0rij5pFiZh2+zXJVNMqyxgtBMVzvhDJQgIZV9HDu/LfjqXCKftWCLoldJKt5DHT19a/0Mg1jB
G5JPbm96bLFXI541SNOo5OlFZo+lJIeJXFMjio9ABCdzUpCFAVrBUEkWB+As19QLIA3rkODQbLcr
XtDOv4IZ94ZYFrZQFXza6u0YXceshoOgYXQ14cwcA6k5IDoT2HyRbxhZLw4LfaRxGmiOqCY/KB2Z
8kh4IvM62+8BSVSz8IaMXcE76JBzUbm3Kvgl8g1p5Q9+PKqNzgiywXrhdC7HAjtbwiVY7A/USs4U
8UFiIHmi0IHIniDpVnCIRKaXu6BzbPf/Tbktfkfe1TCBufFaX+IIH8PJ9QX3vlOHEIXu0ITg845p
0iVGUB4PmPovPq3Vif2c2jvpx8NFy4QTzX2inBTe3jIkyU2nXFTqRgeMGXdmdya33QC5xSsS4zq5
zXY12IFFRS01ueF+uNIxHmC/ibw7uF2E90FoJWhA5Ghqn6fRnTa1mVdEK+CiFtfAUa+j6B8nIq/t
9OJA00FMGiTjObxpD+jdVa3Hny0o6yG1xcWRp0f0zsdATHfg/X9WnumkV2Hfqi0UBhdGhzujmDIV
6e/uIrkdR4faBY2QvrpovUd9lg/Mt6tNoH8daEu6GSePkaSnn6qabfzhC6V3uOay7if6X+yJOIO6
HPpL0AmuVWUL8nv9Y+90okue55GvNG1rdBufuGLrOpgleZDa1cu6bjoxF1m2QQG7eGKw4ircQNVt
ZwlywI67P4zXh7Kb5qmq10vhQ5hI7mjEu3u8ioelLNK7pcG9WRE7zJcyRgzrWkH44YMc9XBt9Q5D
kJTp+qYWEVH/6iQANIHcQVX+iKp/iUVYgCajoF18uHMX4nFJ3gl7Dwj3zjVo2i1bXAyvAtQ6FsK6
vt+yVvw/TmBEHfPtZC2ktW5x2sTZER3OqPM9wf7DDn+nZRk1FsZjCSHOi+zK0xkITfvb/nPVpOw9
jWtXLUk4BJqL86LbOX4E5884JIpv8RBm8DM4gpaOGwk2wfPZM35NH7wym47NqJijl1bSz3zjBL66
3mi+VteAJ5J+E1/pDNvR++lqcjksCLmqn6J03YM0vlYFENiOZaflMVJm+6DSXW3T9oICRr0DicGg
uBWeaUK3D/4V62kdY5xrod6K4zW6Hv7DVYKqVo0B67qrISPPBFH1I4WE/eH6w7CuOCOFrf8+p16H
asJH8364b6xv4J5z+hpbMHlbWLTFfUBI9ANph9Cw8JvFKzVVGl2qoe9GNmTbMk6WUq3RBXMF5nzO
8SI6WXD0bxJS/GykRX5J7kaCCRxFwnf42LF5uwespBDRfrpch0d7CtflZ3TgglLxJBKBNQFc9lBF
w+gwLQd/ENDe4z+MAHnNn1zNGU6xDms5+D1yY2V95QxRDZTKsVcq6MaGtSlw7OV44W85M4mT1DWU
QD3j/kSTo6kF1hxbaxe+vig24YNl7i4IvEzNLgn/su0z5x3jigD8P6rBDR50XlS6o8fGQKD1X+nl
s/mwZK7rPIZLeZoWLmwhES6FnwOL/4fsT8Zv2AJYSh4EqK40DsLfMPik2lrFkEEp3M+l9/1CBlHI
tRkuTFX1HRMoSx0YuFTDc9ev5c/B5a/Nfw6AZ3nkh6J/dndgOqBXJ0OYWE6VLgDJzJ7UpdCVjgJ1
P/TzTHzDa6DDWkmF5oaHz7iLPDPm6TounAA6tataK4amgxic4qB8kBbHijedmBDcYHLUAiyIsguc
UvwDfmMt+brCpB2MH7p7ScLhYuLWKKwJyMeNcYBiWlPTO/UWl6O8Sy4cWYR8STT2Bw5r6Lb0U4yI
e6PPD8+dkxFddJ6Bev0muIz3Pp3oppsKyCLgXLusnu0VDg4jW4ic0fCOhI7FH9jkMYFyftrbf6Eh
KPyhutn15gqKuwKT0yCcULfy2+VnrrEmWJtDRhD8nAMtZKP8pfqahVUk2ffAEBkcCces6cFZA51x
5NruYeg/QH3v7vSW7yhH6pNT88IpdbQ7tK4KvQSLdR++DyMdyM/xh9miIViA2S2/DqzxSXPqbsIS
pkJt6O7r5puvd4O92iQQRRLpcnjKyRbn4JcMBvGXkvxNZcKbB5UA2arRJY1Ek6gmGPMzWuyXBROz
2PrmKl9UXjgfnYid4fQBvYYV9zC6tW8V/pV89i7zOF5urRAf033heeF4dLKHKtcHSigNITq0o4ND
dypve8Oed3s3bZa7za3ILxScw6dszExeh0kEDTX299nSH+PBCKkqeqzUcuYIhpek1q2aKOm/o95F
pVNJutywyvvfdkEefhuep6SSEytai4OaQtzTcT98P8yQW7Jt0+3IeDSc1KaysN/DSGGAeSTH1nDe
7cFFfxE51dMZ6PHlXfOX9F8VzlrNES2//ASq9ewDxTl6oYV/1jtk9WbpLvcHvnqxmcGVvZzDSMMR
cR31s4jn6lv1WaCT6daiwOTlCw/5FThk3RVjegM19dsK7lXTQ5Rz6JerAhp0b/V1CFwv/Hjp9eUS
6EiPAsduZNzHcAyfUCvmK/z84jF95kULWw+Lc9JWZ+yauSCXskga3/nzwzT4zJMrPicIRh0+x5lK
P/m73VETTMk7G3jsc8LSSforOmroD8EJ1qmhFEvvUtK/4sGeK99GiRZ3Cyo1/ljti1uMxxWbJy1Y
UW4DATdiYJd8eirZcCR8MzC39hkJ3wSTkvRS9EspALx7DcZo0rv6ZX1OzCLbZhS/zijNjnxKQinY
BD0/j+rZRX5q/SE8XSjrx6n956yWzVoFRDt3xyTeOBts0FVCO2Dj2qmyZvXZrJQB78DRZS16bVAW
ad9IbEOTsEUh8QbCFrrH97a7I+O1/hZMR0jK+nsoisryO7+w+HN5WmcJNq4fY/tQyrbPhRvRquon
DfYCL7onLP6DvlJbBjOj0UnjbbvvlNbs66C/7ya7CAZS5kwillOF/1lYn3eArR3VSkhWoAjCnGNs
48NrPYMWcP6DAs9F+yn2nyobavNybXGirESJalUEi+/iOIaA7Aj4mm32haRxvKFCZbm5xQxwaE7y
S+5ze+WLKLOdrsf5dHzHFIISZeqWUSicVMXw634D/7ORor6jw6lYYdyORQBI+ezN3gO89xfr6/n5
nRgnPkNPao+G/ozKtfWBoA/uxiWqkK/gUCyfF4Q3kDUiIleatBVnDYV0ZemhRZTn9TJPldxJvn+Q
fIzT9dRmfPcGRFXcijC358VpxTUoi3Mlo9WT/6at37jQb2pW51Dw3Y7golbcUO4mR4XKis9c00LP
xTNMfpkS7u0/ZJIE2rLjg88XoAJrrgn1mC6gnVHLDawu5IrkJzNkhT6R1EONMVq9Wsvmaz9IGdQS
JTIo5Fw79nCj/+FXr/9wJopCwRr9ihIyk1txsXeqbNvz51ENnTI9w/ZzePNfj0/Tww5EVa+SVYjO
KjIFpyhh1q5yQ/YKgha/X+FP03Mah+OwCz3zagYLoGSUl/lI8M7pCrI0rgH/rlQE2nOsH7esbBkk
KxExY9mD/cfNkNfGK6a2kE7n3jp78rdW2haTjo/TJkRHsJZ5EikPo6tIrsRucigdj7ueXy1hDpVY
+gHCFIvIgwZNrATGqV7k71VcpqmYUTqkwLGVQ039+3EJ+O2Sgv7YduImO6/W7693hHY6jcW/E4jE
8xQQNuJkmjkPTmOpHvowGsO8m6KijIHhg7K3jjhwI4QZDgqiXFYNTZ649LazfQUIB+TavXR0kIIF
Ae9tBewqClt6IwQB9jEIlhSn30SM2DE2yAgVUGKT2rXq/+Z4pGaKlM7vG/Y5FM9PFqSq7ameadzY
G/1L82D6sxLcZsVJSfOFRULTAKzBv14siTcnmOG0CQ45zjtnGuK4gjlNK9DoNYVyEaiKGDWtBetH
thuZgp5e3UKRjD27epq21pX2HDE3aAE2tDnTRfaGH/2JT0L428+fISbloCy4cnaCPqFvhIsBqHkU
h9zZuMelGq0fDJE67OGvYgqQDilz48L5KpWuW1EwZwvwZ3tJH+2PLqNiEvVjSowMxvv5uYZO7UM7
ajbZripsaABQVvXN6OuHNDkU6ojtjeahn6rDn7PDHNAWUAtMH87L/RuGu397el0of9vlAff1P1Bc
3y9D8cUgHzR66sg49y6rocCa89bqLOLEpsyRC9Gapa5V5RgEnk99Ki+8X34o69zFwyr2efMotQn9
s8LuxtFvrOhtzrBc4qZJa8zZ6ivE7fHZyAEqAWY8kSOzDswtP+0l67dU4bKd5HtAoPdoO6NiNvH1
8/4Y8eTL22wTpgk0uwOc6z2XpojxTChqS9LftrHhH7i51cDn3ZC1SYCLcYVLT62xhCrmbWk5Ouer
6kyKytavd08oRolrV+32ffGOrGM1lji/sM5IWCjGHnJpJqyECPOLLEUWxiretwfBy8O8YA6GZJMZ
asvTslgRr09xIuIwGYhy+crw9Su8KVMcbv8GusuljCC4Lo5USPardk2tYnS8lJH7qse9wuy+4Utj
PS1rEkL6pCxoSt8SXpe8zyqIUyaqsMXDtc8DeF3v600E+7zA2BDjYt3YAa2qxcAg+wS/UOvwjm1j
a44bjy3iePY4ifFz0puhk3c+ClFgF5T4kaQuW6QQfLmcBOUe0p2MvCD7QWTN8kolOo2LJuRNZgN1
bsdleH0ojkOAYAZ6Y234uwI5s5MW+Db+VrQ8WOlXfLmARb79Fqmlk76oxD+t072uYCDjpmu+nH/F
KNwYcfxNPt6zKsztB4L0G73a85cfryFuTjQY2PXxCXIs6QAi2l9GoDINfOf84A3csaHxsyRZo9h+
8FkDgD+OEUSoGjc/dpX7LdWdQtx7pCCKWBnfEgnu4M63uHjCPNPFP8k0/tt4LE2XXxN3GHbgnGht
EDeyB7JHcebqBB7cQkNy4RDg7fDLgEDE//95dV3WJ3pUGtP6stu+R7vFVscGjCQzekf/qYiFbQDv
kk/5FR6mtTCFlAwhaT+9ZGBeX0eN1khWnUtkkUFF6I16WrX10Ib4rM2RZQ103LTGgENaZQJeteru
mPqtvgrhIYYlph895buda343SxeVrDDiLNOSAR/BlP9RvC+HGLsP2jPWzql+2sKQSlDpp9yT0CQB
m94z3qty4Atp4kaFKItrsabghLs7sJpkGqnwB0h0IPhDEbEyXstHpKTe5ge/7jYFOnWGn/cKvVkd
bMbCUtGK75R627iQEHWqUamgMsOC18MCl5eKS7fvj7W7IvMg9ZYjC2QofyFNTni4LSWwK0gCy1Bl
OgaoxszZXsMpym5Ig4BciiPNNsscHZUqy2VymyFJS3NpGZUtlYW+qEXBrmFD/kbBybPpZhBBTeDI
rOzh5c0xED7kdLKQjvJXxw3wPnEsOF/FCaFn+Ur0OgIXRgBcLftKD8UzGtd6XB97o0n4CeHZ/FTP
TSFMOW6CK/N6J7tgmFc6zot9urk3C5g9JxbRofGVhND/vAqTNYTcUfP3bdr9O49mpCzIIN/ao+kx
fHxY7GWM5mQPihbG7k/+2W5/dZkgJ3tgq3aX4eDlR+1KDkOb3MaOlMb2BOnCU1KnFLXG/igEUBax
cJ5wM5Fx/R6DrrRo1dJqLWlYtKYS7KVIWAp1EbQvvPtTMzlZ/4jSs6KfOJNzrcm0NjCWf+a2/1y3
ahuzUr8txI/7YRYlY97/VtoxzhA/6EZjjMf62q5WB9EavFX1OGnd9lrxZcrcjPI9y34k1Q68vUPj
5SOY4ws33K11ra5OwnyAA4zQq7qOA8ovalRN293Fh+GBu3otdUDu1JtUQ5H/oJeeOh9bJZjA/bqu
2kzH4EJt4kV/M0Sx2D/h8sAgjaMxjmxzkc1cePiZhMFzchAzPVWDvCW7gx2ccr8FyCw+HlD5uhS+
VugEU5CFdgkPleu1RlsRtC9KHVay5Ve3MG5byq+K1c+CX6rvfqfkMeNi0CNeKoOzXq9dBJCWBTYd
ARNSJ/cfmnbFsLTFh0oeSR/DEc9j1t2k+GSR/UFSTZ8RmI7JbHVspfjj6EZ6YqpH5b7Vm8ZpvDfs
AEIQotMnipxwU1X1/MbxcQbb1klbaD2t0VUxSMdKKeobKum6ylHmsfTiqw4QU+MFtvr+V4DaGBFv
wMCPgAyOuH17BpOgMt5hFtNid3o0kPm5Qrm5TI6hChXE+tvqZYwmxO/ssBpun5KWB8DXd0KAjoU9
MZ2Kq03ouHkpbVImcPewgXvej+oKSMW6GHG3rpSvdsK+PKL+ZHfFpUJdQNosvdLjbMhFLUMjRlnS
fcAydSf+7FsXl1vhsERGK0d0aOpkRylO3VBiXIDGq1FVdcjpAnIlIsQVk6k+1irgNxBQ9Z0/Uo8w
WCUN+sUoqU50RvYaidkUpJ3NN7vf3BoAbUl+mTIMfnMp/j9E7WCuVIYYaoRtuelk2ktEsE0aZ7ri
ENiDa+2KSeNPomUsmk/7es8jBlfK4Law+4xMRMCLxb/lirIEqxDKT1C2z0ByuLpMO+nQ6bGA0NWa
YKwO33pnU8dwcvjnsgTjnXRNEyl06q1DlOPVWxd62ysxzQisSQcnND8lx01kxQqveBRIiS44OBpd
S326a0qIuHu3Z1Vqx0ITGO0NK58DAiJinkzTtCkyv8WrD6YpRJskApl58eT1SwOo3U+lF296BLf7
gB7+f9FJfKSSgvod2I+4+y1qiUgC7hHwhpq+gkYW4rDpI0QphWPPPE+FyTc6q2y/hkyfpqRi/y/U
zYHkKcG47yQqn1eTVHVIAw5rLQODK8D0ZH4T1plkkemc1momeZrFGj86ENV8DbUKRcLA0mb2sW9p
MmxapHPLUc22PdVDzHG3rYfkQ4HB0TGEZf0tADErIiVhITSK2I2XbzA5iblLXgGylYGy7w3Vr4i+
CNvm5lDkeHB6R3oXlNEYD2y6uxozC3cmu3zVSAP1xBbAxyIlHC+eEuTDTKicbNCXm7K199xxDS2Y
lB/L8+sw3pTXdmN7qViYZA15drRrEsdgWTvYG9hz0xHziQmbdl2fv2ogO3I7sPhcmmIVD224Ph+4
CoNwwoTeS78RG1DT8k6M7lj+DQH0hA1nYCSaHVBPTYeHhR+B4Yn5GjSsxNtYkSF1XKc7YDH6dH3Y
/xHozcXB+jFRJcN73iRalVIiQBdB3T9jmQHR4EQ1UaCITUNlA26czwFI96EqmQojir1T/hWnnDx+
ZJcgENusn45or2ZnFKCpJ6jOjik02I+av/bFfq/Rm81W3g40N4n5ebJlHIjhENWaTNhyB6dqisFo
em20mHSv8hHpJZOtwzNsxxFKoSH81hbIR/TAYS2+QjDOgxNQ7zJwbRWp30I9HyxMt7h9EVMspql5
3bVZ+kZ9/cxTBDbkOH3aO9oO3kxdu3KOL0zYCy3566wXaWt+BI5fsfulMfHG5GJSkTRnpVc2xOTx
bOQHW2yMx0e+IKxzt2VFQg4KNDiUAg/eDunwvrkgo8qCTjp6A1sn6onq5/h6xgoJ1lSzlBgC46Q1
DbJD0mi2S270XKJqpnnMuLFBNag4qzoLWguA/s+BPmvGGncoyiw8XtWgHt1r3MW4ESZn6eq0/Pra
We53vUx6QUCpWARi4+TT/cMdjGLeGX1pCo5+/qSkSdfA+0HIdbCOsNAOtTvENnNjMORVAHJ4NCFp
jYEdhPLaqlcigGvnbLIKHECIcO0NO/vYcz6oTCLNYbaaoPFSm3sd9cYhXpsRIxSnrq1Y0uo6V5N+
oWRsImhwb7ehBLDKi3U/KZwpK+QY92oP6yzZqGEuV3oLf/i0UdVsw11EDAgJy4eock84gZR0h+9h
07x1/0PD/ngCzRsrHQslZ1+LSnEOt/ioSECyZ3HW9qRWpmUNgCsfMWPBIWl+KGgkA2vAsJ1S8W7/
SX+xk4lh0yMBTIZ7Uss7J81RyyCfhoTWFs362xRD2+dmxMvo/gGz1vDhyItQQ7dK2KcvSDtZbbAw
MhuMDa9Rk0sR5gMApktrpKYE5OW4hFAYiyUSYyKErSl0ijG7JfWVYuNUKXgOp8SzCsuBBgFH1TYM
kW+cTt940LFc9obQqaA9YEC7Px1OZu3CzeNvhEMDUrqvi5BECSZ3Mj8SVRBfmiEt87LE0BP/TFFt
m+Z9srXSldus8o/YAxCBNmA3gJfQUX1802y+0fTBWRmh4dhGQdgNZfFFsO+RGaeLCxd+/cVsdhxE
MjEIhOzEccivC0cZl7gIN3ysxAYfSRXcYmMcjXkQJTLFdIgVy0hePQWgz2UAsFb5Eds6tvjg+/pS
q7JH7kWa+nhx9BfrbNvAeOyrOjs25hB/wT/d1TxYpV3Z7DcSzI/B4oOVBMqWRi+s+bff909ndX6u
Y/tpMfqedM29KozQV6kyWDV6V/dbEQnoQv2hrlpPBMRvthEQrPA34RdPHi0RqQkd7thd7VBREUO3
aJ0VVWChtwEC4lUfoUNI+01hKB9AAeNeC2Oow1AdYX9PvkUT4ErgfTt5ZbO/LpBQSJNrYoIKQ8SF
pXTYRALFovM0bsVSTKNourCsRwzIFAUrXM+eOKz5gh/s67d9jrpnC7hb+TwGNKyXqjK3pEmXzua1
G6FMZFz4cGTwrCNLai8zKKbS1ycusDDOcvqepbfTY3OABFiaLUv1T5qHi2TZsIrWj1d8HgAUkFRF
9xxNZTLEZDWsRW3G5E300PuDB4SwX7vlmHbSocouKrRmae5WqehJuSn/uGlZy1A5Rdak6TX2VNGE
VbO/QjsWxw81c+jWnwGbKIxEDqNJdIrI21mymXbnSfx23/1dPfDS6D6YegoMg6sCWLeHDo2guj63
AOrGjZ1VlfW0szo5tNSWZmWE7uOWhVdcSq1Hwqin8gCd5GeNfkAejntCkrcmMR8SL8WmYiFawhf3
Dfc9JCqtvqDGg3KRFTo/pr1cex4M2ER9VZDxOKse9nq2kJOYsjvGgUvg2CoAUkRc1n8/ncidNFzX
yb3TUVYQxWnYROb07gYGv2azu3+cANhQcOi6bMkYtbHUAx1jnvx+JAxJ7rAti1R5Vr1xbQO8P0JI
LbJlZMv/LB8/JCvMjNd+L16txByJxn8/gUrby43/hKHIOrJrWx2QFXlFUrNkgIcyxB/fcBQ05FcT
raJc2Dq0SnhHOeXnfHFqGE1aNepijbHakO4ae7GAdpP2wdu3wlp3MVznYvxbvkjx6fuiMqaRf5G8
3Rm+PIcwSbY6XD7aHGZxwmSb1pLMxj7hmCyf/pCc8ROBppjJYBbDSHXN8xYGOTQDnUJUFtqcqr50
RaBy1jp477FTFJCyBk03NidTQK+LAytEmP2f6kPhr3yw8XgX0Pk7BK1FXhnHX6T+QnLfdPIbdSP8
SVMOCy/YoiNLHUMTraLa0dMY9WLG0vcfSub5+n39qRRk/RBN0+2eDrTOMojtADrFwNBSENR7MWX6
0Z2oKJlJoSMJ2rAPE+QbQ3yRnG5O5mP0FEIKxAV9MRK3hZHFZ2n9J9HogmXvtfswrdXxQXdf0aCT
waEIRyVZUAJw8uHgN81/2EDlyOy4MXLdHkRq04xPVWlLh8odHoMSkjjYrHZ9kq/OTeUE5e59gvBz
EUtRkPi1TtSd/By/WWCjCLUhwCPA8UZg44hPaPyveT8Mr4RBXY51PCCtnefOoMcgdOLzaEEda2Xj
VehctQZ2YWRRWRzb7xQaKFNpowaqKCvwROEMBfUZSWM4OTGxexDrkS3awBpEigqGNlcCoUBMqMdY
bka0xi88ovoaPKdIGbOXWPoWcMBZNZz3Qkp1dwxKA00e51c6E9yE9t/8lF8adKgkeezGP/lpGJyI
CFgbv6e1SgxFR1UXZZ0iY6BAIjFge5Yl8kTc+CPVmncDT7aHZXrhecFBK4zLUuRYAkjYHhO4yoQc
hHAZupWcGl64Ki2Wq65K6cSqob3WKPpIkcRwR4lKnh2WgZgpEl4sv37Lp7F3UBjN0b0Hn8qnLWlR
5l+8Ks3xbTCCRiv5IsJ8yfVqPsh7PPFla526U0NHiyeUU67G1ExZwmCAz0A7q7Pus+2gPK4d2p0P
D9vKSB9xgooCBLQbePdFu3yjMj85htAp6UrmBNDqlb63yEhyB0ms7ZEFAxpI7THwyZYVh9Qbl9aj
mDpzxSzvGn18E7x+nt4vf6K3UqdofqvO8pSH8juJPaTSF1ltIpRdxs8bi6OkncyalJu5geKdL6KD
s5cO9IlNUeBI0ORKEg/TXChM3SCMNYkrmSwWqiQi4+Ch8TYgOeq/l88tcnGoSd1l/xqytzoHe9Dc
YrgdG+0sXBny5eDNWesRuskshAKf/8NAEYaEenS7WTKjHBsKaVeHudbDpEd8nhjz3rPf558/jStA
CuaDoUC6I5ckB4TkCKrIqKc1TUTOGK1yd7Xp0rjfsyW8ldyAZ4m2pHSeBJMaErByH9+u3t6/wvX4
GsEIeqB8Pgm10mw5l8xTxsa3yn6zLUJpY3Kp1s7bKrzhnHkeRYxL6L9q5iMDOlHz8lDd8h5wBNw+
E+yh8hd2zRUQiXXv54+WVqasWQSHsmcFAM6r9fjqUjulfH6icR9WJxuIA7ojpc185ujAOhkOPhWJ
+BvvcdMF8WGz25EFYdbpA+SUiaN35BRfs8uUk5GZ9dtoYFVU0nNCtUTrOWOcNxi4ZBInEjw7q7Zo
Je9M5LvPMXG0+y9J3pzDUYCKoyP18jUU13Igrq24ykorQisc4a9SUNdrfgAh0avUtJ+xCvDKTEcB
T+JvA9iqUkRJRb1vEmBaohCTY2LF3rLw343hJrscUr2BIm7d7zkuyl9bMoUnUPwr10V59YlTZb8u
dDLH4jZnLd9gUMy0h/F1EdZXEV7ivHn7ZPkmhVUuzTLACqzeYu2F5m9xLgjGhkrwRcyAL2dbcBn8
USlnZ42KmFwDbz5WqVv9dCB5bW/HspIGf07KH1SlzC+bJhBzwE20JgPRSmfHjrZQ7VECS6JJvAb4
FX/pqODW2r/VHoeuasBhim2Ogla3QOzVsbJnycKRsAZrjAueYcAtYfKl0Gy3qWDlahJGlzyj0s+P
QcgPas1+mSsti0fF83pE9j2761xHrgwKyO6085+z7iAJ/DBJ42rNQZMzFbsQwCAFrtgJwVrHSZ6Y
pm9iFJAGOtcpZKBUF45TwvTUBlIiBOjGJ4PGKSImwEkniRP79b9wAEU8t8U9+yebwK5oQrOSsr74
h/u6mAzo3qJFpRQOVb3E+ETq/Lwx29QQm9pDergpygkijpr0TKP36uvi+ItC8hK2BIW7gRHhLZri
3dkxKT1sTpDsx53gfI9A6SkYeDSd78nDVYT2aQwoVOWiVb/wBB7/nUgQieGCFYOS95+hCRTu0PMU
YRufmnmVBn0AG08ug/vWFxrMfczWgcO6HA/2MVgbk+8GyLWi7DeXueBu5q8+gD59Xtu+ykHozabv
cxQKXzLFfeqsn2gYS3RvMEnGo8LNot+bO7jM2T68789Nwb7fq5RvfJrqcnho7txjo6BfSeEOH4Hz
bx6ACCCVKuuHddOy42ADw2IyEpL2HhUX4O8rOGc7rcln91tDzyy7BZXKXPeXfi8pLHpRGdK/lTKm
UDEKGnxEHbw91wo4IJOxYPiv62laX55WiueKq/OPc2WZUCYTppgmLeFz4AYIlVP8OohEnffe4vt4
Pkrt3UwyAJfwAR3lTvBG51bVn6ZKZ20FN8SbQlH46FBbgioDpR/f9yoNWsZ+U75Cbg2sVifi3eFj
c297N9RAJkZr0ANKwpqlg1a0QvJIeSDwbA4y4V723IWRSilw5LnCFXrvXvdpEFDoKu4lpoobfNje
Vt9MVsv5OrX9Q+0mztTG9i1IBZLFWER55UStGCED5SFuc4F6h05iWCHOi/O9Yrtgf7B1ZNBkeJpk
xPTgE3H40y1jU1w/hh1cmA8P8BGz9SG3xJAGl3DLOveCKCpStzUqrUcYTBwUkn/Ib1+o/pjX2435
vA1z/D5dXAhBbtjyY0Wge5VbnKWvbrgYRFzIIR75hL6R0aI+ZxXEK4G0TFt6QhnK6Y3a5wXxYnoN
Z8w4fVB8+uEo0fsOlHzOPYQcZw5UF6R5Y4oARefx7mtDseaXdL1keEEp4+Vpy6KTncZrO6RZnDAd
C9KyjO14dCv7DQD4m5kWDZT+Tdq9VQsfXs4L+u++HbOdY1KcejRrmwtKE4r4XZy+nN85p8tkRoJV
q62Czp+fXRP6ShF6Od0vADgqAnSp2nGmYE0R+P7YYukJkSb0lG+WwybsBFr7CQysuyuv4YdiFFlZ
6yldRQeQFmgxZCS0Q1+3IMe9bXdGbBfUGJBsQveKLbPLyjquRtIHcxgKI72PEUc+I8eQ+pjuNzrQ
76wYZ+w6I3BEA9ljjihCa4ZY8MGA5h2erf4DOEzXsnuLO1EZ3f/wy5aJjV9JOiZvJEF4Zx/h8IsB
+hKdcDMqWnEHbca0LXK0pQ/7Z+a7XOiXP/O03UInMfoRPgtMFsUVWajlgs7XSNJqaQ43SB3yYqvr
TlSMnHp1Aq4yA6tqBRD5FIagdYRJ/ZEdhyCO2+Ex3/Pg+YqaKrr0+fCh8P2+EFN71N5XY7YJBk0t
lW1lEUOB39k5Z1HaRtvOz9fJHa2KeYr0Q9dKgwMC+E4+f0Erd4NyMx2Ta0yx2Vj7MQ41NvqteDvF
bqBtAGiStxgklWPmJBZfJ5nL4uj3rkzxVipcdvjtaxLdogGAowvtOD593jBK0yu9mXYLBQ/JAJqy
RTxrr1lu7fqk987uJkN7obxr1HglCX8+nFQNs+S52MSZ8VFL/ue22lj7d+k1x95uI+K7VpFcdAUE
H/eAqOTzSUGCSMa9FTPURFNd3GbcWYprEmqxKwjqHGOrLL3V2+tLhZCm9TZsrH9WPgWfMa1+A3hm
RbO1iJVV42nUEqKGQdLReZuOHAIL+8GJbJPChcu5jf1a7DnVrXAeJFMCgR+zv0DahTNm8kE04kqG
HRO58YVyrt+WkAIro4tSxc0x4Jr3B7/+pwaRpO4Uq6XQOywQT0AmUnbhfnSV41MtOeWWJIVvEXOs
LuWY1gngqkC0HT0QPoJ65VywAyph7ZnwjkER6EUeutS745/EUVxtPK4ailN1Bdn5M5p8adlnLU3v
vAEQyzr5N6Te2E4cUhzZWB0qOpOtq/aZ+khD12eLUgv8Bmgu4zJm6Pnyp2QWu/q2WAWU/nYvMeD+
b2/Q5ThvwfiSME1y7Lcl2Jq2AJwOC9tb77VJ+9mqfF9m4bVyqbusL5QT7jByMv7eqQAyJnFZum5Z
tBat3HtRbjNeqfxwP8pENjDbnpLMo5l1rgBqD1ruk8CiK40HrF1/lblnDRvnq7FWiKoesBkUa7gz
Si+YAobhLAMxhBSQ4HF9GwDLatWF7HXrGoX1xx3RxZ2Rtac4S2AKqBDKjgOWN+Aic6el97rJylqm
wUl6djWu00lsxM78/Sh/SALKBk4l4KZ8nv8GWx3uXhRLtc4Z1LjYRew01Cdq56+h7QQ6o9ZBp8ZF
GsT1cEAfwv4LsxKk9fvZBhjoJol803OiFgzuFnoDZoYOgtbI2OPiQ3KQ7w4yKO5sbRX7B4xrZNLX
XTbKTNGS7zINS+ZGxLAUm2CYYuPXSEsB7HIY/rIO8UHHZpAqxF4PljDVv1U2DwSsfLYabZrkDLC+
QlMWmcWv1ByJu2aWcJZ3XhAmfTfITWBYmrjNHGauFNuceMVGm7Vs9Mu1gipVOmJVkhB5pf45C4BU
pptM0c8zaj3CBua+E9Ei99SYrMNrNPrgDfy8w43UUHnkCFRgiSnDfHpkd/6nTs46MhzmQmZE18qi
OYs74M54KT85qwdi1VYXeOH1Z2+MT121BfBFCmJ889fGmuTs7OPR7T0w5jIooPermGu+eKy8AmGO
3X/gXFFZCJq3E7sIdm7jq0xIgprAjwTMJLfQLpv6vYbWufU0T3OCqXSyUeg/SoC9DQy7UlFqvA58
/aBr3rfphYq8rvh4OlOjCl+GMKm2HZrx+gY3LoTnI8M2I7Kqlt5nkTisiorfC7UkqWpTFCq+CN7e
htf+zJiI8z/Wr/D3fjbuRXRD4RW1B3VzxG02S2m8n6hfvOQ/O2DbdLfWG4g9GSMdDO2ghw/ajtMh
B2xdyUxKA/yds8fn04CxmDrihlyJVkx57k4V2FxqSzSMokEpkZqtaEiitF9Bqml3/h/3Wb+0bQgE
VN+RXN0bF3yMhy0YuhqiML5HRto1oOSFB4SwfBlQw7ZIzlN9EhjvCwKiiqFwGmltwgKMXRQ6W4/w
iSPmeRzZ7fwHLdCcnIlJUIOqNgxS7Ulx4SvxlhrIO2azsEWqOX8QMRT+Hm4/T2NoZQr27dG2DWOs
NSmsPCJzgcH+4XgKi6mJQr+gJoXmxy2M1ZpiykPGUxO2Tr84h6fmY5MCk9zISsjgENmBOj3DoWzn
X1rUOvCxpz/lP5frsMQc5LHM5dsSriWe18rrUDs3ffOrpHdF4QfUEmwQvgI3dpDYlItD0YZHsj6w
cuOLh65osR+TuVshYn9NExtf/P5kyRYt5OYRSEll1x9bBoHqxNMBMlTssvbZPwhag5unM8fypVJh
ZVaYi2HEUGWY1eBJwrEE/ynHDMq1ukFcs7sKp8V3etIjSN3EOwVV/C+jT6+jwJRpnITubKZuIYss
CmHguLHvjI6BgLqZvLuLKC+ftA5bqV7k+RRDS8LNR2zUZKJsYg9M6nFcYOiXj1S96Xvhx1GVM+iM
q1nuOVglHrmS9cRBC+d+otiEE0SHLws1sFX9Av78pwLbBu4x5PviYYCkR/YrFoN54l1DRkjmEsxp
ZRA+5fhKsbrsvubh4GxSZCPXUJEpupsotUx8QzvAnzBVWZh5Qa6JkOVMnifAenBUd+bLKLN6EaPr
Q3C0kDx0XPoBq7m+w2+4c5B8kXqzJxtIFhV7MVkOq5lIQZF2MwDSRSmrD4XBMV6xUcj4MeFB6C9r
jwIiAG+aFLEsimkP7M+iaKnIlNa12NMVUQ2NDsLn29Y40M6tmzCzccpUICPcuA5EG6WVDXwJjg8a
kLQLTo5TjyUL/cMN2aATywRQJogZKdcaPf2RzRAPPCAFKgtJMKP8txqGBRbX1mgP5nb8vd/EtVtk
VKojP4m/H2lSBb97NpPEOiwrmrnTokqyXZHZ0O2QnOrWaNU176rvKoo3MCZBpqSG0rkcyGtQs69U
7c2/174nGLV9Reqi/CQNzfgMRqHgqnqgT6thE0B+yRDa7Rs+9qsmtskZyKA5LUzzRoRXQk2ybvdW
cALkjflYI1abiDC2BZJzgKRdCsrLuW29L485Zgt4dk+/7YGDYgNAxWooBQYwEm968GO8uHWBaxoh
qO539ER/MnIuGGdA6Rc9GQ+LKZdwx5tX/0jWlQZRgNlevt/FxlkK7khh/H1Fd+WS56YhDIAmCoRO
7PDfAW2bzGPVQUhCJ4+k8GqWN6QdDlNy8ADgWPTmHuUOA5gNpYBRQhNnPBDb6JVzJ0EkIt6HEwy0
qfSM4Fj4YB9xsHEQ3RwBoCqWoerI+fWfALUPmfTK8ITPUXDAisFx1Cs5zM4Tm6M+LRybc4v4uc90
PXWVWtB6wAdmKq6Xpip8BaMd4WxJBI2GWLDmju2+5fGELszudev1+s3JQv3mBe5LlcRfTsI8hSX2
7GS1KeLMIzxcJmTxfvSmuCx0ohJoi9E9PSMKonACpHJip0418lyxZhK7e0wtYIqgOGO4liXPqvAk
JsudDwmONi+WdJpmeJVp1RiLswRil/DzCfim1GHZhZNhzE6wf1vWbikGbIVSQ9GSTEosaWnFVLxM
DAhlYmEG/1TMpNw37+VwybRAgg9KUipYxk5MbcXLvAoXGumfS5q+2D1OPk/JPmlaxuct3sNmZZe4
3Oz3y4J+omk6+OhHeB/xHlo/yvAwFEEmOPWZtovCaKqZgMl+QzRUXCirzNYJz+ySjZMIZwYOV5Bo
WP8qobI2xf5eVCsnXnOeAo2FnW591NCyFaXtoHTwhl6wdmG9DUTKGvS37Lw7P/+bc4IoA+fyAeuC
hBs++beHGBhyxkqA7KJ8GFH6d84SQNPQuD316ifBj2AdPt20P3A9ZwPpWdFamrTnS4Jn3tvPohHD
FpVj+f25lTcHC7NecyBa0rQDnaOKlEYOlLCpuPQnDH2ZdICiWLUtLHPSqkhJ5fhFcFgSgVzrEUHK
oDKCd6ZHJeZzn1Ci2GOmU+SyeR4Ud+WSL6hrXwqk9MsVsZHqfoH46uolN3MqbsL1DAVpByfkOIra
fnPXfygtyFrAAYaM5yol8/SPwV4J1ivNJFRQGUPyPoVcTaJhAbzDF8TQxaxXzx+UR5ZDRzdOpi3c
by/qsHBTm027AcWPSEAqXGGOXnl5uD27H1+9oBxW/NSltu/E3suWXJ8GVIg7DAnBDSsdRTvS/rhS
dLzQsW19rGlenDALrMYQP/BBsJJR7XWdZyQ1xl4LUpFJn6edSU1go+MT9phfdvSzdnpC0wzsH+6A
0OR/2GySPpzBUYWMteTMs4eE3kgOQMemHSjqkfU8Yo7Dtd/tX/VBj0q+xVlSmKixUsgBCWcLerV9
bxUTOwN6Vozw5O2lmfHwOED3gov2jrhkD3KX8dPryXYbScMMeHI2btW0VNoPbH7LBHlFo3yHb7n6
Ad9rwvsD0sLSpXq7TntscLT/bA5/yDa9l/NY4ObI2QK0i4G0oQCLFkUIdjjm0+n0+dhYIzQICF6o
b0sJfnEKsaX4cwWEs7PsH6vRzgulrzHel7X03mumF0i15wJo7g/kNL4NGYypxKHTF3bfZHLmfBGh
ADam1NGEV2zehQo65Ns1rKd83mz9awfIveutrdlZiC7ch9//JrKJC7F0TNp/XTz+p3/wS6g/OeJE
BO3BnATWs47kGcPPVQ5USE6r21bYWPO0DuluVRq+frpAWB4AC+ruagF1OjBvFuTk21SQr4SQjVA/
iZIvTkuJ2iSBEWv5VZgP2plDIjpVFJaGGpa/NJ+jpQs5WAAA/isUP4Bc3bxUPL2/HXhp/diauLV3
0EFrDln4XXVTUVXGa2fJYkt5I8E4PBt5UL8shz2pQhH/SyncStnXSJk9Nb9kF3PQF83bKrS0tVeG
yHl9o1JUdAKjQMeSS+awkjWpx7egeHd36JNcihZK7kb0phewW37yeatpwFlveXemxop6xm4vjIdg
YX1Ywg/pwfSO8MVikwj3iNAn3SIWhyp5mMjiJxk5ir8dC9coSK8cWIijXnZArQiu2DHd/nFK8oEH
3pdXkdaTaDsXfivhKkVFaqoskaIVhdxJrbe9bSN9FMS7KSo1YqUlGi1SHJ9jGtFCJYgwmbdsoo0I
pVLscSCc1GHHAjfJQf+JfEkLEF8Bmo+Kwl0h4CbsXWZ+YyCgLoA64WaaueyqBzx19z6MQermpTdb
TRWfEoZgqpwSL9ylIo/uNx4P5eUQCl70xD5DNEMVlxdoY88bCCjMNEm6F6PHBy064wccSvAH306Q
p5d0Ah1eQhuKMb3zeKa7iyVVUWoD51Pg0q671LGfiu/GeVeKVS0NCLo81QYniOIIraKTS1xDFOeS
ei2v9jI+cTKN487pcKOMKseGS+778LNQW81uNbfj8nljaXpTh1vOWlvMIAQfm4Bh6J4YD/V5n6Fp
aI7xQdtmUybBxc/GctiBUOS8eTUcp9LVVtuJP9AhyWciX18K6zeBnC6BB0e9xAxB3nmQ0kBbMjiJ
7nn0Au/fsuiRqHJeVNkzrSsp7f7bLN5yYxjGxRKmVIZLsgCH8/xyCu2tT0oHA/e5FrdSa+9TPEOp
G4wl233+O0EKUTzQjABP24MZaSmnpDB97nlT4VX6geoeUayJK28yTPVRXNUQ9QtVgfVKQU3muKK8
eGS9st4lEB8S8RRV8uPdwadWizeagNRKpVcmiz+ZsqP9lkmOoQX8u32j2HJL+X3Zh7HcqNF53xOi
E4VF3MuioLM0K26LLjlwBxxah61bzwanK0DW8sZbq4DsP5by6gGx92cp1XoOSufFso1c781PlRD4
zvXBuK+0uRPhRatetCO6ytS4UsHKMYTYorf+s22T2QvWsLswmovBXJXlzib5//+LIbCLuQI/YVYM
APJfZrJtHc3j7+khCsnj4hylD3PbyNj97eN0G4R3pX9+4Wf6DDMQk0vBhvKpu+dnfKwzpGSnf92Q
2lFoxRHmUyNlUDr6HoQmc3+i6hzHU09SONy14wfWt+yvDj2ARWqWL4WXr/Get5pWREGa/MDQ+Dwc
1Ch/kaTDyFzcFXOL+/lEK8Et2MEixOBiRNH2XxNFL61sQxMHc6h3SGK0GDUP5sq1KhjUyCTjloh2
QZOE1U2OAIjrhpabfDirk9L5Azj1Z8m0u6kJDs8NocpbdBsLPBOqh0SMYKu769wgOsySgIcqKJT8
Qrhg0IMut21QWpJLH7JQvUmLMR6Qu1lSqg7toP5l29mimdhTQAL7uRVCSjrXKLqm10qQ2BWtSKJk
lkvQjEADfR0TalVSJA7MvtpYKmxo4RaeXetLLrk7hY3bmCRUqVW6k7fvocI5xHTunEtYT0SQkoQ6
7HdjV3NAm/o4UTjgU84RIYefRiS/Mm+BSYDMtQ391XvadnJ7z6T2LFGrbAaAd/B367wtgPY/Rg1Z
DRm3tySxG+bSlUuCfZBRScMkXn8Il+Sd8c6hIZdLnb/TQLTbI9KQ4Td2PzaS20fVp0JPDn6/3PHt
rzAFhI30TpawZpf6/7+FTZa2fPbFktzn70fWXx8IhVMIAu0DI9lZkFNZlwm6E19MmEpsQMyTdOGo
yzgW8fnyClXm+pNuVDAd1w4zjAJ35DU7W33anlmxkM+tVG6XSb7FlKXmi0oEueS4hgRm+P5oIwzi
+9ExM2b2VWKr3EFz2T+nIwmCL253PCbird1imyK02nuvxKyj51LptgliPd0j3t7FGDgkqwKtOGAz
L2sjmc2+BbZwn7wxeEn4MB8ybHdFDRapzFCdQ1k5ms0SViTlNagTj3aSUUvOwQd0xxJJiOhn9PvV
c8JRtOq296W7U2nbdEUA0aS9ERY0dcRyGxCGSnjhRZjA3oA+gPHSmHoOg4lJ8WfTM7B/4s08CgZJ
9Gl4z/cQGC8Pqp+KHjMCWl/U3Jo/ODW35on7F6SV0698tMzCgFnS7GelsDthEnhxTaZ3C+AQY3aH
+zub0QANW1SAVedNSpljEjPyhbXeyw26tgERoJHJqfaQRKNU1hRcfaOXx6EVzvHzGm34JRSTz1CD
b3vHYJQ2CyLlO9hup9oZ8yYTdvxUIzkvY1LH74JE0bfC+U1ekrriDbx2k76IYVHC53f5xTVIJeFm
f3TWLQRS9WpFeGxAGldYH1iySu2V1hZEata5kuo0FoqYakwuqFNE/KK0DvSEL3yRq1n0J1ZNJP2c
tjMx9IJREGYRwGSxauhRXkSoj5v+haZNh6ciMEC6v74Pvu3m3oufyAvQawbTS93f56L4ChBCpQRj
HG5DVXrjxd7vro6jaK+8vq6sucoFB3oNh3Sf2RUBrfOM+Y2BijfCQ7+cYJq1FWElttDCncTnQngB
Bb01tysOA4/IX3Uw1UxeA5eNzGpmfkmJRpYRpSjtlJH6XvRU1clYAXvKeuE8sNjS4pgIWWRBQBbn
nvGIaBg+PehMlzp6c6BujkNoV4foA1MB5P6d1ab16JKJp453/dNFpQhOxfD+gW0pnMzUNSW7kNmW
RTNiTIrq7I9L+P1g62ffCjBiSHvLC+pwQDHHSshuBqpGEkfZwJ81bqDXAz1P6CAyvR9gsM9vrODX
edK/0dujzkGbMynXFXPrrD/oBB1kjsXN3dzhRA10mLmSy3pxQvqJg0NRl2XRV9CIEP5zAD87ujBJ
XieVttSydBkd5S8eNTCexDgSm+wCqihDx1xzD72ejkihm13yvIevj8vsdsah0X3T1RNaDeZTlgTk
4EsKTdbSCrxYMIvjswI9PKB1Cxf+Qb8FXFfco6dRmS1uhDcTqQ7IRlFTb45n/Jqj2X8Evt9SHPS2
pG1yguESjkq38wExkuMLwlGUGjdKtEcRFeoLpCbFf3e3j6BumVyNVxTSm9dQUEbFXbL8xNiMoN6T
Szr4arLHJNS3R4YCUu4LURvxYFg5iavztFGS83XsPBHfb0JF1gs38d85xQ9FQQii9bVkk2FbdZPY
F11KODpMjlo2nIQvCflvFRDXSdjLHx5ZBI8yatQXMYQbdO5yNq/49yYzXbNtlaO4a56VEJPl+Gb8
JPUZb8FMYkQTjEKeGS382RchiMoPgLh9baAzuUFl6HL2WD01DrITLROa4XjeKazTO/Hh6UZynuAF
5ckRUaoPGVjTYRYyF8/C//g7MKj1tWd+7gK+kWEub+DE9SJ0d1Ix3MG2ZKYHo5LBXPKgbVdFd62F
zSzJkzVAsRatUuutrUBNQ6LexuGMwZitM9CJflCVQDxjJKTU0jutRF+/VFgK9ExMF4AQLX81hTj5
OQzVJ4w4j4NZofoPtCJLukf7JxavlGNm7fDrKf663q/zKGK4sWQo8ZbInFH2FWjmbm8aVS1sUC5v
0IEyEo4VG2nwfQwnbAeB4x4hPYt15PSnnFjUmw4qn5juZjzq7m5HTeKJInDFOl+qbIi7kuhM/ylW
NcfGFlC04/Ss+OL2hsK71NAy/URLCwR4UUj/pV0/vcsvjEj2oTHjCkA5EOz5iCEo/X9M3BNhqKqS
VRQSYZRFIkld57MKS5Pw2PBtTEj9h7pME/Nn/AVawPJFXzf3F3HHeDoXFHKwdjW21jVuzpVz3W3n
sk1qb5XLD8l6xRY7Lex6s2bhUAa1OQaEBYvbpQRQODIj1rslMgByCyhPrEiQdWVVDN1vmy7udZFW
/vltAgqCaX/GouFnHxLQA+s68flPEhkrFNsTRnEZDH/KM3YBCvw2ipJKZOb2QmSikjfKEF6SHOsW
Y/pj+J/42CeXkLB+k7ep4XS+EGFYDDiY9Oi8waZvFFOWIL+lGuv4+/CBMkxRvwUUvGVpMcRLQFUF
3eIK62zZo6Ws0omC49/euF4CCLY35QK/eI9oUijLYU6b/dwgtDdkO8SOZ10lOEw0GP07v/xcDpfO
OWUmk1kn66wDQ1F8T6rp8oX4Q6WMYwUqgztEdbrcLjlT03M67Q3tMpUMEMR/kYa6zh26k2dRoAHw
XtTmzIQ/2/KpF5t6B6LyOTfGXq7MajF1Z6KIC92ccrgLkbWT4pNHXAUb0tO33RdqyBXx9xX3iBov
JazVSwtycDjANhyBOPyoMzZlwPiglZ0s0cZgtla45nQTVA8MwOjWW95AyoF89NyPzjsa1gz9dZln
k6s/kAjMfVTY3yb2tTQlpKBrCqH27tQ5q78f/SnKomOZbOoQOjAQtVjjBPrP3Z4TlCtumUVG5bFn
4W187AOh5z9FJgj99Mqq/ZPub0eE9RpMBSA0oUnjM+CgEbBQ/OPolAPa06NEMRQSln1fSJr6YJSn
Sd2+AkWKtMtb+pxjLCBLnomTTFyaKVFYX/1jPXC4X1TnF+TLzdiB/593U+KsUrMEDEWlBUgZYri5
s+NckPul0F16gb0IcAtJqMGg3w2KIugwkOq3wKwx2+rDJhydMq1i//+EyOQP0pXYT9NAlUbm/hcm
h93udZ7mW048/Y6xv8+nq4CtJ99VDbwcVzxb6GGNtjFhOXdoNLd3nTVoXDr8HiSUxNyi7aLM3xOM
BONnJgspPQNrLkO3Qyu7w/5bQdCuKnUoDZrGmMFlRI4lBMopzFf1/xR/EpCwbmIUMEwrkH13Er0q
R88On0S17fe6ez9nagJCbbm4Mxx3/+AYZqrjvH3FuhHG4Vk5rZj29dAfNbJMOKndtqrfFVHS23sv
w2OSx1XdSfRg+VIKiy52tgP6zZXiNjq2nvi11uLZYyM2defHj3NGVTdG+m/4gZBUuqw06hk31udb
LnH46gi4GYTzjoxMnOYOrcjL4R79g+9D+sKiuebDPlK7LAcxeuCjO095V41Wnc0sxnvkK8An9ct5
pKmFycmB5988UMMpPIiRkKsjWJODhUBsiAH99TsNSEG0rZPaTInd8lJeCOPL8lDF8fk4U05GGWbx
/JXfnMC+JfAfQ3FPzoa+XdhxS0ACX5LvmMoIFpvHmCF9ZrU32YTuG8QWR3LvemabKYMQ2FQ0hgWc
Aqyp9dxjSfI8nzpQUmaDGrxJIEKOfQ78u6Wfe4LDFrqzhTreGlxUmRnSPApLvELnH5umeS7HRcGj
acfs1RQwYfqkL3B/IICnUgVgqIEIFh57VCixSY9oMas/UPO3JtGqsjLySJj5bugWWWOalqrQGf6k
0gW6H/QKVlMzKk07DyZv4/Jnrk3p2/6ZAa2ZJc8o1HXxIAO2N75U/fn4Avm/3fKM9KbArK3bmCmx
SfSQ4V4Fb4OD21eqq3WEP46t+hxsFzepNO1zUAMcEH/+UvtAQRtrDJs25vNdXcg6P0gUBpaRneMW
wETV1JQt8XJ3ZNi1i9J+589GBAI5GJxorfK/oORYIoIUacyw1JVJ3Fypgaw5X9qFrlkCREsrHxFn
rxMvJNm7y8UkUQOt6u8z+3FZyitPQwhm6IfHyglqFfdSnNd42ACQoO3tL4+pmc7+muAE5EoK6nKH
qoOQU71W2AH9Xen1jGtFLCKEkKDf0SMhlPDmRNWi4Ijt0lZ+d8LlNNmSGC7X+zqF1zrd3dDE67Sr
SfPbJuHKGgnjQ7pZmks/9sTcmMFPFuhrujU5Moijy6B5V9/9yliuN1ZqkSRvoywHjbCJaBC+gEsP
K4yzl1fCNH70Utwm2XixRJdhcMcUVoEjNVYWX59f3onYQNS6tkKrmnDUNdjkr15xC4cWY49hnq+8
4XX3psdB6pYxpoRVPF1bYMDQQD1jcKHKdltb1pyfExtergr+zhh8DCV7ljaGHZDjQGv4CjTgBGQC
IqdcqA/VzLSlBnsAMQMcE57//waNMHrq6tH2ECNYKC78hxBXwvelpZOuF5rcyJ1+KFH116O9zJ9B
UvIh6QXEmmNpdyOX1zmsGss5o/RCHaUBfaF9ScxiC1kmSITg/yxL83w1dWFhrTmjuCAzFKW9pjYL
Nl/wBIldlWcHlcJzaf+DTnrnMuE9kOrwb6wteHqt2PEtAoLYiWfdRVsTFgB640qYashliUaWN9eR
fVkpi+b0vID+HRfj/oSAuSX2MnmhQJVEtgDtC0K/sEkhALL/Nv/Lcbl+1D+kRPlPq/338N/05aFS
HzJe0rbVyLzSTpCBe0BZ4H8xuUG7RbWiFKl4AQ1OltT0+kGqdwNpj1zRscPll3FoLs4M7Kn1zKkU
97Wij1MorzLkZLsKmpeyyf41BuDMWIF3X7DJih564e08x5g6c4ltRAdimLW3X2JMRcbEg40jzrz7
o1DId/balWMPvTii8VwHkKFZWvRC2kuSQhRc1E97zDpwrdFmpheS05J3xAzdTM2qkkbJQOdaFQz9
aEFJtaKvsyHzkQv/Pf2pFWYkdHNPjTzsG2nmuqZFoavs8PZ/kooU1K3RJ7TchGhvAOTf4NXC6CJO
7Bo7ij1X0EhebvWvkeNESJKPVamkboAS5xAS8y9DmWm+ftFxqzSpwE7b/dj7KDS90IcgZMTWwOXK
IV8xM+STDfjX3al3Z8EL1KWWLR9mK+3ipQyGDv5cLazn3u33Y0OduZ5yhav9jJPJXB7gskBQwKBB
KQXyxf4p4IvH8U8pa3QVaA2rEIptS16RI4lC6rzikGkACtQsGudpZ0qSlreYtNdRK4DxAv+4Xoi2
noSfkyqIIADEDEoMhdKxquVCBC+lMySMK5zX08XqKiKF3Ho2XwUE0ViQvNBbSxBSi5uOEUgrU54q
KCZKWy0PsZQrnOkJppU29iXwL8lixhWCwhP/RJgnZVS+U1kdb6DSf6F8YB77k16rvdrgkQ3WGBYJ
WfvZ9oeW+z9cYcVkYZ0Cz6awXe2ZdYbsyDeweBZOsvmdc0u+EC4PEMUYNL4xZq2wniq5hEyqwZMf
ebpuhCEGDkKpXSY/Rqp0ZHRduOLVIHmSkTgFQdHCxCctGZcuTY/wpUORZ9i4qWCZKP49Ja5RQZYc
wDb7qc6/gHC1ZGeyBdGRVHbG5nZjOttZEimOVIm2w3TOeKvMoIzfrErZ8k/CUxD5QxQet4BLl/HF
a82OEuESzfwvlJ0TWOeQ1NBWycMGZm+1IT2YbfvbNsOM01VJF8/2eeBT49cWEjrNRO7s39G4rzDO
JSsOQy3QUMk50TabRte8hA4arYjySECPFpuZQi0ZFKcfkGrhp3QYLhkXSQ3MGSkTS/Hhesq6VIBp
07Js7OVVNGkLUgVeFgZOQIIWHK0vuHRuZMrJSuOr1nQg+ajbolKOIqAXv49xMPC7e2KPuuMK+MSX
oAyRLn1+4lt46ibdkzutyZ6wSyGNlSLqeZDjxrAZVR8ehtgORR7gViIq71pyyrYZmydLSRaIQtlN
p4ThZjqbI5d+gFzsmJ8H0SFcYCbgE5eHfTH5rYUOBKFa37Bf8/pfMjpPuN+UMKjbrNEj6kDuBRSx
oqFHHWixLUo3+gdd71f3/9Ge/xUDbG7yfYp8ZGNBRDq3daJWsxORZmVjqxs6r/DheoOVYBPqi5DS
sbIsj8TNw202lEM/C0pFY8cCFhI0xuWF7ZooJMwJUYvwS3O/r67sbbugZ5+0Z73iV4gMosSrRFZ/
YWDXAKy1LwFZcps/6yRyuhC9275QDcr605Vj12fck+5WgIoExmTAZKad3Ud1oa+d6xbSyV4BFANp
gNs+h9RLwZe+qRYmwUPsZpO42h1G5rXjzMsuL/ZIEle8tOfWPyzngeNlDflhLx06QpX/wO8+lBMG
MtKnfYN07O8mVxXIcENdQwbRXiU+Lmk/+qLPyHzcgC2pPwrTSOQehsnAp3g04vMhBhhrgy0xfu0r
jLJZD6A6pvMHS5syKe/pkxCtKyHnuaRiAZrTkVJewp6fQ8WHgwH/ChzGBNnrE/P4gY4/2K9RZytK
lITbbrBwKAqOGFWdhsKcxdraDYH9BeIW2VkCbKHzO2EMuYINVDqU7ndTrGxbP3PTUFTQDjhakY9N
MyRBKb9D0BXPeN3c02JKvhUruzDpxtz84oIs4q6ZVWEMdXcgiXvGZ4hAs0TeHosZmPGyGnpD7jlb
KynSc1Fi3j8/6oA0FdACC9vW3upXtBNLmzY8KP1Z5fa08DRLY2iR8RiLWu/mBgVsUfOoky9bcBrH
2m/9/9zxm7k133VOnBcvwCAc/JprdsDML+NVxcND6OLedB3KORwkbXr4dfgTEmGtR6pvddpgLnFa
9PPgbGJISFj+8Tk9NVW2Cwb2Bl5k37Ec0zgfLcFKtnLt8ZBxtPsfSBTVAEU2YqXcN7w8/SKwCQT2
AOv/A0EJeU4/HsN8jvQg6jUxvzEVNCr+RIEQoM4Y0IisVwTJN4KfqU5z5G2KNZYUjAQrJy8F5WuT
/GWh5aSvEv0C9eDoolBann+1e2v4G1R8r6IRHjJJPlzYprmMnvNwMlHbxB1EjEsgXu3v62clQHix
CHmLWAerx6R4YQJIslrs5YMZQ7XnkNiNOiQ/sAqFKeNTSqT+iKVurJWLNW9Hd8IlZUAjwduR+HIW
Wu6Ragrk2zwC0F7+Om1AAAVVHPyUGMzF2+JE1d8wPtPXl+wAQJkE21vNM93cZliDfLR4bD6IydjD
MCdvIY/oNRClmXjsXqMPGcVlWvm8CQtagYFcuyzY8TOR1yEasa+QmEPsMQF0mnLIz5w3gVvircQ5
9Jr8M4xXe7lSKeGhf4Q7wQgB5xwjs0u5hNGZOeDocIgu/YgcIDW4guC424uUSehkLFbLrzYgOgu9
NrbfCDN2JHMWi3+M7C5XFKUdvpuTPvnf+7gpIeZuX01HO3te9ygdYVZRc8U/trLhs4kDxV97/T3F
t/MyZsQqUKnQYqpVNymZn9QMoYMZp7jMvu4rayGeR7HL9tbCdaneQLsJaOuuXmUIAnKVJ6LjP3hV
cSddf4DJVHR8t2rgaFPuVvHJYqdlPIqdbBblVL+00Ni1Xs2mx8Nuy2rQHA5sCqnucM7R+SP7khUd
lWZZS5vm/kmydIDsk/IpJgVgYtzKgCRIg0lT4WBPaDXGp5TarFkgcZW2S+kSLfkVn45+2fwsVeDi
xTmxmc2bt84mY1WDpo//u92fddjFcyNu+gkQh5FBKT9/AQdlImstgnRBYxNi96SyWiSmn12ELsUN
J3htwTjFdQPP7QGi2Pblfc3Wcm9zd98Jtck7yGL0U4gt037AFneEC6FjiiH/Dsr+mMPuohMpVtFQ
2RBMVHbYoBwbARVOsvEvat5XJGez7m3/YwK5x2kzDu6KsHa+2IGIKanNH+93C4ZTTEi4MSyRHyVA
ITnsl0IDaKObU8zt+PqqdvLJAYsMrR30iDWN6bvpc/V5kSt1YuI9cf5dxYI723McD/B7WTbVRPu5
gvOIUGImpaRBSg3wd8vSigNihVbpWV/ZNHHcMqnzHwVdugKphZT/seTj/UPPPMLhHe7ZDUqebAGq
XmR8KEcEnuF96a8sY9pV7Py9jkYKWgFJWyEqIxhYGOdcAGnwGU6tXJ6AC7iEUY6TDYf6IWBZzmzs
qYnsTqnj/sGndwE0ZEvA9pQWhp8xp++DshToGwFQ5nT4+yswV9/8MjGZpyNjsswiy5H99Cy5cRBV
bd2tuo6I1/Pt9rTrTFRai1jNW/XJMMhYCTeA4K+Jl6+Am+Dpp9L8Gq9fzwojx/qZridNaj6hMuAY
fAY332QMK2H90kFj+HjlhEXCXNTR5tT4ryutJifHfHnUwQDf2Wsc3F4dWvVinPK4hUg4v+BFLRoo
89OpQ5QiInT4/xh2cbkIdxzZKHWGxZZL+9kVNPDigFGXIDDqIHDnVFx6Wdj62+0EyNSkXAWaXGsu
i2gVNkWPDMMlAQ8oRBFFT3w8nNaInVr1g4VteRihRDVlpN2P0K32mw1mh5jWaR1k1Q3mjMLUp9KO
5eJeiA51AjZoxIW1MVcemXIsL9uKoKE6vJg/eYGNsEG5KfBWC02UjyzvSJEELPBFDqDEkOc/UZ8L
IrYPXtQk/l0IXO5ucDO4WRNbpGl4rRxZVBs4DGAENGQ/IU+rmjVwpjHKdCRubqzwQ/+2aCsnqZxy
oshe9vSCFufO4nzy+9yPFNynvBsldvYn8FH8WL3jURZv6XH0mO5YuLuViVOTJ4/zV5PHEvO3Xrqt
vfrYtMzqfGadQrgmEe1sp3XvOF7+x8IUYIUJ0NSoAXMTXu631Ga7112rhUYFoBqccdLH25gxNAOH
eEuGr6JafWD6Hy46/slEyqVGKX+Yxavj+NvRt63xUiqRtMYHmxGDRzIdiXSMErZ8HXTIhIKkS68q
IBnvVcuUG6mJHb0gyVCxUV6wpqupEkjGAb0Tq1JQG5ZpPSIPTVF2D/7e+dVczrt2YWluemEZpSxp
aZK0ybB9JuxcsBXAwQxIbzKn9Bc8re1AcbJ5ybIculUU4tBmIdcSize304hXo38lf15qV511OVSR
4V4Z/XU4iE5KzdzMbFOvmQZvyqxrqhKCi6zN+FoL35HnOoRT3PVUcsD4UkRmAbn9QUPd+FEMOvzm
KG06DvQEu+EsECi3mzk0dE/DnkKtON5In9fq8sI5p7wF0bdnIUX26KIu5NwpEEyHOo8DdJ5sEFBX
0rFjWrF8VmUhfuiFgDps2YSr94gLLQTE8nBMBY+qPWcJKU5OOEqfUgKbAkAPvSM7a9ixoT/PXIiU
h/5o7fm3gySsX2RnVZvahCDgUzGRy9cKoGjDGK2EAIPp9EstoK+fEyZfzqk9V91Wpi4yJMLwGsWs
KTj8QCVysgLCYbbPRrSRZeb7e7P7VhTkMJ8gnHwLFn9C45ryJAaPsPLXfyhu5Ay0U7XiIbAMU/XA
XCjHBClLm16cc1HmVX0kKLtPbH2phbhN7j3O6tefhhQWxoIYqO1hfse7K2hvvUGr8NFc64Suut+f
h2Ltu5O4o2buJnEENjCeWQT5z0TBgzm5Z6Od/gZ7K5CM1YHAzYOEQahe8Bs6Kb22Bqu8+gPGTbDl
UJRa5khunNhJJIQ/ktnP77fIknEXJCjsnyTYDxYOYm7OQqx32eW0eiYaxMqCYuGkcK4sbVkd1fJA
q5pnCjDsZEovWf8kqMVyVETEYoed3LyszbVHtQkgP1ZeFJ7dff7NoLCRL0Zi/ppD7JvBIcTZO7PX
rPGOHlnF8cMqT0JXyoXf+JbcXJu8VYfXNEknfNWSbzpty87UetGg/t/fKTE4hyMmFeIfoY02Sqvi
IHZWs7Rb265Hn35c5z0Zsx6SLiyBU+ilz0WgPiMDZOq4IMH4ebH5irzOBWTSeRLa0di6IHgVe0Pm
UDimre5Z/FQ3L+8a4fzyX12ujyymJ4a6MlEXdLUBV30/J6I/20VmgwN/kzsYX0a6hy680gIbn+wb
AephsplFB6LyhAc7O8kR5ezowVxr6To3fN+85yUuQKt0KEcIwRHKK42RvBnSBVV5TUYzj2jI/5mR
2lO72AuepdfI/4VIrpd+tWA23GD5kFyHgwbpB/joZqOmETJgsUWjLrPewYyUs/jh10HTE8Hd7Omo
59EeKvbo5uNCkBDoRKEvndsdaq2sxfFCdu+3LI2lInw6glRwHH08lb88HL89F4eKSDQEIjj3VZDY
xOLcvGyozIUpFZhxwcuWyZO/l4WyiJABvYrrA2UqwqVhOIkJBBF1wFP9pqFeqpl9Mj1tuSXfCsCq
1Js+aAIfHJZHvsT66FTLeODCzA5jwKeIVWe9vSA69xLAZcHcrY0Y14j5W3nNtUUnjVJ+yvTWjPwb
1qop/tyREGYkxLX6FFEHLzDB8b0ktTkhP/5euRMGSsKrK04+HANRvc2euA/SeVXZx+Hu287Z5LXa
PPO+wbDYlYU9sQTyR33quqOGFK0hBi+e/0Rotisoi/bFoCDXIlZ9PnNghuJZjGrbfbv3t/lrU2TT
+3ikXGR2gmygs0IWsffFK/3UL+uynHnOaTVvW7b5K7qrRBInNuMa/gukM95OPETCjyMYXe+h/i8Z
vvMY3GUqnGV83eni63Bj5SywS6h0w389A/0nd76b98hseTmC5beIJqhGTG6Z1nK2VgCV5OoK8sey
jdXN4rJ8GkXp97KtrTSQYENERWBCB129L/gH0InWzI1SmsVMUZlAN29SZL+TKDyrLW0sf25GKRKD
4hoeca/kqcrwJLS5nRfqXOARLF1JxzaEgmmpP3RnmxJkA+XDa0qCPLg/EbS9tY5+aTx50/8MS1Hw
qPWJfUJsqPLYvQ6v4DwGzI6f9rK5M8v6Ts6Ui5wgLnX2Baaw2g3MBAh99v5II02+3Nl1330xs+Lz
SPs+IM4IWE1ar1VejLB86+i5U6qo8vByhxsEZkg+zAJFxmJ7bXyPfeSPnWD3J3XjRKAMIEXWuW+s
LHnfqHwcWXjlT++91LSy/H8uW1ABcV8YZx1N5lQhn1OxdzHn5jKlC1x9O8JPKDw6I6PV4jY8k7O8
lf3Ho4eRgOUk44tHzw+uZU2SsGp+2n1Hrw3fd8xAkceJCpcZZ5uGgqUokHFQedH+zOY57iRGhkuQ
VUfIhxs2IszMpCEvcvM4djLmIbwI8WhfI9IALS9iW6wggeahyU3bnv90KUZkGxYhWvbFaIgoJdPU
PHkxrgwHMLofjqpCXoVEldkYDN0Bwiyml7EuRK4FlhxwD/uIYtN9XL+DVRAtPGt3eurO1MZkS5J3
dGw4cz/JNtl6jrLUFizb+/XJDNUINM9Wx4HgwT/neokt9WAGPaMZ9t+UMY79gZbzNSIZ/67GWtRI
4gS9K39zT67hJXKnxkhPzUttHmlzr5ceDTzRXydoWfPfD3SqfK4m9giu6J7ZGxtolO5qq+tlJNju
pQqzLzJ/24ZX1m5SFovhZ/jZiLOhSLAZLP+at8Bkgnb6vl7lKty4W5ca+Vg2ifJYXvPlXOvncifi
ga9fHiZkn1FVCO1Nuzs7KGFDUtytyobgm1vt7QeVl2vJh0oI/Rq6gzZHS9Y09HizZPClS8ns6n0l
hdAi8fTfqqlhPjRohnp8kKreYvqU1Gl9FEs/4Vi1NcC5VLqUQTZzzRtXrlbMvpMIJXUMooSW1Kvt
mOiajZEnfcpPHltZZJdwB6o7r2Woc2/O1YAmTtUtrdycYNibu1iG1rLDGV50bfDx4xS+JL27omCK
66wbzgK566k87Ewt90p8QrvzKyLYVD4q46+nY9g9Trjtst4rOglFf6hyO0BzmiKHEdxa2tgZ/9dC
X0SKfGv9izU4A2Kz+eL6EZ2zp1uVTELUNH2rJbAmwAoNlvLZfV8J7cCt8ZfuH0VwQ3gQ95qPozpD
EvcvizJ2Tos7teOS/RqiH2a8kq5tTnCP+CZk/M9fr1zh0GqLGKD0zkwHj9ghmrfvCVTjIUVAdQwW
mh1rLqaeLEzGCluGY3X6RO0bVHm2mhBuNYBXvaMmjTfioWgUeqyIdGGTACGlphvbCDmFWySo1UXo
H/HXmguHFrQGsGZoUDFBfa5kMUxwQzVmLaNT6fh2CN5oy7Dw6hI83JBVUr0QTEf0CmPTWvzjzcm5
ENRlQmQ4CIwFQVNSzPJp83L4Drya/6B4zabY0lzVbJgsH7lVn3VfMbFyw7y+KK+vCrrVRUNd1PoS
WpqNay5YwAlveVl71R9Zalt9ORKR/yGNinPD8ZxgkNFUfOMgWQ7ZHgfri5lQhprW9jcMe8h7U29u
qh4uQprOIcHegnRN6a1ZXURzeO21m5uPPh2eQte8zBj56ydY10VxowPM4wZJ0psZVbOdK+0emx4R
P+Pfu1Giyp4j75m6+KBKAJgoSbYHTVT0P8vYG5JGeilHyKtwrrpDzdlNdrFBNAuMTT6ygEj41MOd
2IXzKcBxODWRApvPqgWPcKMddRniECkzDIPsW6T6DIOR5TM9MiP47mZkTn2cZ4rmgtT8e0TtD+Wr
TxFo4PrasJn9aopVRePOhva+8MCuxsa1KkpqVUzYFB74MeajB6AjDl56TXefBjSeaLHLh0DWJqOk
gG4OhgKYEKb/L56vEtmI5I6zKfJRjTXgizSDTIam3gVn1k8jHxwgJPhc4UQZT7ZtzN8swjFZPyVW
r8SdWWG3dwPWifHcYT7a1wH0z0lX+I79RR9HGJBsn47eNL/vIZiLYxl3V3W217mKrSBJCbJaEDo7
Vt9K6nFYfblejMScvmhCj8vuALU3IaKPE+n5zyNxHv/5HFvSqusZPAE2LsL+kd0L1CdoBcDXKkxG
Isa8Slx3/woOn+2R6oe3IoxhGJxou8Q9wuLZ7/JuXv5LR4Jd9MLDcmAuFrEwW/28onOCGUoH/1Be
b+N+VD2qnfwpgOpDZB8bOlKGp/B7Pf0rKrOfxyQfqZUP0EekBOuczuhcL968DhfyjP629SWV1ydE
tR2y/M777o5RRcwU39eGHFeNqurMIwDb1Y1e0dYD5kQL8qm+9trLvw5Eja0kxRfSPUcowuGNSGz2
yFCA5eVsPJ8WzN0L8DJfVUv0n/xcacrn/Q4Q4G9nLLTo9+0edcQcZP5j4tvGwJzQnEC9S0FthUps
zcnZBZa6SYS2+Un10KzOQ/j12xjoCduEo8bq0unwwR1GtrtJVZPj1LIZMRIDgc2Oqm6g1ozT3Sli
QXz/c9QnjlU8ab5zsD7Wd+/TLwdNY2AuMawHaWq3WNGQn3lCWf3rrFo/sgQ9kHeWuf6Yxfnnpfo8
31CCNWa39OO85ce3sm61FTLkpkhd8aHB43vFJm0hYPMNIReKsgEK8l3jSlTYY5CrjmQsZbn7JJgp
N/xkEeQALVfQl1drPnmWWglOgPbAP8HoX2thNWgNW+vk4uUz888QVJqayVWPy1ibYt+engFwGcar
3+acLJUIpQwdpbTu4TwEbEqeLLIf24/cHf+VMW7aNm4L4P8EHaH9g/k82YNCJ0XbWmm+VpIhiiJB
654Ox0baA0yc+p1Q81Pr2NDNsJ8pzoZre95UV4WZytgZ00BbaOCbs7zYQAgTakPhgUpXGjUrNw33
H2OUltOzC1Kn1JdsMcqU3AIsvP9cjDo0m27zH/9kwG8tDerDzVq9wXlJN5W1tydetIYg+RCniAv9
D+T8Y18brEH9oRV3TPiEDLBDDBMs9ASsQdin4kOBuDV9aOEYFaxBkWZSYc1GTP/epm0zQUbIY7dM
1T8UhF1jfNb5B3COp8QGx0eJNLx9Wyr7/a/KLEl85YiruO+0H11VdFiGiIp21qxPqWCPUdreFOjK
EZqskgBo625f3KTrZR0NfwuW8vo5wJd/8AdZBr5LGsZwYq2hQdXpr6b35YatE+5xRfkauK+OcgxE
zVBFRAOZZu3b81kOB+ngCta1B0WxWvjcO5eSUUPKVbzkojT4gKXD8W0rTpxfYY+6IxE6KfAPiM/1
UEXpwXSVj0FAJ9AgKGuRTN31VYWlA7eA9C0RPf4CAuI+7dh9nd+Csj6eJ9Rr1SMrfiX7oLLqTjA2
ALjrneqozdatiCOMnfkOV8JKR5KkI7gtpR3kDxsxV6tSXSr2+DdRcueRDtJ6wMklzGxpxqDXo6R+
jqfkkM7C4PFH4z2I4sxpouV4PFjab+f8gxGSL/eVU9+QXSOBcV4vsCnAi1JAMz9FaXa0DyBDbqXs
MaSxFSEIClQOgWHM+l3I0hTAHSkIDf37fZojvFm0kbNXV51izIwrND4/pwsHZwbWgecryWksW+Vt
LOLvZkLRde6u21E7Vw9DLR6RaJMSXzsO358l9QbC66wxdO5lRpeUif5AegncqdzpQGjkz+QY3BsF
JHYiAeYvd6Bq/GId2pzQUQA4cP3ORxciDJwo74D9ntQJdnQryKtlHnTrDSYrto7X8RX6Jgg9JGZs
rPwmN0DYQvImNDEYd+Yxp8t1YE/JPXx4s+b7ON4C7l6VO+m2h2nvRBjzysdLdLuwxoGPN1KQc9Mk
uoUK1W8Zlveh5AP/beFKY7j/bNBaIkU8B9kGj4Dfj9tsVgmZAkQqXRuwoTmwBPFFV60tF1z29i6M
OHmXkE6lmkzdmE3wPFtCXn28TqeLpulFdmIUjD9WUApaHskzYiZAJhYP0wYK+xdWif5JfciBxXTI
fWGmRU2eZb1WYIkl4+ECPkHMynorVISZ7YHp1G31jrZfgT0dfJdeXEzi9TYTIO79SP3s2LprNNRC
oJ0VGGixHAYL6iZ1YZH8C61OvDSFCk7mVZllk4bwpZoxwnARgWy/7w8DXa4FR3U8gbfpgwJ3Zfpb
UFZ67RUHrXv+46/cN0xE6Eq2s+5OYGLrd98Zg0E6fWZXIDLfIkOPEkXsxx7T514phzLzOdJ34tp7
12rgzwFtujdteb9f64eAMSzcK9B29Qq17+bd4SAHvyHn9+i7OYSdRVOyVzk9kXWvQ0AWAmwrgaEd
qzsUfZ9FcdoaFCQXMWSvCJReI0sh/L4V5HCPASt9hKRsXUWvL0oIAHCqY97rG2G1Frc3AsJha+KX
S52uMLjHIvc9+FZjQnX4p/4i11X6jVBX7YiaI05dfD8jUCKTqDJwkFhlV2ChjzUTr6ijRNVhtMeB
QJwORL4GMPvHbjGTpjDweDFHvPxAre21PZ8OZ5RCg8z4oWmMDZ3Ym8OM7H7uS3cj1KbP2MJWuLNe
QCX9qpamR1XcC53U7FzWoaooxl1gxKE6C3B/sOS1e4o1IXexmSA3usqp2W7px4K3o3DHYpyG8+Gj
b1DvGzCoij3cU1dnP1OAnCEIAan/bDKPILIDBH7ELJOHdQlToJL1ijUjhVQtfWtRxFNFxFTpq9wd
f+1vWJ2cJ9GVN/OcgnyIO/ut2fuqgjopiOoMxZGdnicG59cs5mvURbTqtzdRzedfnBDXbl4P/pCv
6ZLn8+xZlM9mk4TjP7k+ddKWHynojCkTwm0OBHlCq5oqmg8b1kJz8ZtmthiT2xOl0o2HoifbrTCR
NDlR4FLe6q13EnxR3+pkuxvuzOzfg2mdDb0oPVqZ4TmxPf1viQTTguAJTQi8+hX4OK68aW3bGcm0
MREEFmFyRye5Qe9hfqYwrf4JXgYz32DsBUfpJbaQc0VzgGdupMXTFvjfESSlJnRffJh3gqoWpl6/
Id+Z9VpiXwtfXpI0rRTytuSGdXWETBZ0Zs7lQtRI6rwA6pcQdOCdFtUSnHXMR/55uUDO67o5Un6r
jD6YsohtijEgQqor5FSv8XBQ71HmxJMjiOLsHLH25N0DbvaOIlRA5ZxReSijQNtvB/65+29H0p0c
X65pZ/zYtz5OO3QAAhWgibtdxka9PsKZw/VhR+a51QNpKE6yr/gPqd8PxV2chcaA8JIl9/mtaRGz
ATfseKBlGftPsVIoiUknhQFJ6hwJEhSYqXPSrY/ogpAQev1MiWOIxKBCl8cRLmJvNranf5Fq2vIl
1d5uz5rFFlxgtEZ9kG59cN34ncszXYy9G72bEy2f3nGaAfusLNqbwIzGSFXak+gWDBcqS0IeK1kH
4WsY6C+5poHR/hWbD1JRw6Kma2WP2/+qYFSp+hufaz7Ao6G2iad+W/Gf/t8783WWCZuNp6HFUCBm
QtYEptRHgN/jeyiyvvAuXZqknmicOaZnCUQKYkc9FyHgVlFxrnFvQRpOA5b+boldT9gKzB4iPoUW
mninnc/fLmIGM7D8wQ41qy255KbdwlgT2QGxIHyRBgQRl/p5REySOrmtBvV/RnyU8Ppx6h1zRpOg
kiZ1g+LDNf8SAb4R5CaH1uGHxip52GSrKWC+T+m3FWcr9qipWzIvIdirRh5mKYBo1i4cEP/uwTl3
P0xsmFKBehjZR2hAgnToNmIM8+lNC0I396gVVpQHzZbd8WRQThhSLllV/OI6F10YdF5rICF94zO0
qfMAGzi73fhaOlxTC3qaqP9l1O+PX1QjOd1iHS6AGAWDUEaS4z0vgxfLBRe5GJ+YxRLHYidnUvcP
ZeIcEq/U0uQcQBL3/d0vy+vPorqJARrmdvRN3Ha4jYefhTUQtRAV73rknv5M/VDVJMg8taFUzoHo
N9E7YeIP+vsop+IHYGNuj5s4KUc5XTpC0MQr/pErS1IhZvEbpZxnrLNWBUA0lqCJSwYhCcrHCi7v
Nkp7czHoEG9v62/yzsOyYRgPmN3LvHxztdnwR3AloJNxHS5RH2HBGvxiIxL/2wWknoWblH19jvM9
gaJCAC2M5WMqICk+uUnoqAsLZZseCLK9gVnOsOizqDU5T6meEmd6dlKgWXe0ER1QhQdfgnHTeJxc
CMEmFIYXKo/xg4ULMbhL+ynQiAfzh1ouDNhtLD0W4IDzGtHepHx2sUE3NBX2REhVci2VuA3WIqzc
5dg9OmpXoYLZFX3+aAat1vAgnfWc/kam5m8GCAW0/JIkuTQO/CgZQWFUUYRNEm7JPiCYTC9i9Cjp
AwAYR1WlbN0Gl2eJ/z1Xc2UifdwvOc9AyqC4XgnZ1NNti5AxLqv4FOwCS10ig65zW5V7WCjBWMEF
TD9XvXORDrbRmCDUOiojqH/LsVHmOU6sthNHML/R7J4IgenGqFoErcVUg1ANGon71Mli/zImQ8A3
uvg4xHn8oJSYOSWVru/YOxxWP3yakiOwdZbbCfyTWaF6QosOXzOdhDEcOSS+uHbmM9zCkWZuQt6P
YywUKqAYlny10rgWgaAahQeqvIOji13NLDDKYUgJc81nACEZ5ION0/+gQXl4u40N23zBTmTFeByA
B8TI8zhCtiUflPgEyeO9f9Zo76w6hlV49xgocbafD6SZFeL38WE14rmeDAI5CouwjdBZKN+KmFzy
zEjpQPspIlxPULtTUFfhm+XsD8y11vZSlziQQEnhPWWQRAeqXEhaAdVZ0bU9Jr4sci5By62vidb5
Bv3tf6uMFRe7vgSr8Of163PPVkOZKfz5aapJxQEEWrj79PVGKF4AULKKWuzc4zobL1MDTh5009Oy
rPDRjwSWLJ2uGniZy+CvqitzodvYgG/X9KHzsUto+afOjdbYASktRqWG8ew1qj6kfzCin19RJR3h
elI0g2PybBpsp+Re621zHVeFcyKmJAOi6UZxNigFG0awwxZUzIqTkPYiUPd5WlPiSIEjU/mo71ln
TZvH3CUMK0mhkoMxn90WQMopFip17VAoX72CLv+syXoCwTSjHO6MscqOSfE73N6uWE/xnufJIVuD
X+LR9prcW9J63ulb2Okr2olBtVLUpNJoU/FVf7WL6Vz57/3wcOIfDY1hpuLyrSjj4ZSdy5qNUyiz
NbaktFVU4GBq/rtqEbVZXGtLYZrViP54SkLMZkK5/OTqsx2+MQOvHc2C9DLCzFniLqhvlEO2s3iQ
Lt6eEQY7WAiVaQdPMJ7Q7xG6MWoG2priJWkmL7iRPvkEGLqNBIGF0B08BtiFrJBoNMkwmK/Cl0lq
cG3r9IKk2BQxnqxJOx9dBuasWiVmWMrAlIwYUKMHlz6lKrtidByWKhW1amZzrpfI8hx0bsHZSQCd
ynElhqlBNzSL/1SRWpcuJcY2rvtJyille0zYcT6Pe+B1wv8vU6nJQjaXPPcNqqrJiNt3in0YzHn3
b/OLBiv56kj40NP+5hN3z+9leePt7dFuYNxFJn2Twz2CYNLR41gCAy1CMKh5GxNY4U1ckT6cp0UH
C+4nsJYsNffJOr7jENsIwQbmBy8Phz4Q+/OdefwVc87fXK3XEPz/AtgMpsIFUV3txi4W20/mx960
26ZFktBcrPCsM/+w0nlPjCMisRIOg1S5ciBzqAYOuYRYVOOgZ+XaKFJNpgNYArunE5ki8GSWrcQh
vt2kKzAvIkgmauc95fL/OZZOrDbKws/zX1hsGK3EJDdj7g4aUCL5r8CrXEHja752EbgCL1vRmbtS
nhH4HS8ROhLL7hsbsdIMwfRGHlguyItDew7YLjEElK9lYAUX9e4J4EBDlZdzWYUp9saDN4txEaSA
JKK51tbBI/HEpk/2sp+nwuMDtiDIKoZMN/cuQyNRF6/bx6AHCNs8E5e+Oo6vOcX3yL5CDNV3GS0m
sVb5UsDS5znikxPgb6iIOaTG42q7A+cW7trK9bceZJSmloty0sXNUGACgGM7yuAEPABDo2oKghv2
HCtf7wXAEiGnrapxvFViiWkWXZZTaHLayeOUaN6+pHZ80DHsDaHqjU3W2ShYxg6MLIhzAqvkZck2
uzfzsc/LEct46K2xBTLMJxQfllbny7a/vE6SW/VcXNqpKVDR7NeZNKpw0UhbXk+NbWCrv1KO1Mkm
dHaCytniOQ8PDGXMmlBSZeBwr7UIrjtGTdMnaK6j7Ab2xwAyEcj1rvtIhfcOsMZyYWyIMyPATKuI
lOhWqizXYgyGWvLZLwSxRqIpb4rK3fRKxaIim9KDw6gEkOIoIwcyM2McHP1np8ZiwoHAStmLsXYc
I6s6EQp9V+i9EOV49DIHZk0K235xBW5GDjtnt+y/+bZ1/g0zDzzOKmhJj0uNJdHspArM8DlH3kuo
nJclALH5ujPNJP4ap/ksOFviHolYi5Qjvhel+YRhRAgDrMdg52HTJ/fS6QBVREg0srUmEJBQI/uZ
suD0ZJ3U2k4YG56OSDpqnmeqsPDX6VQura4espFfIyQSPbiAf62iZYyVTfkGRguF0tSj7Jgn2+bS
5G0VSqbr8k/KLypFFzQRBFwF2wgGYIX8XvcjrRQvX9yxp/sxnTOUywWBFYwMbbJpu4BhvUmFc03g
+EFgU8vIvf8AIy+vXjzIMw05nYsQ0xM1qq8WQjoon8L/d8fz98jutfs5jcfphs1vwkUkI1LD7N2N
tZ49KqPiMdXo5BcRIxouVAuM3/PYFpSNFK0kzYEpwUqKp+ROVqmG5ZWESeYQTwyjJNXWdfL2aC+j
A8YtmlUk1UdW+ciLgfNVkDQvEpEzrwLtrTEd5lttJq7HR+6Q24JycBEvAoKTRvRlQ3TDK4DHef2F
HjqOQhpjfmcI0rgVY1GvyalXv+4AwIdBCfy0AxnSorE1FcYUUn6ilmWUNjR8/XHHmFEg8i9dId68
roOpudQ1uCDK/G++fe9CTSpb/LorkbIq2MR3i+98eyCDLniAlOdCsINBT0pxu1DbdlRd2LJgBMs1
bWh5rxtnO2Irjn1xNgqsUBvKi84CoMoXG/2WaR9MRQq6xueh7TuIWrO6x7zU/IDdkBHpfsIe7+Gp
xwvDIFdDu0liui4HqYe8aB35tfsQT8NaRB9dD0r7jskmPp3TdrvIAi+Ll5RnFny24a5gCC4fJ6lk
7LZoFAN4sS/FDJHZvM31SME3bEAvqR/JYso6LGc4UKYo/OgC1IgLOoQYikm6w8p+hGmTXyW7R3Da
lu9A4QYzeuiDPc2sAHvTYSKl6a9uaGXK2FWjuMfeWvRqaaWE5YCfDpBU1m7YMWRGHYJeF+uxjvGE
/DtAR0bHs5maCadQ19cpLwVCD5MWAURO686kP5YYGlKkuclpu4FUWcQm3sRCmg718zfOUIeNJ7hy
d9C2RtLZpCarCoe54z1IiRZJvVhn+EmdCEAmRMMu4TDiB0NiEIMsHB5LW7VrkC4cY7TTz8rylhUa
Rnk6YhU3pZtiSkqSsdfrkcA7uaEUTb0bSL6A3j5g5Ys5L7K/f/A26GAprgvYzU0gbrPEvG6V6Xkq
w/cnjP8c4YEmoG6YST4AnwMSKw5XoUvLeXB54EHAXfukDgUBnM5iYdluEG/J2LJHmkXMIj9jvTcg
n+mDVt/b6kbr+jcw57TukMyJl7f8v6Wkqrt/bOO0bkDiM5oKaei1irz66UEXBZ+8T2Kou9gw3ckZ
tmTztEiARfazdQ5Fe9+OCkZtkIucjHSIWiQ7yO/eLszmjM7bpqXPS/DjejtNeXx63QfMXk0YOETM
bpsB/rMl224O06+Uz2juGagmOwxQk3+x04OOIK9zpSuKu+49JDfOf4km4vCWW34jD7rhQliHtzAn
sPWZ0TMEAr17vj0prKbe2pkl/F019G/jme7ezRoKpAObmPlCUZYIs2spw9sOkiU0OqSD+LH0n517
+aWfrhkmEehgrVKeQ7rZY9slB/6coqgjF8X33QEdE9ULQ40yUQtjJPSIRjlUmg7KADpKl0xwInHS
6tt/hdJKNUNvjYQgowQyxjv49aHWuvNnxOWu9xU4Vo/PAwZ4szTgto2E3skFYU77Sf2Uvzw0rqjT
+Pbd4m27CpYh1i0n/nMBqGlyufb74eRB3tDZzleQ1eDL+VCPnFvVtlK7L9sCMrdwLEJBWMh/KLDv
JoX0JL64+7vDc5SHdramKkts4c7HUDS74MmQMhKovd1VldvKVz62QNiBRhxKAri3twstjvtvc9RT
FmMOUJLq53arkaF3K5h2jdGJL/fakQMlAl662oSPhSBn6sie3W3jJFDken8CdlUPIxea1d9WZB01
5lo42cLkT7/c0TtorvvH/qjaR1vkpZjPd0gQFKGBIP3k2vHgE1tY3lj+lP0Gl0TjRk9enRuud+vb
AyEJc61v6MMhTx0xca2aeU/IWEeDiqoUmp2/KkfQGSN6tna8dChxFydpC/6XD/A7grNkkYOWrI9m
q1wrKfyCg2rVuVK5mmO2uTjzbJTi5ApKCyoPLRnqE/SAK63PX5DJpgOf6L9mSTvI1CQjzkQZpPc4
E/HneOgecnAyfaQYbhqD8ictKlUewEDMSG1qbMi9urvbvJGI43loN5wbF5aRc5YSmkeD31A4SJq2
1A6wzo17LwmozO+0JRvlskDWxaj1/dvP/RwhewsGHzrpwtogdFEk0q8ir2AQegX5xLVuAT5C9xb9
uU4l6wTz1KLNu7rb+A932MGLTqRHZ4Ifg3nfOb1r86aehwBG3fZXjIKxyUHCW++Kk7x1DDFid1yB
gakivAVmHYwe2WB6Me/Wbm2kE7mlx+cmHamMMes9M7Ps6NMCYsqcryDQUElQEdFHqreAWYFua7/z
xLVeyh82ln8NKgsOezYA7DUA8prPPGa1VHcbXA2Ed5qnW8QEALaixrsNZucTSI4qnJr9M6VBEI3p
dkVxxb/Ff573aUkv9UIlE+1toW8G56DYisHuEvkA2aEqzDynmiXP5hDkdFax7tDrzmgSIWaczMKL
WDL8ECRf1QEcHzhzzOp/4hml44koY/0OyPHueD/gubgmwY2yEWcK+Fv4Ii/RYG26+k/9xgfjN/HA
F18llWxBaGUn5hpxj48o4lRjbC/vlEsiWV9dLUN7IkH3Ru0vA6Ku6lMBAmjFQXe1kpckxOcF1/8/
0aBBO69W6elw23cxV6/DDapJrCx8SEq7/2sLSNuL9WLM15Y+PRLYlTPJkZOXUCyKdRA0WiA2Xn48
sAQTA94q1k98lkzKAqcJwM/807rhNblWudlN/7ohZM/FWVG210yQC1KdhgP1EzaeN4lLMPPagEky
wRYuCJfLflB10H6t0p1ah1XuBEfkNgmeF8Ub+DRbZFnHMV1XNGZb5XAbyAjWb6gVe5G0z2NHv9H7
GkcDTQfMd5xziNO/jqtLxJX44VSjoLxLaIRyApJ3Ju1cs2fInJ1Y21bzXAl9ZRkEvF6l9tI2wa/4
4uMD9BcoOTq/JyONSRFFZf4srliyKx3NnZ073snv8ZjDC4/NmNN/airPAGSUdt+m3yq9z2zlhaKn
5BFtFFaCC3DyRq9ViZz1cR1GYEVFGauP3fwnjJQULgOBg0XcxCcL9ABIqCsWdlNS6s4imY3Bcs8l
zMxoYIPzletXUUo2hjO79gCI77O3V+p59JVxdVhGEnbyH96JpKbVWgjvLX3M5PzNToCpzzD079g4
+/vqsppfkLZfQ8NbINp6Hc2N5mhG/Ap0Mcv2xDdE+52MDSsh1FzcJAb3LnT8+C6eWP2g6dWc5DPb
dIC3OHGTkpVxvxtWlxD441EVxGatRtE9PB0o/lXiw/ucNo8qgecwDTUlUdoiL5o3yopjG5NYDdyG
THbyVWBPR+f4nB15Pm2Xlb3tY7qhbYsMsiVRPr7nGC674GqnjSKik93st9Q/vyTZlgQP8Rucxt3E
fCyWcazt/x3Ie9W601+bIaL+RWQDFrnesr3gnEhkGfvFp/S1MaObNWSu64K2g6dEjilEmUHwClZ0
X/iwZmLNGHW1ePRzlTKycuJeV2zHIbMZPGiuj8skY2nsHOnBqe0bC+7jwDmbKS34sfldy7uMCm7O
9qxzMKkxZxa7xEgCwIITFX6Q/Y4G0R4kPd4iX050lt15lhzSxxXNcEMgVtQsgxc2QQJSD9jzP9R/
dQ2DF8Lm2GDZI8/ebfrX0nDwpLcbBk+Y9Y3XJgpmL1LlSHJ2hBu+4rwHMVPtpB2ULSb35f4Ijxq6
2Q1jp92nyBifl50klLCfjGcnQ2JmVYN9M9PbNyAV2OsyunT06zuxObmfXN2PWhyajVE8iNUZjyb7
PUNu2l+9JvetCB8iwJH+kcDJ1q43r7A6uJvyQHekTihnt236DcPQduK/trUvk6S/Z4AGnTPEP6dI
JtHXOl7Zng3Mk8PqFHysw39ubBkub0cSCFaj05uRP82Vijf2fVbBNZWTlY2qm8Ou7FwFYTLVan3D
UE4eBL0hD4ek0xFGF3KxoeWkqD7jzMQKO9z4WhrxVCiv+X5DCnKNsDzYtJKbhToVA0prZw/CwMWm
QGZMogw6PeRppmzlFmSBPc5ynL8nx7YDODQy7wDozzPP/herzYQeZAhf1LlU1G1VFzGWCRH17pJG
EH74jsrXCO6+uvmj9KO+OFJs5K4vp3kmfZBMzfFqKY9RWyEceEC4LpkOUBCPKSt/N8ehvr15yiTr
9lgCt2TT7eVHltAhRhLgeVFRBx/82UyVWfYA621bR/5x/wC7dnedAINUPKqDUctgFrktXVsv2N4s
SpoeFiiJWIk/3SgRRJB6QjE5cTFmrgPoBCgS3JATwIdW0voMnO0IyqbWrz1kF6BIabzgkFGjC2Yy
r3ytxbSgCvOq2765C5xMua3Y10EkpRZRjvA69C3YeomkU1/GkYHntx61nlVKVyqrgnVI22WCxmss
86edU0zzygMVDoxICOCyG5WFO6Sv06fYberOrzvsAMOGZn845K02f2ED+KOeXn51bUCAjbAxOHlr
0Tpy0tlfz9kd70vfWq9Kn3nzOBaC4QHF8L13laUXqF0G0tE+i3OarD+Rf/H7hPrEKBffoRULaoyl
/NIlweajkrSpkPeciW3TyIVHli4wv8lrSTkv2kTM34udNFvJcNDlCzAKhU6P5G12rlAmwbXgryTU
wpGt1LYO56SiNSv2weehY6uAV7FGUFpDlY1zPsfAKQLbM86PEG4sPyi4owazQCy1P2ROjlpaYTF6
ymfAdgqSDbJJtBCEKsUYxnmrGtsv52MHmzmgvX94DY4mLnoQfE4Gk78vKADC+oNs5bBVJXPAaSXs
vWN/LJwXjyiUq8V2RJc4aqntZq8T1+rmgoXUnjY2sqohGPM/B/WIKJn4W0xhG5oU8UvvaU0Ksh3w
H0kw9G7/hna/QhU1NT4PQZ+suse+AC4EprUrUgL7GSFfsxMxsfYH1YpNBGK0mOCLJeIBHLq+9ArW
Ii8bkLKXzJnLyG5XpGSgXS5gfcrv5GfQHWxEaNN09J9f+Fa+WGQqQ0PuwKGZ+2iI/3M7xkz3cckz
IjTRw6C2BIc14Au6PLcV6iRq7yepf/5aDUG8K13YgxTsCVLc5jVxmL339UahlIlzr5badHdwSBue
mMWAjL0CRpZvb9ddcsC4JeLqZUkk8VmF/KF/gdGefAGFPJy1kcwtN/o2ucT1pkqFjFugS4fsEjNT
fwzegjoUJ7qFTeHMWcQlPQszAKopPZU49YJIwbOnoKvQ6kaAGMznR82K9PwPvN/1k/2TR5hlw9iq
jGgrFsuCR821iddNNJAMg7AK+zB8plPzMiGxPfObWwt6leZFx2vEJqDGN9HQMBhkYkIa25Fx0r2h
XFusRlf2FdGeaVrIgHxmIkIT8Ohon1D7NexeOV9jQjMkbbxCFNVfFQt/nYlUy27IVN3ohNyb0w/Q
2QCx1U6SUoX3tBSX6rmnPR5rVYh2n2jbj0Vmj0/EfOjmstVgcGRl6hPWYKeV9CD3F31a3Geh/ih1
vKhHK42Y2VKt6tSmhnaHlcXI0HWLU86VBEHuqIT9ZWArqfNh/B2r158yuFzifliVRbhyp2eI64qF
APCvvICu72QQUFH9KMfCIRcAvyjZnm93nXeZt+r5743yINCMuBmjNG4kNhk3GiFy5MvxV2kWaxEB
5XmBVy4pJk1sP7Yhv2e9uMJUP6nIvkflJODcJ27IX1qOK8FNztnE2KbvK2ZGGNtriMWSfooFiEm7
NhkZksBu2uRZ8K4DbowgT7svKW0tegR40ctiTA5oixBSnoEVySP+PHV/b1L8EyJpvrRABdRB6gHK
+PstBErFTT4s4RRC/dejYCv5wOXDtABFgkd1GFCJO2WPxDCRDQzE9vIq8KhNEY40/bUhRQ2W28kq
nyk5sec8dkfFYfy1hdEfDxeLONVxcAqcHHDwEUSFZTM4JIo+NxAahfL9kVmG1rkAOJY//3qj/+HK
TLiHCYguHRvqzF+7RACRlI05NcKspydBWpEccSqgRApBE5C22CekHT5+5orOWXw+h3g8JXDD6o6H
8kVAcX09INd6skrUJNHis4VY+FVPNSacg4a2azkiBXkYgHnMvs9VXPW4jUazMx7wVwl84nG10Y3z
tloHQG+gX0Xn6bNqJyX+OUh1+gsX1M2hqRvfJA0iKFkc/NDG8ufSCcwDcqJu5+DtkKYOVlSVRCCy
VWhtZ2CNuTLc6O/2SGFugBCHbwPdmpU0rhMGAyPhtdxRNVPM1nnGQxN+vUiWYDBLQucnCNuoQuog
mwvKVUgYy/NuSGg9ev0TnYKkzwPnlb8d8GPmLKnN2zlVNkA72WH68rUJEdTT88e7Y2DYc1aKqESV
5fm9EyR/H8y3TM+sqk2hxOtzOxYT+GSdh09arhdoM+K4H+QjlSAL1bJwedSODrD4F7B2FZVZRY7E
EjGRnS5a3Q05x3wS/2QoFfaoCilGtm0ae52J6xA25j4VEQg9U6IsSqqixYqFVyt6KRAxPPKg854T
+RAZeNzjtw+9CJk/R09ehoi6Hj5oJ1R+c0MFQ5uH1FbxZp0b6aqQCatv3PltSFAX7ZV8uCrUVm/J
/vEtTamnS5yQ7Tv0t/7XCPVLeKVp6NNecDph5bnzxzTUnpWen36qGlOrmi7W4of5Cmxw/uXBzvYV
YnCRQ8rlVkeVKn5+27DEMSuKrm3xBWJcGledsFjrn4uTAUlgudGQrMxC4qEYQYQFEfCYaonzLcPo
US4kCiC9lfbOdmESt4mWW7uM1j0xHne93p7MTuWuOKvw5F9YEym7TNBBp0vWPgg6JymKfJ6JOkOG
AG9feeYys348TqSrjSIhVGCY9KQuZuGC23kteQZudYy8RxoKhdCJfONN8IqGJ5vOZV4esdc1cqcv
cw/SLRSehe4aAJjuZAJVvaUYSI3JOHXuwb2lgUt35f9XphQEj/NKCTa8v6VPq6DOyTRyJBA0fYDV
kPiphmRUStsl/Jv3Ru08fo0jQq5zW1BY01atNOKAfyyQ1Iq9wFWEK+8Rg8x24jw3Pb0oIA990aJA
FHCJHhM8OWdwgWPFG/cd90NClRbpV1sLxM2toH1S8YWFR71A2EpzfM4YQ4k916dJa3Rb9/NU4iU0
iceEtwoUkKr4Xa+cojpayUIWHUoQWxiewohPDhYur6bxii+Gq/L+qihnebajgMG88e8G0IgxCPPp
g+PWGk3XqCbNekXzOWDfvTTWVjzhoKyZtShKmIl9VF7UnMAcuh01TSG1S1YdTlqmNf7YYQaoLbWM
6HripoDn69PozcChGjt1ehS8p7nemwqLu7OcTylEhHlOgUElPM/gOWJgAIuSr47eMbFFaotwnu8/
TEKBhmd5IX3L6HeQu68i9fzbBhaODKGPznGTQwQioeKGgIqPaMbQ0xtk8R73gcKWOmWopj/k6jhQ
DYPeWy9GIIyynE/UtDNazYkSSfomrrosZSAaRv0++KwOBnR5oMT8PT18VZjeC6la1es0eo/8Cn2K
iRrlEwhjwIaCwcYnBGhH72JxTViVrtjM0dVzR7kXDenrHIRIdxXScl+i9080x7+tnIg+395LSwLu
b2fNTGx8hg9V+zZ6hxQuJN4Zf4GTgbEToTH2ogf3hNEtCHlX+MUEXc53bkDkKTY42C3OaHKk0AaQ
afAKCkt44PRMEjxxe1RI1wiVVDO/t5zjtZ/P/w+HxPuM1+zUlzSDfcQ+ssbby27jzBRUK296JD22
J+STIGWY7iv3CFIMXjM0f+Ojt7Waz4pxT2BiKBcQLW8ha2QRQd25JuwuvmmDyqTXpwi08E/zvbyt
tyj0dbkGLCG24ppWFxUU/tcOMNuYxin2nxOI13Wy5bCFryI2KCOj/VPYTtA5kDhPhXfSwRs+5hA1
TOez40ZX7iMehn2Cbx7b29t8e7Zb4r7wWBE5VugEecrYKkLQCRBAIw6HMEWJLCcUxHru1g1PsgGz
P8dM4Lt5feEoMlIwmXyZUxMNFJAfunT1WIhAAHwqpXCSWjcnPjvXKCDVr/RQuKLhWRftwM7Vi15B
eqJMwlb2CIxtUiW+1aGvAU6nNgSjoT1wPFaVWHNt0eDeLNMYXc+MeP3U7CwSBZrWZrYBhrZ+27WG
NdRS6aqIbwdIVC50YIlg894maLTPyt6U6T+TBdYKku/HQmHig1Cvi4fy7lHQCb7SppXHO8HcSWg1
uzuK1cZQ1KR0+o4KYGDJYSc/OqMeYydM3+YbAdLgSxYbnH+P0uQaKWM5mgPQnaxllsDrqV70sZU6
6eZOaA1FjMYfKQpZA58sFZTMdh2hRcf6EOBXAfKNPzj6Wuu2+8y165F0dabkdYpk/yiozcUSqIp5
UkuukM3rT8ZnjugA9l+GFKT/pwS19IJ5lIOjhTi39xwz0B50Utpe63pzNYVXQWdQtshFhVGBc+TA
xcsWs6BZGvYw6PhvVeUoi8Lx5OT58XIQGHlMw1sJkzoXOLeH85lfrjsD2Dpr8isYkxv/oYRzlgHn
Q9Az95Z7pdogSNT4RjsePhEUhnai145iF49lBBdPzlHcFP11trcRib5nDuqtRxwiWevgjWpYweOY
rBpQFIU6Rzt0OQ+PRHHaAtt76HgPc9aH8TH9hGtu56z4uTQAqSM8jyDWTTzUZXPngprLYNSTR09Y
eQLca6fsudnYXgjkDwnJ6Y9cs7If14SbZwHfO+JtIGiaojaGejpN/HXtTAl4ltvf/wWH0ix7uVoG
zo5Q5118KV3EFi/C/yLC6D5Jr33c6tw5zjiffhTQXiwpWmnD5qzAsa1FkVhqgJcUafX5g/L+QNJz
1gGH1uDCgniemh/YuMilswTnpEWVSn3lvfl6WIhQ66VwNAU/rctud878W4ZhJwm3Weg0S87vzSzF
qIJbQpIBIR63CuEdcEv8KVFCiG+wye9noLKgplbIBk6lvdeKm6p5wrmALELL0c1ZTsmdbXtQk6ds
Ur+e6B1Eh5+ErHxC0Zb4uSGlLMwZm23oMxFRGhAjG15xWvC9MCIADVw70fuBMvmwNMk43P7uWAhN
s/BSn+mvuNN+vCiO5+zkBVczLrYp0rD7U+WKVdW08jiocsgZCqRIWz/h28AW1Z8opGTOjmMzl1XS
69hb9IFLoRpC7DGxNOyAiTR2LOiTTCfM9se3QUR7obc2Voj6VcGWi4MZHyDjHicXldMBoxrORbRf
0f3DoYBZKx/snziwQT/x6Uqzdqpxwfne02XK2Ud0OJKJITlMQ87TYtXqciJ7hJDyyC9gVvPLWqjs
0AzXIRjknx4wyPn6slEwusHCtdZzQk3XwVc5iJk8zTGy2I1JpHamlxbV0bNINxtK+zthueIWuuek
2K52CrOS65i6N5jYNSGgQ81A1vXzel5jnxlmVXXeo3omfV7zFXy7rSiwb1MGaNtbIl3Hm0kiBHIG
0pjcCPpdE1UW3Z/UBbJJz2xZeYp2YrLlXFUYB2HcOCD09KRM6Y7Kmh5mNVwXgE3dsVdDU8WCq5Ey
arkn1xKDfJCHwHIMjYG/pPuUW9Ckl8T09JLjEqN/I+1Gfa3SqLhqbVLrQwIcgtjJ8/OPy1AGPClx
X3kxMrDG77zipRxG3uXtvtdrvx5bB7fAKWWmcick333GGsaLXJ68pKHeEsBrTHtExg+7gZJT4Tix
qjHu+S6dYilMm/Q203T3Nt3JJcRxorWhIJU+HWccBFrbKggPtY+Cbz0dw0MQbXqJidGkbtNUcwPA
HPzcUWa0zd13KDabXL/QILPClwMyWxdL0jzJG7lWJbaNqdjm19ew8XKj0yQPviuoO9qOWHuCpv17
t6sDAt14P64d/xgyCnuYwMhQvgrvBWrsuC3ApQDFERsd4MYaARvOcY9wDNv7qMhFDwaP5pmVzni/
FORKNpynkKY0F0sePMPaRA01y6dYmj9En142f8t2zvXyOUiWurtp5oD0Hr0kxuTY7KP46kxVWXLA
NOb9vVNSWiQemRmb/vVjeSzQ0K/x/2s0UJ3icdO1kq3rLGXrUQtsALN3Rsd+3bB29yogAKxOjrj7
U2VTjFRsHbrLvXqOwBlQ9UtbYAUqyoYLa4L2pqtjBnXqR4dvYRS2d3iVvSpgDpygUXfZLXd3Zu3+
xtC2guCaNU3Mk/UschJDlpt2OUV7O0MZLApo5Hi0B/qVRsxeDSKt5zna0wvm/GwBx5AXZx4WmUun
Fp+W2K96FqzDPq1LAS6Tod4Zn3m17v7roSzByfEqbLW7h0NsInw0XnzKsk4vUc4ueH6hx6rAmaUA
4yHViFjUKjFHFdpfc23rdvs9/tliHqiYeSmX/KRmgqVXPg06bmTFYyA4ZA7ZbTMA44ri+XM1J4FH
XD4U2Br17YdmBHRJBSjLGwhfqqR/rTnOgeNJzEETNgJYsctvZZdI7g9OABCuHq21ZKcojWpAjpOd
rtjoUSBLPAuyOjJ7upapLTDfLALszReF/Vv1GPTljo0TJsxt6eemxlfNYLe5p6WPVywNxDJmmNjz
PKvZYEtlxB5GthuJv/t6P10azxAt27yBWujCjrEyc8OSfL572KzQRq8NbUmVeLJquc01VhDf33rz
pv09HE5FKbXm4UhxomZLe/kDLb5bn6eSq4T9unarPDPYXCk/6kH+0m7WKU4pyynLcWwAVEhicwui
ZoKZv7ctIkIKCLbZp7HcyIqgiaaLNuhlEogJUWh8sUjEGOEjn59TGRcC5L4QbkxRoApA3ltJEsUQ
R67qx4l3qKRHeEiZz8efJSBRIiYk2jrc6W4618OV9Ye/BvkX7yOILrcAyt9qrDjeYnSNQtIQkt14
zo9miXAjUbQzRJv2ZR1i/hYzo3+YIWdiroeyC+xy5aB/AbTtICJDdWB7A1M+/efVR5FOhQYiiNHb
RkFLKYwFwxylyDz2JxMlYPOkJGHKklJTbFKNznP07+aazmQNcUPAiUVjg6nWwJwp8IFhYAOIOE4K
5cCiSkSIU7PnxxTBclwb6UOlnQSK6B/oi7bitJX87y9YsQ2Gbu0FGhAX79l9O9Xcf/SlvwT4/KsA
qgGmbhCtfCow6/YfwPQBaLrWOlYgudMjh3kTcHKFe06SNhJ76FRUJtNYiSSNDT72QN60CrDwxGsD
9WXhK3IJajWgQcRWNV36AsaXId7Jv5HIxnDdcI1/h9hopobpw9tpIhlBvTn5kLjuQUy8+2RIDmJI
MtaUdAVltL3mjY+wIlVePI/q+Ocu7u5vU3fl6vsP8+PsoY62ajuj+knmw1rbLS5EiJpGPjf0IGc7
8xzvMnB8pSyzaG3REIACKgsh6UEI7NHx0zfv19ZTjHRG8GE6+JBXUqL+Ir0GEEKFnwzAl+kQzjcU
LCOSd6wdH5AncI5bEDB9W0rwTbjtkFfTUOmTwG8azb3nycZ7gUwwEIt0SSsjEzbb4S1hSUwoPA4K
Bkp1tA3eBA4Ki0GWX4x4prJusg9WAxm2RD2k7MhNRzO3NvHvTwUYGiD+HQjEEy1b7vK94CNKdSqp
3j05j0ApgOaljhymV14D+BJvelO2JEbhVhXLMJ0eFjEPsq6Etk11Mi4B0v1/3T45O3apJQW2mn0s
y9m7Ht9/P4XmXNYl+WRec6GFkOtkI5gi+XIiJM6rcN1VGqvHqAhX+LXIZF6USzXNT5XiQBvs02dF
Sw5rqmmcB6pcKkQK7WA5RW0yzzgYcHkYLUd04688Fm2WCyQzAOvSvy7g6ZAayVIA+0t+YgeSLSuk
N+S2/9HUPbHMKAwQRG8ObJJ2WVo71xpD/uP1ghTintmvk2j9r9ehAZrSK4Y3+JFo4B7yl8sxfodE
4M8rpAT6MAYOBxbHj/Jr6nqE2hHml0rC3MIv3hYs90mSAtnXaa5dDeHXAWh3t+KxIe8NLBfYl4eL
KBpXYPP/uk8Mtvw91OkoR1FqqKPFabSp1leZz73KZbFoIdffWfPpb1bMt3r115qnjdLnaXKNJCBg
kqM2C4h+IxqVOMyk9iKxpsQuvJbeAV/LRqZuAtIZOtg8ncp22C7W7rVU3z2ipnPxHAFu8IqbbtkJ
Iz2NXzrMra9KX+xBdB3CQxFeiLChRGsURhtMHxzAu1m4uYOU0FmooQL7Xw7D3hkmvbd6IK5UnW7B
v0+Pq0J6DsclwvmFcFV0YD1E5PcO/CifWmrM8GDAyXgQhq6sT0jto+O9tg63/oxEm+vkaITY7bII
nLsz76bziRAEbBL6OIeACD27e5mAKPAdce2i2jhTaX0c8vnDiTxX0H7xPQQgcrm/X0XlMN2Kkav1
azt+DZ5LUSaixD+GM/pRlX/3NVuUWc6XY4XNoLmO0f7jiyc2bqy7k56l2pdFbZ+8BqMChMCE1N1W
9mKiFb+5vQu5Wt3zBMNtjvZoAXnCae0ZqGtqKxKUPJ6LWGwYMBAu3crQU697cOJGHSLB6aUhjiel
PrSgHxTlXRnAY7HzsjbEBzeytUPFukOj79AK4Mid5naxO5Qoi1o22HbeRLkjzo520PPfLruycq9s
m5L8EvhVf5z1q/FpjByXoJX1NKWXQ6AYf5VWE+DuV8hy0HckoAb8qDhVHh9DS9SK9GJUpK3pHnaB
yBOnkwHLNzriojTRUZ1TnH9BQ0EPw6Xbazt/zLKnxcFPW93IVYSi0ULWyPi6RhOkK47pVWuhu1Kq
od1UuKrh4zvwlLCR2cCqrDIPKgLLg43Up/umTUQv2VsR4xSTT2/wWJ0maQ1kXPCjA1UO4wo8pRFS
vQwF7mKh3Qed+n92gqygpMTb6W2NEXxC2PuLKRYecBzpWibZP8nqfkpZMcMvxRTK3wOnF6j1ByJK
wwkaxfSxwL0Z9aDpvsgIfVTHkyIIYmGV55+r/gXOGgv+pZOVNJEgGKp+RMaiPwXuM1v43g3glLhA
v2Pa8Kzo7GHt8nulhzXsWJ8wFWcs2V9+kjE5b3azM0v9ZvwDk6ECDUCa9hY3wrcTkM9fVVyl9xJ8
N1xOJoXzYIdBEMJNiTrIOSbYsD6d79Pl9HL3KxVItFZzwYTWzNVFW9YAfD1fVoPxh1jgNo9oVFVh
9IozMWYtytmiw2Rwrsg2ge/qocYOrUG6W+nbDoru6/R9UExFlcR8ru1jMjhS8O7bylgzeGQ++W5w
NVsnlYAc+VxCSjIcenYIaIWf/CMR5Ql7m3oCl5IWGaPMb1TR+PfcpvJLTiHKguPdJDFT3uVx1y51
x55gfBEr4epT/1EZHcZs4qbB/blm8WQJmM8PbUOdfp56Jm4n89Jt7CUAzTuUENugC7H/zvY5jBdb
suNURTtIXJP+8vrghWihF5iQDiCLXeY+wpCY2PZx5d52XwGCZZHTYOOLiZNCy2aPrnJHbAl2eEnI
tdQkj0fkWn+MbfKenziFOF1XBPUIll5fSf63MFQt197v/Ja/2RmMgAj6Whxlp6Xd6kGalUQNasmV
bk1+h26Q9ZITvEDHog8QUY7lgTU9+hXhrWJpz3Q4IalnAy526N/ecDra+KfZa9aPO4wmRvS1xL8S
QaYsRB6nKbKu46cS7TdBZTvb1RRbL6+ZqJCErlbufH+8h1KFg4Rt+z/p+/5doknICosXXw1TySN2
S/C95L79ijbkxPVQuTj+JP2+WRp+J7QN/hYXM0H0mDZjwocWdIqgjGSlB2ogTbgOulzxhA/n0vkJ
qpB53oA8rMBgVaJs4ogF1CN69jWGaJnOzdKFFRVSLn5+vUQSy4ev2BkrLSlM9MRFDmspApnoFJkh
BsjR2ebRPgPh+lE7eE+QjzVKoQoUCZAoP4GHO2ILgxE8GEzz3inSgiATgi2EBA9WHy9T7z/0/ViF
aReB6D4Vm9Neke89EFZiE1bkQjJrdb8LEUQXN7xbRKkWt/N/rvFivmO9UK9Z1f1O2uQ7FEssumCA
62kwpBjFf9rgbt4JSQwOnvMmjqyegjpU55Mo7ZAImpCn8wtra8BaFb+iIsrhWHUnNww1ZNBsnq2Z
CJzZWVv8ONQCQmKqpeEEmsK1A7h+9pbwI23SsTsaKClI+esS25pkxIFt/gT9lcSB2s8OjOzp1ph4
kecy3s8WMX8In8vQYOq27OMnRy/YOzJBNArjLp350ND9uzwkwdYmZO2lthT04uTL041YLi1Wx2Tw
vwfQscT3XxBwjPe8AmfzNJeN5KQcXdOcBVzzeTxgZX3RVHORkONwilvlpKRt8pcI9Uy/TWDWtHhf
U7KS7DC81sUJGuWQofEBCEsp3mYHSS/Zm+DeEvWEZD1v19pwtZCKaiWzM8AQpE1xtE/8hXdN5iPe
ySzJVqUqqRpXKBjSOKTDwNLccNWKxv5avwcIIILFIpF8lGoWuiR03Db1xMLNXRWTKkJUTy/PuhnR
+Cv2f92SkFfxIy5umPNKoM2rC8qzA6tMXmkeB3BvvGsKI/mcRs8KmgLsWvh2ANuCuCLOxeRHYt71
ZwCvte99Xm3T+JpFaW7+01BkN70pGxiEV1GhOh246NVzWvc/oALUZp5l7XNzR623O8PU08yUb5dN
Emqpc05crZ3l7dUesD9XNVKY044wgOO4vfNlp+CICUbFFu4dSSEPrPDgFVCvHGIfF6crouc+KvzU
GygDDGs5hReym1zwT2wOs8x0Bytz3D/50H4uo5uKJuGSQ/JGKdSG8LS8JnDxRZVc+gzFZQ6kszzY
ePXlicEC7NqrGmInMVqiOjeHSwPFrMKMyw9/7LzHaX1WnjIJe+AW7yQdOUeIXEGI4LRa1XpSPSKy
SvekVkoy9JhAFHObJObXYIx+4zhhMiQZiC5MPXd1iCeg4nweH7ojGeqUtvpp0Hyn9IlYGVNdpbCX
zvKkVKC8C9Ny6tLpUgAzzwu0FoF/wrD6pYjK+7QT42oWsrJMHvApsKUegnIx7bk4v+e1a5qxHj9V
RtpSaU9m3RMGChcncQE3SS8nUkLLIGFY+9Rpb0iMmzW9b40EZdS5ZXAkVwDLv/RZvxskpOpVVfyM
fz/CXJeDjFfrdAQdooMjR40yYk0YSPZoTISmxtIiwzVCt9d7ZImZka8w6B8rhle7+JBDHmxkBmGx
oEeYIda5AbGbSO05DyERVT75g7kXUBBK46fwYjwnJMgs/mmKMc6Jyrco/9CQNKqHKvaO72txwDwk
8T3u4PAf9v7SusHvRgGKhQ6xqtRkg+up8dPT4EnPbeV68hPuXkm3TaD+k3zIkQ/JcSZ0PLsA0SkG
K+L9g5leY5eSyRc8cm4Zj7ga5hr9WIS5KfcWAVXuSeCUI8FCqUjfmJsRQxn5fN1NvbpaGr3fcw8D
YNxwbAZ11S+dFvVKCvuB4jksEQdtkGo4IO/pG5oEw6INKsbFJIdgecHMDBzmo6B7tHL5GbifkoOZ
hfZtaqG2bB3f4vqEL4DA8KLppfgD8JhKFwVfBGi2LdvshCYZ/GxqFUYhKIeH1lIxP5tYqchS79X5
erARgzdm0SXQYx5VCUiCIsHccFX41je+JRRx8csYc5XiqmpQanZH8c/s2LX7Lz6Poeg7Z3A0lk/3
wh4GZsePqElgk1him5ymF7SEg3de4SOWTS8Nij6WXiAq1+Z5tskWj5926Yz0pbMdZ9EQ9EzM3OOZ
FePIf1FwyFwggkDeJf2RwTwtROtxF0v07C+cNSOm8MyPkafyx3BHy8AKH7hJgWvs5Rbe21kRuFj8
k9n1oRC/mfoLzIOlUvX3WxlF7EIpGUkuqUaZc26ASeJmTGin9lBm4cb9BTxnJfVnJ9h1zLX7P11V
wxvfK7h4hG6iA5/l3RIrkUPFxd2TNNVU+5HjicfyUjGD1N9zsz7y9A8jB866rQbCRKliRgAuQDx4
ygRFuxCcbIQ5xi8tL/Fs1BplIOyDXS2Rur2h9mj6peHCaO5TH+sT3DB2shtKiX7PT5remcNSP0Lo
qW/XFw47p2549rlHBL165ki2p4qionCd7K8y+bfHrMZhqgoy6AAcsj7jtQVkXYfw/JUsMjtDGIXb
riFieNDeWB06/TU8/bITN/4M8Np/4vplHwsbPngKtkAx20CZ0eYx3cmo552K7cGGEnz2d1AanZQ2
oHVI74toqKEgvfMrUuGD4hJ72oGJjZ7khG84p2KvCQGNG7eFbaUCgxEyx1OIH1vBfOG19tkKXnrd
l/XUrhRE5G3u6cBBkiAz4LIWsw7/kG43EXbTH/QVoXXBTFE5PenksB3TpG1GbdSHj0AtsurLFi6s
ZNjQxyxqUwc1KTbJyCNYfSAycPXtzl4/h27yu3y/P9LtwWjzNdSMXVH6eu85ekOtysiC02mvFHE9
QrO+W7Lgy/sREp4BArTsLTdilbIPrByVfLnkm8jSew3cxqRwGL22EmWhnV0mtiqI3dcf4QWPFNXv
PBqPkaYlabY8IYxSMtOk0M1zS0cp7cGRu0Vuv5NmQfPJxRyX8I8hIwxIatVBkUk/FgEbDA76zK1T
dUfzv7lwU5yVff+8T9qQWClXRnxIBdkmv2HijYoId04vNFBHF/wU5urS27zyuLjLQzpNvjfWvOIk
+oM907iN3iojtXz+jpiJhg197nszH0QzBHdaAdfTJj/89s5u5gmtJJ1RF4xFBk6yHzuqos4lJPPt
6pYLQtPK+3137WVS3w9zIhPA5iNdlsmjkq/3tVxKYhc771AEVQXxHRyx85Tj4Z4d0JUOf6ZtRcHw
rBPP77v+Ejql2+JTMvAkVz2+uPGCrHqcSXYol5PmdTEqnW6F2oop9VxxXJpfqwchUlj9IH7wuNnf
+l7Qb7cNj7q5DUzwPvjqM4EDh/5q8uNITji9xTSJsCfqGDPCw79TTmVP5XuEAvwUl7iW4c7dUy33
TqkwmOIpgCJE8Q2CZpsgh6zMMvDjTJQ6blJJ6vhKzphVggqQ0jH9bLuWS+VqAltodJEF56VTWVvx
+Y6edoPA/YrlDVbPlOsUarCx4db3GGz/5kakzqh0qhYOnp+616daWTj2zOTpUnSw4wqiqKs+FUdj
drc9AqKx8kXeIck48PlYmTy9aTyLXHgptLLWn8UMEwCECsBj0jJBvECVEaTGCarZWSJ96ZLeTSWS
omroCBYMOf5YjtA6859qIhP6Je9z8EBXkVK+a3hQ/S4GyCWzFCMC9WhpXU3cPHb/1H8STGy08Nth
0TA6l94ty3frePWOuVcWHqINO59P6XMPMyH7xzm1L4GBpKmzAC+oeN9MDqeR9tNm7IoakAmqbL0j
HyMoUKdBfToVkZwWLuFNo5O408/3Cu7T+LuvnLlDHMHNx9JbQyUSFM8vZH4nsUzpG5Umq1CGMc6/
UMgbBsmlwZXs8bTEVvOxqYO3kN4vazzRSq6MYKmQ/75PrWw8dp4O9dLc9Ch4gG46h/WVpFIuB6wT
90YrPbGw36EO3sUHmtbUcWm1UWdvbh5l/sYo4MUXfTQhJTAg16MGukFDIXp89N3Zw8lz992HzIfX
2Gkqu9gWiJFxB+XqdMjFh3p4S95pIKJUOU9ju/bXXA1/yaslXc3cqJEDIcCa/bN7XvdNQCYq7i4C
cL5daQ5g3fqXkKT/B9gd7Vez4OYzDTW8UoiwvdDAN6ntdnfyYPK+VeTcpHieix4IKY/PYM6PBPIp
L0TQFX5iFx8IqBYSBcbFDjieOO7YDxECKi3Hrih9yFl/B4sGbMveP0GWveT01eQHB2Ef/pbGRoNG
nJ0kltuSmBCmP/8HXLfTATq85BqLuOsjHwHmiW79EkUqJQeva/pdCII9cBk1mCDnnoQ3cWdJ3i3x
Wu28kB5ZyWJOmHPOMRNQmElzVxKCDeGFZdX2VJ58t314+La1FdvmlQXowN+C8ZkJ1VsIuAMlT0CN
zlJjoPFoCtPslM5JRa72E2qGJHcO6c21CtaGm1l8oIJyC96YxigSGu/UFJJJYGu34RxG2eavOHby
o8EtugZqB46you3vcUcWc8toCmFXX7wuiROVc/9aylippE+09dgvhyTZBQ8AOnsg4uCSz/EvOraS
TKQEnwEc1GJt53fRJBDMYiH4xeCbUI7LUJqFCYCpUUDWWAj2MLaX7NYtsF6K4Uq0CVvnmBhY7kqG
lZMR4XZTGgZohIB2lm58NeepNRplfKH8kKjaGc+QaI43K96u2wVQjzoRi1wEjaUXwQqdwDlY4COr
ddMHKucui6Te5tTGCpKb931ZNWdtVz44LDBvaNUZAzybxHtxwNuiKGnxnC43zmJiXKqHYsQ/1ma6
07K+jlKpy8SOfHNlrQJTaS/UncNW6ta20D2rAgAl9fEusC2mtQsPdt+nO4EWvkEEmdAeLO3/KlxC
r/xSbQUwAeq55Q/8t3BC/75AzBNjt8ZfuZU2vnaFuhVFhzIOaaq3IwoMYHJ5xfmXwapuo+qb0Oxx
XJ2xmFtvQdLXfIpSEbAZLYW1lFl7ePqWoPKrZIQ773nB7xtfYVAap60Nx8H7HCPwRJg6lP4l8KZd
fM6bYYyULCyU0R1ed24qaddsb01es/baPdMnrSXsRo8tKtFy/RpkNzy06yIqXWXmvl91f7CQ7ngA
eYCK1emo1wgs6NpLT7DzxypXDfv+cdAT/DgKQKVmZ9kfzfkrghYg+dp6Dh22p4B8e89F2Rh+cGF1
zs2eEttO9BzpVme1s5sLt2npjV1GGlJ3qBfZnx+Sv5iB6nNyqM5v0aLyJTkU+a2PCc/WIYVPKOqe
8lw/fnfVQ65z5t3V435L5w/EruGANu65HHe2ODg7WiDky9bIPm6FHh0RdwXxC/jQbWO145wS7NI5
7/q0lR4VjpQsGYz6V1HsMtLzhsNbr/FgLCFCW7VTrTL+xFmnwFUswSDTaCT4HI/WW8fmBUL2HOE1
m69Y0qH2I69SipuUwiHBolXfNn2bpJT+4mi4tKDE21Bf8YBUeXxYEhbIqnknI8gQR2EFNKmY6M/T
FAm58Bza9qkaFQKMjpu01ZgdicudODac3F69ULaQurC/fbdkqt+hLhtDqsWAz2gD1G6ds9nOobfa
Cqa2vObDmAh9UQ9kRYImoOpbkBym2RXiDiGJUVhlC+q6n/lcSjd3ReQoIy/JO7i3v7k/iK+OaLwb
DoPJoacUmP6fKESxojZe5vPsdD1D8qPe5jDglOb5CbXaSouIjzNLqJMOiydGbxN1IdKyVYRzjQ+9
mKr0KHe2DWEKx9KhQGntjQysurjwv1BQSnOG0LAlElhHoCfSzPAUroFOWUCbRdWrS7fqURXjsbLk
syefqrP7/qn1Al6l03OH5eneoykSXvQgYt+Q9UO+6UDUrBoAMfdc0nyibZSKHybYDCxtzbcv/dLh
riuoq1E/vVVjyYfhh2K1zlS8/MBUg4lDil7LdWyS7b3bsYGvP15Gqu48UqBAWlwpyaMZZBHSRPxh
J32LtPExuwRQ8ZNIds/HLe6OKB13t1R9U05TGPq0pZvGMsenwG0U+ialxy+RlOI0HO5ny8czq8Y2
59NKSY6fgNIk+GtfmU3pYyqx+xrRmiIOuTmYfSQMSCNchrGMFmobPlULPfDqh4yLVCK/IwrC0Gk4
ToZ1PLEi+ch2nmH0ng5yaYMdrUsTcXx3Vci8aNZ0jqLO3dz83fjS5UIEHvKV2w2P5QHkL2ciN/7j
nbg3ISN7/7acB42M3is96u1ZaRlZ8bWJzZc6nfX3RGUxVCk7UluJSwWglSCY/eqBKN18AC7GVZGt
wnroq6psajrKGnrznjDcfeip0d4amBf5qRuixRKYTGCUwMnShCFrmR4Qqg67rG5TnN+pcOREj75+
FuXIk3IDSl4ahe6ZiXpZQrGUb3zStOSxpO1L4rROWqyx8ilptEhIoa04bVG30AQQMU6WRuxgTKfk
2kDEQeR5B/F4Us4rVIDlRoornZiDIrN+AATGg4xL9lZCG5FrtsUi3yBlpPa9LM+JpNrKu5fi1iVZ
CoTw1e54eZBWV07AhF1obOdL/GJkgHjiduT+6WePIgrpI6Kfw2y1eScNMhrHN1B7PEf8wN2n/hHr
2xX5r9jn1c9eMLWe9eAnoE6KcwXC41gP84Kx/O1O5PgEfVCWDYvlYYGkcsuUph1Ti9GZoALXwZM8
pUR+L9096kQgmPHnbCZGbS8x4vhha873wuDyeCVzlCC5y8DDYewCjbvj4ICCWkDXFRMfq7rrkaOS
fqWwiSBUo/FjnmRRorERbF1Gjny2TC482wuCY/htAzZXsiea186lhkZ6xGXMPtO6H9Sc/j5hs7X0
mBsNOs2FbU43EqdqURNwHe3CTYUBkr49+2dgA8DlVO+pd8SR+L6PQVdda7JfO7Htu5vdGI1zgSQK
7tmBEJ6rxFaDYvfavM42ZXkMXBijlaL8KOckuIRw67v9saTK++CTiiO0GZWlXhwfsTxCttqhWqa9
uUbjZGdVu+InDnm8OrRLO0DwKn55J94O88NQ18zNfJki2iCTPgCmahRV2WYoEsu2XHNjTLGi8ZTD
dciMpyjZiLqcXxfWy55CLiFcRg+TBIj9fJJfJxkFVpVl5YVQqkRYuAoetoylZJuw4U4qH0Nq3s4v
TdNcKRBWPVxBkNdr9aXf7f+xyOsvnZzvOQq05q88LAex9Wsazk6yzk8ryKLZc3ZVxyV5Zu8yEEQC
k1IIuu7F6OU03wJgRhMGL4vNw91FoEnnn6c9a0cwrLduO426lG/VmFq/DN1fgg0paI2Iws2+Wah5
EJ8zaTgp2d/jeSqX0TEZNf3B5/wTRm1/19s/edi19JGNBJEcMzuvmV8mrpJv7GtrF2tFPM7x0+tq
HwivYFR2T9WdyBWkFdoWvrv92K+RqnHXSH0H/3t9q8dvvPnGUscUWxcikIH64tkw/n3CPB/hBo7E
rc1MEAG9+QeCBAamD6GBPFIE81/hyFlEP5igDLkb/ljpyX36tk4ygaFefXxzKaQ6pCSRCVnnrneN
Yz661q1+Wp3StyDME5D7YWCb5rzL6uazWYMkk6HoFEZDNp6V75rfRQAsku9pPv/sX/BNAn1WRWyz
U42E1IZvoBnKYQMFMqGbHOaF0eT9sIE064ea7PB+kpkqt8QJc0LP1XOMhek4hbieL6DEbczjyL3F
5EsYMgjkF+RRgVz+tIH41lEGk3FelnBRsyJM3RXZ1+jjq7jaQzGtEjDlxqLL1ZU9tnpJf61oJLE8
P1hah4dLS5fT2xUyfDf9bBMlp6/toA7Ba1MdKlAcO+GD4OiyE1fXeMl2SfUjH8dkd5B/DZqVSlCK
aX7mQXH4svBUM/2z4FGz1PWG8jio+m7zBtwUMhlecnWHZ47DmY0huY5VplqxWBHLLGXGJb+0GWeI
D6QlPm1aA8ornrREgyxwsr4QrzGV0uuu8q5CelKViWpSd/1oUrCQpG3RgvXIhlK29YHVZqlewIA7
3fAQX+do9zU2pIHOnrjWozqgmKFx9AQoxLaBDrH/mvV7BeWg6mk2Z54Y/dGYqjRZoGjr6R6eIxoL
aJ5+ymnXiZSgat4jUerPMAt7AloKOUMjrIWLHwFkfN8hbm6Sbdu1HluMsi7K5ydhgTd+hbcjg4rC
OjzGejNOjxVtuMd2xaOX+ZoWbUmr5QhWij4vYkKKDiTkoROpimFYWD1QJU682dErpPUzs/vJ10bU
kFlHBi977PqituVnlQRCm72gIDrqWj2FzkHHRBBqZCi8gIytEN42nGY1jzUmvsXs+K/Hm45gyhSB
pdhadd0yH9Cc8PawdW1BF5bt4B9gTqykjy+CGtN1wHIfHJVQiagqvT0EdDaso2TauTGl9YKA535H
wOAGJrv6ESVJ1zDDItbl0AWvoLd9xjQuthCZjhMqEbb5NrZOsJkOyDwgLtII2gpjRbjoLhiu0v7f
6E0HAFj03q/tcZEMfhGRVkaq2LqDKYLCrdVb/hR3lWCqWjfQMzDv8+C8W6o72agWkWwJYLvTxyz8
6doO/Rv2o1OABb0T1wnDhdu9FHghUQV6YBUmmYOdV3FPdWZeBSLmVpFXMMzisSrqVRIs7kArxF+e
C8/XdLMH+Qwcj1EsubgOMnwkxgcjeXchyNds5fWpIvrvm2856V3db6ZR9qJp0LnA6GXun8dtALd0
iCIuRuzLgj9pCaBBd2MO4FwomDJwCokJEzD7d4u3pD90UytLVBoOPUF98fDjRzCymcgKYXevqiaR
IdHf+gT7O9a/SvFR6kp+HQIJhdSV27GJ8FIH4kQCVgRVePJ2t5ZbKqjgbp2JVAlPZggCjsWiv811
dgQm96BtxOlruH3ac5ksp6nptyOIT9e/ASiGJnunZBfp3A0/RNDSgpwMn6IrU6zCU1wEEiin6JBb
FMcec3mUd1OZujKTkhEAuEmiwbZ8iG5+PDiMs0Z9TAFpOZFsY606WDMI60LUWoOeflAD137rwEIY
qQA9ZT7xXt4SreM4V+6DbnY7RReP9lBeevS6GuJrdHYLNNltyhqHwKL50PHR2Y9qz7p4kIuu/tEx
GgfLEE4d4tJOH3CKtNhoydyhJLhatGzxiUUs8zD87XauOHu0pNB7eci4GFj3EXEtpkr4yGmxbqSS
whgiVY9DWGsGEdS57V3NnI0o2UfIxHcQl1+aQOq0s/94YuoQpl3YbcN0ZJtQqXRLJa0f6PViRnNI
NOMwA0PW1RJaNB3bfQuW3v5HyZTcUFOzYcu/cfPrqCsV0XS69rsxUbJcF+Lgg2tkSvMPim9fScxO
6ljMxQV1JVm3kk3kWHci5LPqcMeE0va2OTpFJ9ehrdWsns6F1F2m3nmOmTgR/kDBhSYLh+Ocy3RE
YYOcDQMZsXudt0J125mj6B5XItPvKPUycYth4BX00mChnNPW7UrFvVyrvHDbhHkAORG8s5rmH0S2
MvDK/7rLLxk3ViNVdl3XszCYiFzgGxpRzSSousrlRfegYBE9lh0Jl7DvuH426mKE9xa0oQtbu1gR
hPhxAUyKewigWcuwIO4gkiMukvimRtIy8jvvaZSHsHanldp6kfbzrOESrh1jXlsrOrE8Y4q2uB4t
CtxH9umVLbPGe8f9fuzjglqBubhVuH9Ag74lfqN3gnq2O39BFjeUriCjEtUSv+BwWIP+hx5NExbD
BewB9onO7TWQeiU5XpQ3osqolQS0yADUqL0AksDXq043kknleBTH9aI2AzA3Apviej9NIUszBbB0
0DhWX1miq8UaZH06iBuHTHR7Ry9qp22JE9yy0o7wAyQrgbsBwWxvhISuMygadIJsonlq0BZQnDmt
iSYFPqnD1p5CYDrFPUlqciprBTPXyOt/1+uaKn68MFkCXWBQDJpfRvfJqc3bn3ZrwgXidKlg8Hbo
/aF8C9qEh6hQfhJ+Hq1xySVSUANWoV4MLvH2gMiMBPFYRgFkE2ohUwu5xqa8SoBNa4zcsGOOg81J
ssGPmqf2/qU93YZOI7RIT/ACfoJ4Njdpaf+ImuSMVPDgKnSqPG7VxltRfvpH3pWw/30rXUPiKfI3
am9SAvxw0OhsFqBqd6/bbrC3bXD2ihXJ7J9hjpXCWUSyXW42HYm2oAIDrW7UUioS1a9cLIWDOv12
QWnW48ga3Zw8SxduSaVUVb+Xjy6yNqvSY2CKdW5o4PTHKwbeNJEUNam5lYD64Gln84+IKWHKuhvm
0WXBBfj8gwqlCSe39smF9VvHeu2Eq3Khw/vVIjCmRzbMnbZ9MoYqLF/IUf9YBIgSQUw5Ikg327tA
R1NQRC3oBj/mAw/uPufYlw/je/lhy/mIU0/CZagoQtsJ/pS59z/aQ5v+fIqm3ZFBzBwtIVKkH1iM
/2ENdq7Hif1ZOPQo3OboP55Xx+dEzQe6tCDnLAOtbtVad5e8LWBy5GQg1RMVqrwmGNRivP+Ib0g7
p/l9wYN2ZWUIaiS6X+1lEMjKeKKuT/LBW0ZiMEnsQfrTA4Bpbga+rMQ7TYKUsM0bBz5rBNjpoeqg
6c8vasAl9sdzHgR2pGotUocrKH+LahNhvVJqnEytKOmk5GHPD9+O28KOiQhbSv0rK9oHWwQk+pCV
swI697W5s3F1RA43GeAqTEX9z3LZPgTzNDEu1uNoDgNCTBzTPnezkBScDxyQaGhciQbZHhTJR15G
ugRyPTGG5af5OMGbXyvcHleSdSH9Tmc7taIlC2c009wwmmv3DYTJf2CWRpmPnfCWW+mTNSWU/t4U
jb7lne6eiBH9JOULF2KnVQYsfHDraHjRofEDge6MzukfVNwml4u8u3GxdswYIKvom2o4haNW1dIn
hLju+6n38jyjC6x7T31INXjr0DkrBLli8Dip97FE4/N8e6FLoe6v9d/Jg9Ml96bzmzLuy11Y+aQ9
WyqLkZ3+nJLOzNekwav+Qji5wsvDmfoR5GAxy2mtYA90lUc0bzvaj0IIBU3sXzwrdKgbFQhnUps8
B97pEGOXixWzeBir5k6MDSDiN3fqpuLUMFq4tcsXVc30sZogNt/r3yU4tMgBxPmVDgygxrL9Afz8
DX/Aqp20k2FrKAQTeqsI0tQmNBE96yif5KY+oFXbXOKADEvM+O5Q+grctFUCRZS36ei9MwayGs2e
4LDdRdNQDCkjZE9vh443T0NSb7c00wbNcMSz4o/VekyeiDXsGqOFB6Aq2mlXRYKDB1pRp7QcQCyB
iZ/4eenT7O/NL3q3N/zP2Ggm84t7tPGjxEv2qAOhPyC/w1RrPoy8LZXKekNk9B4PTI/DtMetINW4
g9znsDx32bCFODU53Ogd6zpVTOtPEK3fWbiiP+bEU0NNajFqF7q6nW9/1JJu8Pxyt4o5aS/sq02E
Os5drFEdb99ZHQP8TUB66NdszSNiGA6du9+OWNBNRBgqCt0G1BbpSKbWY46YaDFY9ZxgD6KqHzuo
HT7SD7RA0SUdr/fYenH68Bz/E/SMzd/I3N9c/R6Req9NuUFBx1uXiI0DLNjjCepW/SM2gm+QpgTd
0qp22lD/HX3XjnMjtVaYIBhsrio/W1Tk093fRq0rfHhy4GDHYrKQ16qIeoMlW7ZncSOotoxyksqB
E0qesc1YOaMPAGGL5Ehj38Ize6ds5WE9VLaMwduXii0ws6L6tGaG0TbLa8ddvWIizD63sAKw8GD6
bBKqEh4P+6ZjZ88aWcpF31tSZhReODTUy84kSVNuTojZwD2RK8O7ybSAeiSmjOvpuBbGHf6Vz2U2
m8Lzo0wsk0wQ8pAeCcFAf0Vzpy0LkUA6Xz2U1rFBF2cKQyTR+vEfAbnoG7krmqGUfazX+jSVi/+o
do2qyY7ud99CJqqBZNidRqB5sjJ+tCmUl3i23A5/3ngjnMCM4tA1mYWCnGEcxhIunfPjfisSVK+I
Ld4/iIzgdu6xAiTY4MuItYkoVr7rhwPGYj0bQ8jZYL3Fj0VcqC0Dbg4e57qE1UOhc9BuwIwweMiU
DWSEpSSS16oL4YRmSnB1AIW7T1tk3oV5ZRIeOKKPbwCpYuC1iO9Huq2oc1YA/h/qecySxgWf0F3J
pjG3CGa7h/vCeU882y7iE4iPIhsBvhJW4c91ftF7D+it0pp1/Z4Y+k5ZhR2BNVTwXqKL6w3w4gZm
OXMYr6ZTVubOK1KSH0IzuOXIBtqopEbDeGGMcpblX7LK/Ui2ykpFx2W77eAWZSkeG5Hhwlh/r7uM
4GkgP6pSbAzdEc6vamxAAozFMuny4JHYC3E++fo1HeEEv4+Hiyk+JzTIGbdSg0pJb1/88CUcbyiD
jDZMBDkizKCbcqA+oeFFPTzmwWnyZmHttwfq3Vkd3mwUOheyuLccCheuxsXvSccMUJYVk4lpYNaV
fU054x2vdy4lUeI6o6O10Tgp//n32WFfDGs7MZmyQ+cdileC/Ya/nGbHMjsG2eho0anG2LVL0VSG
2c0Oztj+YuxjDzztXTvaYAI8zE/Hk5c/rMxJxrTfeMmC/0PNDr8EUf9pDS3ndzaOTkJtL3xMLN9u
NQuohPn6xQ50Lm5Bs4r6jfcE+q59B0TehxHvwS7/3onyd1AkA0m4YSkFLhcubg8ZOeSr1ARGd9SY
4Lr7PV8dNIG5zyiIGqpCCZU7/Yd8lxus0yKeEYmfYlAbp05fmBizzSJQkndBtr/Ybd2tJOB4EGzk
jtaSL5LpsjTa3XvVntbQ3MzgzxFV/F/wcp2YJtmH9cbdwBdf3jV6T90drV7MhsLV8cfrhJsstaIo
60bgiQlqT2JkBBRi3SnG/Gmepc1HAl/hXRKvCyrp7571cxT3Fv/kuIKi+GvY+trVnl7gD+i9sesO
NlpPL+sM5ma5H/9NAO3w1nCb4Ryh9EV0mk5xmp8xcLHDaHx35lGial29s1o9gMvWsJxkePJvDDRJ
Leet0gUfIw9d30msRky0n7ytCwI+MNsefB/C3Vy//DPfPX/wd3XxpKcK6HJtY7B0B/JgOn7YDS5e
HAPgrht+GWSIDLJroYnB/knpXxf9ol9prbNkWvXRBMqjQRjERRIN+xdLJbWEkqOGTCQQ0ykMOlRr
JyHFWmCqQIf5rOw7Ht5UhLIUWy+Rbzo6EyblI6U4T5J4KbMW7Y90mVAEXk//IVJVp0A09uNC3DCd
UtQo7GDu7H42UluhD48Mp378AQzC+Qa/Pa52a0uiu4w1vNbKcpl6KfN5IcV+UnRUfTcX5Movko27
xlhQOrHt0ekhsUy+bDO/wvvgxKvshNV7YBqwSNRmZpldYIipG28SgvPRMWzRHcgO28vI9bN4cPn7
fXsvXnXXu6mqxLmi/zDAZgt6nv5fzNO7p9H+EpMTaB/2wEiuVuv36oqbm78zTMC4+4VseFHE8yxq
oSUs6PncXGWZ/66bfeHrkJgq33fHR9D2flhmsPQOwcRA7son/y19TpImLHzDwSrLNmC4YFlTwZdK
Jq2RlC4WAJgo8ph8pcuz1i5ScqHk8RE5onzQ+hGqueDhnijccYYf4iSfybVi3uEmVJHVxpYdY6Wq
x8d0hVQWSzGtBICvQp91bj1E9W/0Hn33dwmy4qtLmtMDOhA4TdWF+YsHaeSgMUFeBS7vPXEDBsV4
Lzv+qqCKEtJ8M1Sx12OFIL4rYIZYa6OP5ZnZXI7njxVYVX3odTV36wSc+54lBnb68d1W0bInVlqt
xd4Vm4n8H859iBY5V+MzXTL+SEqOK6ymHk8Ln3T5/sdmK3H7yIr5PU27fWclH8YkMbMZc08Kc4RO
QQlLm2Y4mepnO6MaZ+Jrz9PARR04dngTj22U88MT1UYmMA+dhgc3d/eQ5rJppWS3ITNA8/q3ewkp
9THXQVgHHPTb+VMVLb+A3amr7suT1sUDF132Y3M7QwvR0acr1+xUsLA0qusRfB9cNpl0BJKqPfvF
4XtfXgowElRApF5w48xC+kOopCKByG0fxZGZOd8P0WCMgR46bEuzt3W+TOHs+vPm8dlktWQD3XQf
tBYm6sz2ZQHKMw8pPtrk/EYJNuYuAsmuG+vukYxM4tZl0oQkeOxRH86QzramarYWyy5FOY9wNlVy
bVexrHvdk71WVaXkNU+OitBDTrvN57ZFbLN3AxKuW+eQvtMYGyW0q4RWtBST9hcbyo2Vpq/+vZfX
Rrfzw5vu1/nzfi9z9yCdlOL06QABMmqXkQpZyhA7B+od8MWMaoOtX33mwBQQ/amSbg5Xibn7wIuN
9gf9cQPj63FhT5Csgdtm5h8pbeJZupUsx9bBkzNsyE1JasyvGSJ+DG6wSdvW3btCIm6DCwUXQLWb
koHjftm3DrRi0B46w32iEqjYeArneqksnWPJ7DC+3M2hph9ROluzKoFeXjIeD8u9RpT1ZMtTav8t
eXCdag9QTPVPyDPzJEmeX2A3UET5zUxoL1I3sX4GZKuR2bulxgJMVWu2dVGf7Cg2x0smwHMV7p77
JabcveDH5H4P9gUD7p7sm0Rp8PDJ63TeS6EAoCLsbafYOIrCaMYY/Vuzd7EiwJJ6qRThdWCrBgrz
pQpj0VLBzqxbKiKUbD2BBWKSADl7qQRY47Ika/OXrau/fQDyv3zCFZlrB7c+qecUK9STkGPfRNzx
lPiDfh/mUzjxFEZRiWeFR/G2ISR/B2lio2uIe1KUoEHTNx1p9aXWW+Anud2Oi3HzbPj3uzbRC6yF
VNdELpSOcbx+rv7nmS+JaxDhu+PVMhENx0T+1iFpOG3oJpEUFfBM/ypmUE1BtjWp75+eDkBEqMLk
FLKFQ+zD+0p+zFXsc5MZdR68Et0sMG7d/Rw3u8mR0RQnD9dfS3xJzg+lJIYuoxRh7n9sSajlsdsz
3TebEXPciVuAD1wzSJ+lRJ8p0ZIJuMHq16nAEMf0hOJI3CnSiRwrjzZuSfF5dAPK1KMn4Ev4a+om
CSYF9aOk4SPe3oWSpou4o72/t+G9hDvaIgefEYq69V+kr/Fjhf01dJqlMpqzQrpm2XryWaHwSoI4
V8q1VK/BpLkv1fLSqpFuTriOD22hae3G847pSsimVqZ94WsOif3Ce3/Aq2S2zoEIcdyP0NzIR8GG
H/U6TtIfhduWzR3KGW9qMJeyrNw9KbaGplN69JVy+zvUemTIH8eiP33j63Rvd68a6zSm7oCXdFDq
428A8Bc+bv5IWzFNv0UfkaMgF62fcBMOymrHEBxpKuD+PSvqL45rl/es4VSI+zjKYOil1/v0owL4
jUm4zSzd6vR71soA+vj2cecrX5gYd4G39RtpCD5fQn9xP51ccfrg6JW86Vi2y3hP5A5VfHP8KZLJ
+eWO9GW7bcuJmx/3i3Dx0s7pABjXSiqmYvf77pbsNzvuphDY37M3G9RVwc1CsQbU7vq1H668OTR9
BHVwBt38mDhhfz+BKhtb2PZL7eXryJpbk996pH053LMFTgoXEbUUE/pPsRJAjhp1G3QRVeNfOtVh
fU1EKxtkMgb2w4diCMtbhW3dcpf8BhKmXatjkXcgNdFgpC06i/L7K9f5BaaK/U8Fwoz9b+4p/3jW
2R3no4i0+V17NRS+VaNMFV7juWIjv8VrWN6RUXDwcORxEi12pxkvLZeA1lJNt4xSNqvy8ddybZ4r
h6Uv5tMOeL4hrmIEXTOcI7aF8w5rcXq0HMaA9KGHxfS3HQ1JwcuGdWCVqtl+rF14zlenuTPb2BIE
80JINgkZMciBa6VbVgX9NYNIcE4vf33BRnXSl+oJrRNgF9qDlvDQqv6YFtEWDkzC43xkxjl0tVR9
NHVZeB5i2y20IiR5fOSgef57Xan8XonecCnqQ6mDUqtZDh/ZlHtdq+mPFtzXhDXgkcj5ZuSGRNLN
1vM88hadl2bTICL8LffQrjT4KDsJbApXnb6+4mNjsm5qA9WhcTJOebk1BYY1uOdx+Utli/Geaip9
3MretMi/o3NWzmya7i0qsVNyUzy4ipKmrq0uNDPZSSK8WYFaCPwLmkH+/YRzcvLVAXjz4i53dPi3
zlyeZcBu7GVQwBU4ndVxU3qTcyY7q3M5UQb6+u3xUDAqZLsZZK+n33OcVYDjLe4vEZaUh1bXVtEh
p+ipSFaiY/7KRluFw3oUXFgmV+wshrrpPSc6aix/Dt5+POFTLG8AuJrj4pB6W9RXFUUCy0O8c718
et9yfj7x7ze+hFzfqfVQ0clO/gKOWP2r2qY4cTCUGvMI71Yw0WJ1FoUw4pVFACpG8KTDXa3Bo64Y
+xi2qPAV2edQHJIcAUVUTjXvC1WZ6q3Abv+ewJkX2hW14T6EEddihYLJRBgt79dbmsafAVVV2YGt
2lQtXAlvJ3OBMs0iIdzeuVjzimNQZxE0GPnanaYO7COfuPu0RMkbOEYN7SOGX4JcMWH1nbUGv5r5
0+bHDvLnfuqzHRebG14WkQZq7181nCZ1fHqJqdZ60xcmuFUt8BrLy+CMh5xbj0QZdPD3AXif27Vj
oZlahWkDNUfBXX5OdeURvfMBsG9hzoGM/VXI1rDSZV2nhttvZ+PyA8edx8eLuQIBWXy1mPX0ugmd
H0Y/vbsXlx2NHKoTdhNMOeRtJDs+VZnQUT1dVJczClYwrsk3tEsPZ5u/tPXdBBhLIa3H1mzzaBkJ
7qZJNnEj+qZJ+QHgU/IoKsPuMkn/Jo3ZN4x3UGyQxFzYfD0mGX6YzV86jEQmhJhoyCbn3HU+VySy
GNSP48CAt6tJ9ExWo7AyAEbpbBd0/iFxPgYwueoXPPSgUUiOQ1W7LM9Vd4j9jsYJFWhe90usci3G
7t1VcbPbTHmPimx/w5NQnehMxG5cuarHT8m5GPmlY3rsGR73did2K7y5wKV2TeBXJHInVtUV5mmb
3eOw+xErxowCYItKbfLA9I1fTmF2FzU/abSCm8ySC6HrGMEFjELUN0vS8GiZ1ZDPpJB22uwZ93WA
5AdB8G4VG9dRw9vr0nwJlC9CX3NO6lHnLYF5nplFPWB3ip+HwY2YOuJ5GrEKhteKeQoRNA07INjF
2bgO8GujT1k3s6+MCpBVGcAtntu2DIXjyCS/b6bOlAI4LDEMxKwyKQbhehW4kPyQwAV5ZRcVrViW
pVoFISlOyHCkwTNeEx9hIWNk7+1oRRvp6B+PEavORHTd85nsht3P7xtiyAJ9Nuwp0V+Jjur5GPsl
NOouDbHOtCFqt1CQ4Rj//+9y8wujufvDRbDAV4Q4KTFSX7Z5bvDNpJg100ZCTCBziFwsJrP5iOet
z+Bl8YmMAf8f7+1B+N/Dpnhl/VXkGRGlXOGwWuOkmvpdsBS+RlnPA4Ir24zMDjQMD7WT9QAhzDms
dibY5lW4zhD0j1Ejdb3usWpMXDI3Hd6cdeaNHP1g7bXtanIJxsh8EKTnL/5sgIaxCzSBVSz9Li9T
Uq2Ywds6YkjUBck0Ewz686FFUKhRsAN4biTfr/kuiQ7CgjBk2UzE7lRg7XnKsgnckJw/+jmKatMZ
xINbQvMoFucfsj1u6VMOoylE8hTX2XnZWDJqi6yyDIrNnsRYA8ZKj3Y8nTXN6lU/aLBiAqK7EAK4
gU5Cr567Tj4W9fg3BwoIzwgM3u2J5PLAaKbzsCW3EFPBoPN9+HHfWw9KTATHLd1A3tCo9fmGPAfG
lqxQrB8hcA5j3waxcRZ0z+9RsrRVpXUtZZs/64m3XUOGZ6NnGcKepyab82oM7Wq0MxWl/qpbE86c
QP/XWmMw2/xJbV7sNg9PbBxSpg0NSnAPMHhGtjvZBpldGXXJ7NVyuM4xqHw6Ii9qPO+EDVdsS0pp
FTmFJWbyfBmGJQBZGAw2h+u/wpVGnIivqKwzrzcyclo2pqGY8CZGP3KKp752swyDcaJQDBszqXBx
AhpyHhsZwi+kGuoY9OroFGzJWeEFVISqLLE2fPlgzJsEGdPhDxi5pNAbt8d/m9d7neAv8kI+SKYs
ZemUhQwDgO+Jin+uh3BDIWoynTFHLCYaAL7tXjqqDiEnmjEbCEoQuRKUtr2amOS8wmWHQmXJP/vb
hDRq1zgquAdWsZ54GWA7Y3YzrpAAt3Tsgof08wQec1IHYfFy7pslf0/o+86JLVo+lE1iduyomeyS
rgbyynrDdl26IQj1qvGrwT0YIyD2uN398fR59vaFRoUGk0D7fLb9O6QR0la2ZEho7WiC3w4y02uh
AEeVQ6Bum5+b8lQ+KUGrzeC1hMteCrjPogrq8ioOM/lZQLYywBV8qzK1nITy+zRRY8tznfD2H24i
DUDPhwuD4TXoP+N8Z47QTyVTpkJ3xIz9ikx+2EXHll00jljeqO9o5pTi9S+cG2refVFLlNnH8XS2
//YThnCxJ6cgqp8E+srgXWQ/c4dn5e7PfY6YxAEZSHMTprUJDu3670Z0wBUCF6pBC35ufYkLO5J6
ZldKk1p10VODwThmw/3AwWw7vaiFsAgypL34ZBfrS+R7zUK6TL4SqL9r64v+GSiQHJW2ePt8Ysy8
XzLVtWt9EMy/9MQpavjyv4ld7XEifOC9H5zEYcvqTnsPuch5wHCDtA6+wYE/4dcR7oV4eKM6iR14
hvFLGpOAo5na7HmzJ2zfIYTt5XG5o2+lY7VqHmLZSMM8TX1Bj5IimKoccpUIfrCRMyYs7qM66Qjm
ALESdzSkGIY+Wk3o/5u3mx5LHfgC7rXBOZnn5NstBL2qrsG7GKijKOU5onuBiORiDNm4itQqrurR
au0nyaHQgnfQIfG9N4ngh8AKH4tR0EB7fnGfjJjkreHLGP5LXK6eZuwlkeHjdGImgjfNpOjW5RMw
dwzZjYo7rKlqN5kP719kVICYZ98OB5iuYuVnH8A/TJw6yETCQ96JlDqSGybPGLj8GXceIsQ5IgpP
YSKi9O3u1Xi8iTJzmVZ0LtOgfO69eNeVJElxKC8OmsXUNbZiXTsKFE3AbKPRYUjyOAyiyNoi42Iu
/MSGKgXF/fu9lDlDkVcNvYHI24I0zJUA4VRVKm6Hdbf4gq4tJ4puoJFERwLCbHRDdk/nixIKjzD+
avowtW2V7HfVamdX54qIkOD2t9Pg6JpvNG0/rv6JjQZLYy37dXznxhg4KW1Asmj0GU8USb2+CmD/
5XbEw7Em3p56lbDilQCjbsCbnnLeLqNBG8dwDQAFKzv1D3CrRcyEmZTYlCpCxDjzxxpNOMig09W3
48YfvKwNGhYtgAIHnQ0H8eLxKYK7ouUBwMKXNnaYWL7XPyJJb4wXpIceV0h1UTlAuWmD/37WZ3a2
czmUZW7h7DXQDL8rueEaURl0xv5CG3TsBVlXIrvdsV+wnijzeTL/ukP3WGvlLCdppZTNPsgBFoSN
TKvl5QGaclDEvHid8zDKo2cSq5PjZ+BdxJudFEENSO+1oFigxV6nsP43cBkM6fuIkQS10+CuvMmd
AWijMcKkMRiPX80JhKgulgwr7KLYL8p+22Sdc8k/gYMDG7t/O1uk8sOGUn8Hxf2RTFSPctQoEtGa
QMEXkfaTX2bsDjsQpbQ0nF3+d9H+eKfJFr/0z/A+Y63g2OwOpYaU3WU07gq/B4tpth0NhneHy8dr
p9QGlQ/zkpbf2ju2XtwV+Csge3IG1INoKpBkMbJFFdwr72DzGKbzCzd+Z0ZLJulEJ4wddCBGhjlE
2DEBv0BsXx47Yw4kdDSKw6gG0dw9KaH5qfVypBiZ161MvB2LODFSCXC6dULCCYtOqAflS7ROXAGi
kzRTEXmMAK943l0W0+nL0hm7IxvGLqYUsYxHI/SK1C7j7a0yt/IliI59zt3rvfbJXBlINaJD+yx6
X8aBiGdroho/0RZnjFjbwKJ1UPwoP2/bEudgu2HE+DSV2Lw0YD7uRoAB+I8jhirNM7BkARs1mrhg
JuK3fT2r3VbiPXIIrYngBo/VWGoun9bnQ/fsYeTUKHnaFknRujyFWvrZZnhT7zf/j76A0RXbZVYJ
ZchTRNd0H8BMHMyNHOF7GmOCXq+DHQOdWRssFOla6LHxE3EauEBhjqVcHnVHrfoQ/FGxUPjP36wS
AJAo63JcAJ0x4Ok83d4ZQ6mo3r9VV5IZtxcILI+hwkIwKXj0VCnkiyzTth9hhvPNS4LBAZtmMlB4
8lilxAAAnW+s+c1wQ9NcWNOmUEUSyh6Oq4tXS3SpLz4g0oCWEgSKu3V5aNXD57pLgUEU9w/YIlCk
qxX2Gh2JO/rk4xaBJxKI1CNH4l5dpbuvxYUCzySnm47qebfHOUmsspQDnYwzmtDQV2yAjMiERj5L
Nh/Fh0VvgWPnSFC9augryS5Usze8uMFeHoh11uQ3b0SREobBUXXrL3Lx08hfm/fEjJbnAlLWSd+c
EffD4Fc8pg/t99DvS8PSN6SRS1u8XztUWl3ab0Xtm2uBt5r0WHiF7ijINEoPyl/scg2VxhxaJM6T
1AsUa9yGi3a9qPVVBYD5N7VSi6qSDtLey3vpgmIJ5Sh87bxdqa+pRMetPZoEniBKtA3zyAxbyKVs
PCtaaVMfWGZG5TLhlZq8g14f0DhpEQCC/FVXiz9XXVE+bHWCGEfDCCK2xF2rhmHGMH4+RuQISsfR
QtRylbj2bkBrs47PvkYL+I5dr7SXBppB/HEZSPk+pScw7DOPbZniQN6qMqpzqF5FSmAKlGQQRdPb
7P3kRaTK0bciEnkywmEEdd7X4YUWR0y614bnUr74viI4bQlgnv9Oh4pbzHMou5TmPO2+zSKxJzaL
oEzz60c1+Lh11Ko1rEw0++fN35rbg1TWoLlQwOGQIPAIJ3LMLz2Td4ogF53G/40K8N7NXW5TfNgf
FPyKCt9HlvKG3FHhi8qURC8ilCRup3UncpBHSkuyykaercPV1uRdZzwaR8RK6NkTIEANW9UO5jpy
JDdMFXwRR6Fij0KL2ZNtYuZn6Px8+kBG8HzUW8x7Oy4W4N9rAOMIYxUCDZ3MXawVEOHK5XN64zI0
6IMuThPleTfP9XTsKKebmY3jPRVM/DckSc+3m7J4BiKuXnLc3lQHEROcrB6fl+TR8KezBqfDN1ba
+FJhf4FQfTm1axXEktfIYZgMSnU9X3jTCxzEBuml0nuJg93CJNNmEEafOz+cGCM+uPzDWSrI0ziG
dhRdP2sgDeQ3oUobV5wk7pGwgaSERIvD6WcDcuOeUHPEmbOHikyYgamXNnG+iTCd3YUnPylrgC2u
tPkROUssRl0TD5iBeL5zd7+P+3VEyWR5v/+t4MU8nsBbNTojH80Vci/94Md+KZk5r7S9XwXAXUYu
SLZtYSGrJPRkpp2QVqkuNzZGZKeJA7lEstM9q14TNzJB608mTIHfFkThy+VIfmYvAlFKCi4jFyV5
tstFWkvxLfK8Iq8tTEDEqLLsMiJ7QAWoYVd+bYmoBd+nEieLxnEZRHavVTKIs/m+J0m6sydYkJHa
Tvhc56uzitkfk86XnDwnykclkiGHdXYzh+F3ae2n4iDc67MGG7KTnUfVBfG9nPabzHPkMwdsVZSG
/FtrbcsYLqZJf9q3oaWZVAjn8G2MW0xXwHByIP48QXexX1kao+LSbuhJigQAgSiiwH76IduLFxqZ
kmzts+SeFPJhRN+qkz+sJybChGRGXtPrKSWpF0WUG7tecZUJgcPWq8fcUEH2deP0Wvxa8miXzCpn
bdRC5fHYlfh+Cl4iJaWj3sjrSe8W/WhKMVJu0MX42dbo/rC05LjSM4lknKXElEeCPMgAAb40HZSO
JVoQwhb2BEr/tKQqU617obKGkhDaBOUAWsNX2vGnUoIsYLAyz7yfPiWEPwWXT5EgZ+8mGSAmQ5Oy
iEkKVMcF+qGggQdSYfSUDRCb8pAnVQv45J5rdpNr2j2bATe+QuT/Q3xF7wpbKJ7lrAQ9cMroHwBj
9XnWM1M1ds+ki/BnNgu52yFKfHhkkie7ZSJftl2Ww/3wb1+F3x4SBDDGju18LrXUJSQ5kPMikiMc
/sKm9UpKX8cvTpKTp5DmfJd/RC1U5rCvkgZprEPP5XMUDPiCopzRAWeNa2lfWmNekqcs+OChBLOx
Ogxo6cTh8vTFxcLDBMt1JRy2hjuYEYihiY2kHJB8kClAvoXjinyQdvogDz6OpheNmVqLzzMkUYuf
Wklv+pLVSPUo//36nA2AdBByAeyMA1p574JGTnwJTVoZZq34+EocNTHp3obrp3VrdxwiHekzg6vo
R+tIJc0nbHKx7xkvvyYbey0NusA5bQe4ZPoRmmzg35g+3EHHIDfMHH60nZHssB76n+picPp87Hx+
4N8+nAmPIqBWd2yvLBgxn/cfn0LSgmelSLMFQoxcPiGqP+0s9qwaXHMrKo+U2O4eq/sN1uhKdFZt
14tzLkjoBBzVFg3Fc0hmatF0HyYDMw/14/tgYC3nhgrwSPctkSwpVYP45oRABKqhiNzo5nUk/VlJ
FVPaV9D5d9Mp2GF/ueft3YDwmVd2jigcEuPYErDmEsGLIJX5678fGiRCO5s1jerrMPylC9Tw1O0m
RAxr0OBmJmvzMHTzEnAUq9FL+dY2OwkDgyYJtmwH9adEyUafHMnlnbnHTySt1FocInd5iE4LrHUF
DCyJkDEiry4HX0JMHQDmTEe4aaFnKZNjS3LItv9eWC58KRPsWA5t92Nz9eD6dNc38SRbYcFZExlP
qZUaZzVeH0TMJi8kVMT36m7Krq3d0SLBtbpPuYmcOW0nP02t4b6Sj2t6wQ1J/ZUX2aDH5QfWMr45
neIzot8+a7p9JPoe6trCYMVVw0pWzuEKPm0B8syi6ImFtT35EFCkiqXcKp3d+Av9vtlVXPC5EnlH
2S0Vo3E6UwgG4/bubTY6lt0bLWEoWl+KZ6QNu4Xmmvvm2OurrDwxWsU4UcVyC3kOe3RRFQoe44Xh
GAkVJQLuuxNOAfrdffgp79zOT0WNMSMXj5+ymv+vLnpGjVChjfS1fEi8Ur8G1+qt8BBEgkoNCApk
TC2H3Arbrn3abOlR4F+HhAWMynvUA3IjTPJqdvlW1/zVy2cMcWjhBRbiOmM3Jw8qCpIazHj2nSXJ
3gYqL/1coCyXcgOqgNt2uL5EXpZxhqQteaAz8dn5OQqzo3INeKKCFxbBwd5gFtc76gckmgs4SnQR
pUmNo7NQghdr7VRvVk6gyPyHOdUgRkobp1ap2Cvrsa/EjBysrfhhq8BfW3tU4UHU5WO28dIC70n5
UHeYe7Y1VEqpphdsoikfvON/9ofzTWhbYe8LbnDe4lQ34kFYXeCPU0g07VPk87Q08Z98aEnbGV5f
8lXKdxjfdz84n54frjiodVrMubLmUwnK4L2g0Xwf9YpvLPUK8ipD0VXsGpFdvTT1pwZh9aRhsWtJ
iZw1BYnDNRDDVptpJW4b6ZmT7ix46slnp6om4nlfSyVTZcr5+VfWCyCqkIOYe0Gi7qrS0SmEw62t
JF42OAkDgkMQXxQX8lXy9cYvnrFFAUnbs8n9CXSpXKYiImUfb8yESlebePGt7NGMg3ZsnVZE+Hsm
3Ak/yg9c2QaxKB5JF0kIMCtHZ0Nni/W099qPqPs3lk04/0fgTRIv/lChsAlOgaVWK/+V7ESHwvRX
ltEGYLVpCdhiH70coaPsqrsKqGi6eQMZpvAPb2r55Juff4uarVk1/xbtyOh54zEzUDkhtMqM95EA
NFPV277fzHivHdtgNHILbtUNkBRUcuf4EtmLzJsQb+gWLed6rJW0dk/Ra5as+3dkKEPKPjfVkmde
/UZZ3VUW7xfKzn3OCAFh4Am+s9XxzYRObPqDQzL1LsCQaVSkmXpgL9mu/eCi5TO9yQpOgl4PAJY3
nOxPQbBULObJIOrK+KxpQ4rPfPOSsZihTVbeWhcu4Y0tZCREKyrTS5VSAIkWHPfQnRhR0WCIMhDY
rffoH6BKjwH02KGzH6Nxeijeo9n+xyVRkGaDmZa0dcqBljblnhKgtXJqog+Ui8Kz7rtpG6mfXNLe
2W3EpGd2uOUpDu050cSQq81A0IfbhvrHLJy+miR93+9M/Ie+ZFSjKJBGD2a9G9765ouKKe5FA1lR
nNV02vh1fxHMaQYruLJz/NNTAWbzLF1dhLrzyScjN7/sLIohG1HMs8pmGQ+XkHPI7/jJZxfzP0Fp
3Ys3PMWObJ4+OBegOWswdign/1wA2r3Q7244jHR8t5s14HvhGeJqH7+3/SWthz9NPheYs0umeuFF
a2Pn+yf84a8mmvSyPTCMA4ne1Ca9kKvv82x04jjFZYSF9RID5QxP0EyaU0tKVEldWdz6YHX+N73h
3xxXkK+TMCuCR19hj62ZXTJYMxpQpeLivDJSj5OmvOqSdkoI1e6NFF2n6G723aiDDH62clePCRvQ
kOxo9DUud0uGTcM1KggA5007YdXDTr4A02uYNnMLspu5yyVxhudHR27QYeXu2+jhc+pTZ1E8cU8+
ktVa0gbC7Buf0vnxgaKSUcSPV+3VWwyezpqDnZaypZthbGMamrC6i68ZMzRbvkL87MtoNaEriuZe
j9IU8eD2p8aGLb/vW51Qh7RMU8g3zsKc2dKH4R5DZrBmUkmadiU2PEXZXb3X4IZ7Q6PIR/B0uqwK
XPcq0YtoX8b1jG7pMYAnw1YKtgWA9iobXRrh8kM4Iv3lOXJa/faZrifLi64vft6dI7HfQ7Fp9ePl
jg5MsWOWAdf56ktZMUKMj7g65akEUUs5I67t5+GGjzrFJxQGZ4gfIT8cP/Myfg3uaJBzsst7vWXK
viajem++58b7wg8hmpA6i4ou2E8WrGjWaFBuDEbf5E9Fqsgavs+hJrb7qzmy/CYV2Y89AhFVoBvA
cNevpUq5NtYlTpS7M76EKeWsUSWSqPlKNrhQ5pEavW/ivX22LvejS81QKIVhT03kzVkW9/pzM8We
wKNMqUfrxd/MyJduPt9KxNJev3zaP0cY/CIBDpOC/Jo5/9/K87V97kTEXLJ0RHTRTJJovZDzqmxv
HoIH7OKYHKl86pmDbFYpIr5LilvMARMXxDlHuefXkBhxipAUtIJyq4LRbF8TGTq1irWJpQWJNWq6
A+gFRP2VF3JPkMcO3INidy9G/D4MaihCLnt08CI+Ms6Wb+de61KqUSkrFo8jVYgw2KNucYLPvlU5
RUO1vb0OYRxL8wfBGirD9eLo3S3CKLFiqaIfuJQ3nzD+t2FvJYzpA0DH05KAonTUon+t//6lStNa
MKsJbHXALja7jtmenhAptFqUFiYsID5zha+I4RBhVqPoYMAJkl/8KKPc9QxDpjBd/1qv1uYgHCKM
WzUZ+LFilTKsD+Y36N4qAtQYcUUQnf4Dh8MJcLQ1j+Arp3+3vLEBolmaqqd1CZVnkAT3Jxbs9exV
dHMJ1tcem5e5pl6ITZ9mUJG77ag8Jn+il3ay07KkUcR+0HGfJ1pg6lI3RPwgXyYaIIBAEYMRPHFx
zn6+nHM4ItLnMs9IrtVUiKP9M/QLYntEe1tKxpLmXlS4fGmArAkALYSVfmguZjbWmLHvd1TTr6Id
mm64C+6Ir1rbEzt1ICi8+ys5GoAwBvOXr8dfpikg9B+fhGfeEosrbS8qid2+E6giBqGkF5yzRMls
cr23KpXDTs7SWmgHHWExLzyOZf3BiFbNkfAQtN5jjOyp1hK3FakVQsDCZlaTuSDAejWVGnFiHHBI
c2g9YXDY2h/6WosyknhvllDKOHR7wqHmAz+0zP/3CCN7tIY18uOUTo8QpMLKnTxGItjnNa05c4DR
H2b8aNo47w15MuG/SpmDgZqw1foxdk/x6W+MrbjCRf27ERVvG1ehHU9v01EUrW45WxEdxwFMTrUu
M75TcD+dhWVaI3g/bA3+sP8lVGRx3CBXcn3tGdrJnvlDLEugZO5SZqZig+1Jsc6B0jy7pbFiEdPE
UeUrRSYDKzAKrj7ahLvpwCySgFn7wI9XPmr5SArSAM7bUcXaU3+2PfZMfGoIWSJYkd9ZDDfopOid
sbi7ZYceyapq7fBxMvSLY2MxFXfDaVgXEgN7EO1WD7aCn1LCXQLXPE4naou+2OOObq8A2T5JBKGf
AZiEFCuIwBK2V9pjkAsenBzSqK4ZB8ticfsPzBn0MM5i0wSjnle47ADej+1Uedqt6KVYG8gI9IoR
d2n4SRdCy8ZeTM0LloTzF8yN6XVHR2FD2SkCUbUwVaVmQu9XeTpk95S3/BW+HCjfGPlUx2U6MpRR
IE2bIR51Xolwx/2BE7CSKVcq188F0KH+tq9Uwf+UnWbk/ra4L9kKdkORU030grR0/gWbUtDhEE9g
kMQrzBpqPoWNNs2ob3MBkwaViPa9doZ2ELjCerARkQDMl6GRBbxWmOIU/Jm5ufUQ6tUNVgQpqw6Y
TEyM+4cAo1+XoCKrowalUf0S86C8DkO6iDzyJngBedGGTlk+apJfbn4T4oC4CBmfXHX8Pg/Cs69R
PNMq90B5XivVO2I6GRx5KTX1rk2x/3CMjJ+UYOJ2ynrpDA2CNGDvlwujnALD92QWZxdTKmf6fqj9
M7VAi9LjIA5uwu5pFe6GVhuZZsU+36COO00LFhRfS9IN2mTDy2TNXQwAEOL973/yiIjkIF87vAbD
nfqjJ+00x/hzKMTYs4uoMkJwQUN941uzmwLLnKqu9+uCy9o6GmNy3jA4CO2LDyo4Vz874r8hoYVq
kiuk77sIbRQCi9vLG1apF13tFHP68xqYmhbTnWpbPEgSditm5HryfBqa5R/afTNCV/GVol8r1bdM
RsQykDxUQrzdXHAymYxHIXCMirPFPTb9i76/bFtF9oUfAYOwdgsC1gIeJfHZ7qK8VufsStWTv1nh
/K8pnvi2it+yq/uyK8+VNBUCGxcc8gHTAPC9d4w6qGHu8zZuzGQgG8axs90zWI7OnDwjCs07nq6y
FeMgzhSV4Vx6UFrP+T5H1osaYrBJuQS8LzXvJzTFS8E2WTytixmWEy1Dln/I0D2HgfYsd7cb2y8C
3IkBFx6s2JGt+ivN4LGFn/PLOk6Z5rC9/oPlin0GWJ8AS4xOvJxAJZFTica5MsFkp7CQ1xs/PkOY
MQnDx+dIooqKxZvmfXZFUXqW89EJcD2MfY2Hr1wXdDDlTcwyrKRnWf77LGzabebFeFPboLxo48/f
+YsimS7hNexNdg2Sj3Gr7fNRvLZhcInJDNI7iLuFKNIXurAE8sFfKJkGzewUP3RqozB+m9Zxren9
tb8SKnQQxZmDEubuHSqBeyRnDi9uEQ9P+j3xJtFekbQaeObiWq2XjHCwznGawhBWBJCzxBRazCvh
6JdOBJJOzZp7Z5c119Ta/rw+XGNt9S/6J5+EzOLh8t0k2SRTtZddcCVdgk8GL/YagaO5v87gzZth
zT19e1uFX1agD87sMMrG2xx8OgzV1oRcJFBXv5H+dzUuVMC5FgZdHzLTW3QTV7FV+CQwnXz8Wp6a
vOmkFAhhzQw45+N2U7wcv47VlVGFXQXlPA/LLTsIiR7JL3JjZ3BlpsvvH8ZyCORPl+8eDVAQC2jA
1GpUxueKzrwXzH9IZ/dowW3nFvVt32IkmAtoG0gIwZdlWs5b7zAgXskkXonxGLGQtiNfoDupGcpl
pypsvwYyht7fQDmzLanRtVxV3fC3AhIcAC6fPkDJtPE3svN/wlWfHN/JH4EfpgObrL97VbcdTD1O
cbiwLugHYuwY0MF9dFMNcV6s9+d5B7lb9/m5TemJ1Fw59ivJpqamKjwt2ulxTo55PEbZaoRs5A+V
R6pxmctEpO5EiDYkRZUmD2glZEd5SJnLEH70d1L3yLVdWl5lyRsAtn07DACHFXHNbL2g1Tgg9JZ+
nQ7s6UGaPxiBLWh62AsfVdWFAirVQu8LFXmerrtkH5jzr6W3sddNtHNlDN14n+5CMNbXwyp90xjx
drKQn2GsAT0Vc0IW0DMJz17muVBNBgZmOS8Odns5hrFGg8WjmEVrYGL2TVNgk6dOB2iVmjiS862o
2vMJLWyZpFSIU2pkyeHV1Tx22EfnFJ2DpsT2sKun5OTwU4BA/ozwqHxBzZkYGgWChug266eSNRGL
p+DRzCpDuZiF36YJYav9Nmt81Xn5Au48Y+Y7fKd8KD1r2ICT5j9179Ce75xbBW/Z/QIGIEDaX1tD
LgTpc0waPthZRS7fw9i8oroaajIqjVLMlJ/He9MJ7OFBW8/NQFbgJ0Y2J8PabW4UTIzD2vwN/cV6
qZFnTqCaZ+yy9AsTk61fQtOeUq/WG0o6CFvWnUvtMCq8nfUGKooDoevPr2kQTQECaZor5ypeu+Hc
0UlpsK46DwMzUX/pOWjfsbZJorLMokRgkbdpby9OKC89ps7vDnglxPHXQb00iWu0ty/sf6BW4CDh
eL/v4q6GIclmYtwhIFizp94X1afJoaxpq8h4nW7+pVj3sKQwcL/02c4vc8DvILWwUkOHjrK0j8Cx
anYrHOGsgMCGv50WEkgRA/DrllZRWXt+6TC5dYkvvDWJCzzp1S1WXHLrRfMOLOgcjBh6l6Z0vmYf
TPv/faZDPxJy8+x7vpsojltd3G0jVtEogMzYMUe7Z5/IlWDl4gyWG0nMxfTgMbFAKiZ2FQY1oANV
XMPxyhmXnMirGgQzluXCURJV8LfJCSDALcrIuuVTl2HVrIRBOlvq37OgAZfsw+0fsWFYX0n17Qbv
7e+71XuwaNvqxOIlg2U+5tA3uN1eTuvnNEjmqXbNqj/o/J5hUFkzb/HnYge3jGAjLxn8lfTJxEsG
qFQaarFEorPyuTl8cOZjJ7a2sEMahdGpzmpjKklOie4bburJ89rRdOZTQVWwC4fewS3Iiy51FjUz
njOUReaXbhhf7tEwSQAC8VtUhme6VlTvwdlbH4QMNU1qlxtmZaQqEmfHjQ4p3occ9J6ijfsaqZXF
AyNX5BrdVgaqhYC4eXdCVetnFHmuuPPh+fbe31HyyLjq6xJv2fd4W+I8ljXL/94yXDXJ1AxDsQXs
R/e/UuujG38Yvw6qo9n/C9kPP7DjAABUvZbQxIBtMN4aPCY1Ltt5Qem7/PS4ANL8/gG07DOwhjSv
fKNC+l0bK3Xl9Ucq3V55ImENfr+QHv3X3xeOVMODgq7W2W3Q0/WY0REDj5hHqYqsiDnx39rctwPv
2LbQIQxC8uDw4/ICoe0ra9o4yFhw7giDYOcBERe32/KoImFISp9tsAZeE2zrOwdEPYEZ6foofIOd
IsCyRWrbE2oHgWLJtPDYez64XZIqTSrjEVxyNCRvwsRIPCdFiVYhQmSr1X0CjV7u1UZvMU4Zb/tt
lzsOshn12KYEDxPGJB3/pX7UDwX9OfQa9aj6IbeqQ83rVFeHyhc3v4yYnO3PcBwbpGXk3FF2Qaj2
vppSnOiVGpluOvl3pIC4NjyEO2vvITlfwovna1sDSvwBlEjGYa5nIGyNSjt6cxTMELUTewKTUn9y
Cof3ZVg3xhwALzJEZo50lInF0uNm6eGd+QZhuW8F2TsUFTpyg4oFsAv/1nM0WPCMUJVE0cYcetOg
Gxrbn1kKCdZtBOCxT2RBA2Aj3HaidyyMvnWy1Ur38nifyV02Coo5i5dIlhwF7WjYoMbS8SlsiXWK
fxWGszjbj+endGlkYo/rPWLc1SH36O2WPz9rPHXk+chThMaMdSZrgeJDk/c6WF/AZR55eW0bRbjr
5i+COXiro9vYiNPEyn5cGH/cXYo7ZJ/hko2q5ApNAFrgTbEqCG9gzKKkUw6DZqwzzMEsmX/JB5UK
1y9xAAWI47ESfieRuTdAajJaLblGQVQZLEx1kfH8et2XjErXrH+qL+iqy9zsJvqBTD6EBCT9P/RV
TvLZgzxrEHFOTg4l83RRyM2n3AxQ1MQ3OcYn9yNpkibgYMJAUCelrNsOdDloOs+17NdVjeGQ7Nkp
PxEFexaDQrlMcZt+XRyU5DpkrLQJmBeFMQ59qcM3TX36KkbnJawnq5CFAYB8y08Vxf/ub4D7Dm7s
kE8OitUh1XEMiLYZ3QR9fQBmtgKDRDphVy7n5scJx9ycTPfRsU08gRt29jNYoBRVGf1AeRncitwA
XB0k6NuWVK+tsPUTCTKigJUjd0wUM7nvz0GPuCif81csUgsLrxnN0g47Ny7dqK1yRiOjAUqu0vgh
zbuGA1bw6Zz31wHdxD7lcyJaPB/oNgv8AMsOhQcIAV4rF9Fbgeu3GlqJrXS57NUdIK4tZyI7trFE
oxzMe+G4SS30ySOfGJlkzk9ICIlh9v0UNxdhjgAgQ0JQLBRxg63E736i3B/q7D30SvPZW7WukVGV
k60zT3WR1kjL3ec8uCCenGV7b3Owyqvsw8pVfhEYEv15UjFXA0Y+fY4iZqK4b8os+7BVSYAmJDim
Nn8YbdJkVVJN4erPlCvqJBI8iwmP5bClCxsRjQMKVJMCZ6iNe9mFk6Z2fL8yai70cIZbiuUJwh+7
DjrtxfwJncwPpYYKywpshf8qQx3SggVF4zlTWCWkmYj2Z6HlJL8LRVyslk/RFfBMJmeNcBaiDbsT
8rz2AMuJSiW0q91VXP0VtfwFwQI3YxIkftxLB/GLKzExAidMNo7Y4TFXRiF1KlYN+3DV5ZYUJ56T
z7oI7pVCXkcbDpUARuTvAcBzlAY4Y5xUKI2uo6dad3miQnIXYQFs0RqLpAsQYCdCV1okBzc30oZG
adfHXSz6rCrAsj6Mm3CDzBKRaBg7mNeIu0eEDFcwLBxjCDFqRdWrKqayJP7Di7TISIzBDqJKJlBz
qnu9ZBL6x+hLD+jPbG+m+bMnvbzwsiZahYjWg81h6/RITH+lzQu3EeBUBkd5hVYNhYOKtfQggvZK
l0FKEGD0++eNP9Mj1vSR5pnUnS2h5E4nl5tBcFqVtcniNJEsCaxNoLjFHl3NDzhQsF7mnAssoJX6
7/ubf36xNsLKQb3df4qfbHhnO87y+3KHo7kebCpdtoQtXokY8I47xc6Xindq+j/DJOET+4Z+e/Cy
G13oiflt+nW2JpgVGUse2uaimWCFOVeOJyL8qw5Ua5d4K+YFeDPtA3RZWAkJUrSEPTUfLZXOwQhe
fsKUh8m2vkxrHyjOdcsKUIpSfCLdCbasXvYoxk20lzFblMPEUPrCbgA7vrZOPihCAylPKwa8XIY1
Efp2QcsB2gUFYyf9Bgs6DKat0bv47js1oYuK5mZjFnpCC7Ci4QYKw6rqgKnYbgSxtxAkyTLOSnKd
M1PzqXCzPNbZOxIAeC+ZyrzVyCcCbJ9Rwl4I98BBA9bSMAYefofbybnDqoO0AR+M9L7GV3We5dqV
FsPGoquH2af+0u1CEESWhqmuRkwLnH7ppgQa8v10nrj8YhV7NBZQR+xwYPdGjhCauxyiQdYWvpUL
4OYCrfH5eWoNrgC4zOsBAhaaVKcXsZPzrDtCYX/U5XXwl4ag0iiO4opgyb2f2m+LvYsr1I4XmprU
+mG5nyJTJPrJrcnTNcvahvZWivsmVRTgSwWHjkK48rjuQmhoVLJEVGGTWiUqCpUKZcFmWOEa6R1j
jNRXrS6YGZWham4PZCCD+Un6h5lqidB3rGfzrbI0BDnTdntULbyuaZemrrsSLH/MyFITnga2qcAM
3ZJgn62DQUVGTmLabVwFsOweLQtldhGGRrXHN/PoGiiNkVgayCm94OarzAb9mTgrAqCrWx7nyLBy
rICP4xus7IRXQMx0KlYdCmL5LDBdKH5rR20xMJHXAsgEniuI4Bq2xVcGgoOFbvLDzi0wEh2jRGTv
94chBRufL/OMWadUWw/KYPOf0n++iukNO2eObL5bkLBx2Z2JzTjfx1vmG/NSHGyUybdpc74p1zx2
SLicUpN+xevHw+dS8wJLTT3jsMV16yRtDn1G1ZUvVpAzEfywtR7B9dZVZkkNfSTk/65qA1UGCq/9
GojDharXVKVLPo6ezykXeO11PS/XpBpJ3UdpJjENK77iann64z+2uH6ps1h4oBjnJeFhuuLX2yOx
Qgl7+WPOdFrhyLffCnibaKBGNMkmA3/KQiciPCmYHcNyvZWqrkzMNEczWrUQjOOy4Hwepl94oo4V
/TzMVaaH/I0irEskF1uR4o7bjLYxoqQQmOXhtqM7yaIPOtrIgO5K8gmKWHvnf/T/wjbDEwStvfHx
ajpkNy1KR9b48+dy8JaWwwtQp3sAuOEf8QxIcKdrd0LdiymYzNVkZTmIlNt8K/ymO2u6HFoza6a/
kVPtNtSH6ZhymuJyyK0+D882uFlFbsQIDur2dRECRXoU3zXt+pts8uQLdJabNqF4DZN9/tyZZtUN
6M7uEiWgQMRxT2ll06HbcwHSI4A97v3HawMSrXLqQ25tTRGL6J4YBiQFy+GQdtd2qcVn3km8JWfU
zDDPmupKerU/g7xh6VmyAEAt06Johwhd+gaQCHyIrhQaj55HL1xrVDWci0R0h/ejbBi918vNQDRP
Y2IeIb6WvVLqjTek4jTRo9V4yaDPtEYSI7YZ6/NvrleiZCDLpgRBsFFrATlhF9Npvk7K/Do/geDZ
/cxXylGUJSbQikAzl/FImmT99jMLslQOuRM+tPYcYtV0N3m7y4zTxpYFyTfA/ymxbKdDf77t3N8y
5iQIFfsd2H7EsxEBnkVBq4h+VSwAC0F76CE+aIGf8HF49kMLLTYrckGnVDMhC7BvdtAjYZgCbWmo
8/eYSFqc+UwtP6kOh+Sw3YNkAmkTKSl5BVunlxFfex5K7CIwQ/YoHY32fviw0MdnAtExGcosuQNa
eeRwtpjDF40znjbmMOH76pqUmpn2y81xhXCn4crtyumglVDojzWTlexAi5BW4ZlUphzQjaKczEB3
znwmMt9ZtnwEW8qWSQJDiwQEV/mE31aN3lA87+R4Zs/iqUpLGXr4ITY69Ohg47Q2iYFJudKam4cm
Z1IHkz+/t8OzJn18eL9NzLTucK9leo4a331chSLAM5fV5mjaKx5wa1PoqjV2uVimZqL7GhSHE+UM
w0ZB/ilfivADlRa55sPRuwg5WN1h8L8LWeml2s04PdOvzdRq2w562A71vJPMVbuWXWzk4OseTpy8
0hdwGLmXAXIH6F06ZSYL1eC3ZHmI1HlcrDZfV8uVAHvXxfyAEJPwlOPWqToD3bIfKxmZJkblV/i0
hiI3Vp5RXCdUAKITbSO+27HlbWfyP2no6yh8clVxqzqwuhbmtZSWesu53M+VH4Kudjw/rIKqH1B0
5GnLjUxctN8kzErefBe2wJHpEm6vQA/e5neX8f0bOPcMIn3tT1/VlwX1KqOG+AV6G/sMe2BCHbJj
Dd15f9+GEsgO55U55s5fg30zPne9YfPtb9Ezmyy3P09m42ty2yK44ISXx3v6B/pcej39YqLqPPVE
Y13MkvYS01hdN+gcclalRoS3KkF/xXfFqi6c/sk8pfQsH1tPornt4PomiSbHaAlPQ7oPVUaNAroV
0WE1URgZd05zJIqudRfPQQElFDTEgKDMPVwmPODytfD7a0oPMh2vm1J1ophS8EZV5dml4MdcjSX6
lzC5us2n/4qBnZ5bOOfFzaSOdObw/litA+NE0fnB0YEq4vPpg6opiSQccHL4ENBzSIg67yGLoBqj
HIN+0Js0Q0mTf/AVJ0/aJCuB1JUyf1IG49eqOElj7fGU3C4/LW26Zdqy0M3BHjcxvqqgR3R43fES
EYapIRdaPJSkcdXeQZQ/xy70EiJRr/2Qd1V1PYkmuxkYnlvp5I5Uk9ZbPzWW/6hP2FRzPJtG9vLQ
Yrew+e6JOJrN1Al/cah74JJWpFkIL8lb6QjcxoGesJRmk1A8N2yT5GEeB70iMGwEFBi1Dg1xUnKq
JC1ONVhKrydQ1R6VkVGCog6R+EK1U+zU9691JpH3nKBCXd7krMxML2JjhFfEzNSbYM8Sc7vAmqKJ
Nz88/gocKYueSUP3wExkiFoV7PNcLQVbkRXJtLY0oYNxh8ARakL+wKqi7DtmbUkiZX9KfYQEq3ow
IwEZuEzH3HknPkNgpcgQuFpKf3YlvARM8YYUskg3j7vmrajMjMXFgHOHHV15bVLS2tbzYBkbf38r
rKlDDITnem1TI51xFzpro1/cFK7HWW2dqf6+JS47BrgHLYsT69rc577zWPhB/i+/ZdhvGLXIJsd7
ahgztTLiCV0/OOEK0SBiopttLfevoSAUrA6/RJT63qkDygBghqc0KQ58xyVhdL2Rz0VxoYGukMd4
n9Xv7XwI+MhCWgEuL2p2RG43gI03YwB0dOy01A1CAO97aDDRvjA+JCFCQ3YgKZlx9AJOD+uvj/px
un9jRfru4X34MkYJ+SmfUQNNfWIJPqoR4BHoIISayR85ZpVwKzowZccqWCpzRnvAzi7dybksucK9
v/trOthjstKCvz8iZ87yEWLq8Ir0hheKE/9tIyrBUtvfV+wi45f6LtaG+WZraXh4tk0qhB8B/TSL
7TJR+2DnXo4YnJmv9QuGAN/nINKsFEqV/GmXrsmBsfYZAo2WBD5euvc7PoGwLRvMVn/UID9sLXNs
zYsMqiQbMJ8fwTlFM/ygtMMs9BoS/kChJPDwyQFcs7nzmqt0GgQk9GylT0WlRRTcsLccZ3kTNn3Z
Hu+5zHsaO3aqoucXzuc6JL245ALwPth5AJ8lZLrWG9NQzoHYJ4gVWEU3DIzLfVy/1awmlCvmQCh3
8FgFo6Q2nMNA4EJYOO3XIuOS0QgETLlQsJcoWdcXi+TF2vLQl96Mhouzn9x3My4+bUvUtGxExCJ0
9uUzIrXZFzifiHbuJcDG8XQTf/jnpiNk8rjI0IsZz9eW6fkB9HW97GoB6A+6+YmnCmLRSFt+HEbR
ueZXn5oAvITzYNfcTGDYys+EcXazo25TpvPo/3Tgaj5vIuXcuqve9kFiDScDkDkF5l2UKhwH/LNK
1QW09tVVl2dx0wgFORct9ZXA7hYmsTiLnAJIyyvoTjo37dNa59zi7lN6+ayBG4n2d9DPfbzwxIxR
yyQR+cUyi/RLgSM/ozN0IDGIZto7bxlnoYpx0OTwNQGyci0GDai0v0pcu252txySlZmGgPjxP3zz
a2y47GE2wgI5srnAUN9P41LC+wEA7xZLWGmzSklUev61DabNR8Nb7P99OWhkqeeqPW1qz3Uj1t/j
rwoUfq6V3qdR3D3Tju99HPgKVDf1HOUKAPXm5Ff2kl4/uX5MqRba17hJf7yeaWvz3Dq09oVOxqnR
nCP5fMARa50l/q4rF7FoLcTINhZPxQJAlT858ycPhgQABJeg3wtqW8iAj8y6gRsMZw9r5Iz8d1ME
oYweCfREM32y5i9se1A3XS5Mbl7WI2PhRNiftxQx0la4CVJMVLyV1EQerLq1WJ28NdoxJOHEElr/
ZqtMF9aHVKQUirAKMX1nvXWEJnJF/lAb+qX4rLX2o6j6EMDTM5C+NAWUv71fEZ/5n0/GcGpiAAbL
WyoUZ9uSynszXKTQkWVrMhuzru009YOl7/xaYthn8I/90lH4q7sIYKJZO8O/ZQz/OF7a4/4p/Qw4
7xs9gkHWR5dOJdwn51eVBa6glOiVYZk0TRIZY749Uwmckw1pNlDFGnQEGF+J7dq1MA3hYdxVhyVu
xC1qnrLoOYeO5RSkV7hG2Khj/ims0WrJ5PGB5V5yOH6wN1NSBCzbcoXpCVPcIjo4YeChVU3U5Nl+
v3BHt9F3Nfwn9O7KjYlnGbdS2PuB6p2xa0fcUxdM7EmPKQGECFpj1rJ2tDe2Rmabun5oswQlW6nz
q1LTx7JvB0ts0XY+3GYkZvtIFMU7X+Js7PiC0llK8ZOxIqdCTFxpju5k8aW1u/FVQBDflNTco+UP
3YFdwPp/2w8dAaZJwLgQNqwDgFL+DWtP3m0bY/hXxSTIJ/lxUKMqtpRGCtbqc0uKnabbF8qcYBge
nmKFnwmY/rNDbKajz1Cx+4B1hrvqcIbbK8H5HIkjhtGFljVUb+b+4jPu61leRXG/OxWNvytDIxp8
V1DKcD8TktZ01I74Bq/GeaSGk4tzEuIzYf0/O/ZL/TWi5GBXeepAFLGdDo/hXdnlaWFsdMA1XTj3
LuHbOBLY7SY4CgJbKx01HtzbrtG+pWlnQXPQCy12/tRywQkP71Zh2BSsDx5FE7gPoylOER00otmX
JoL/UE3aZ2HaKgSMHxIy7I/Fq/k8gywMco5Vgo7gPLWfyDZU3tmgPo7rYgIm7GVv4u1ENzsee0OP
TaHe/M7nD7uc5sXAuZCKuBA38WCbmnElzIz2E1951Y3lgK7xCEj7IUFUIpTG1GVdIRPPDT28XqEN
PmGOnvZw5gS5nJFpQ9TDPVXe8WrjHvK0gEFTQBg5ISfZ5QcR1iY2JHzV45WhbwSiXcMz429VE9mR
XjSiu5LQLuM5IsaTksLFtt2hNOPRTdqEyDxKI/HeZBYJWPc+14O8K1hbu8dgXhiH0aUPgDGs5QTi
SOJ75mVx26T7a0NA+KY+pYPGDVhIq6ulRkyMvTIY5NyrrgSJsu+4aim7XUsVClcNpIUpTOHIHlu1
fotpF0GI8HTTZzfeGFAIEXIev1lT3LtzdOoAbpyB2NZzwbABp9Ldn1xWOXigZ5HZM7u2dNYvINOq
C+3ifZLtyv2H+XXTTz9fzfG6LysPBlyBHV0JW5MJCD5Rr5YvbRZExp98aUzRviErKuxLq/8oNZqq
0kTvNcKztHpDnUtjMB4LvfAvxfgsMMWKmPnlAv9kTHTwrsrGLX9TB4r5yuQE43L2cFdvyYDzSIsT
n5L0abfg+IFZMnIzFOuAmsiM90IZL8WYnDJ+RlrqmZqQTdABVCMil8/sidVzrefLzQLeraRyAC+p
OhhuyOCdbOvo+ZpdChfRWvPclj1GsjGnsxEfCSx7Xl98w/WTwkDEEJCs1wG1ELSiUUX8KWfV9HSr
+XNEqoSuJmuABGcCkqFzLPsW9wCAXlb71DYLgcy/q4ZWUD7b8CEkPSpFvCO2d8dj+EpugSg7t9tF
ks0XSIleGHi1zNhykOPX+E93OhGWg+0erTbg1WRgn0B8JlpPpja1LLfSQCsy+qOYhzIhUZjKxuD7
HBnkljlmvHNC4TKieK8NiS9VDxyIrZQbFrP05ZJVxX8lbD9qT/evAz9nfuUAw3K3Re3cr0sbKg0D
5rbCK4LwQ29ntvQlBnmB1Z8rtm5wROkGg5aVBg7RKdNj5cjMemetNdu0esY/4cEGQrcueDHT/hv8
OtGKpXqOBU0a75P6cuDitb9Z8LHaT3bTV+iWGwz7PN/mSalBi6+T7fq91gJGo3A+qFqzcFvgmuzl
8QSyrQWU31AuZkpC6U8mIeXiF/wF4BDLva0MaceuSWzDYSGpR4BsO66wovMN9iHT77bELA2Lengi
0i7IndHQW40gxQYTws3rRJqmUE0EELQtHE7d1ezjkiCdB5+TJ7c8tza61W9BGlMrFww32dEnCfsk
oclGxcN1imgP921AfPJtL6ciWxMUBcOitz0wHvJWvd9y+g1xmUzVmM/aQyyyxwnm6rbTZRuqVj90
g6JGFo4KGA9bsbBv5u80LYgalG1R/x4oZWxc+S4SnXxYOcwFsOj7CGSr2Snj6YMvNij+JusbV8jG
2hunf53ZsJiDI/MFJCu5ulaooL3WfKGFeDHYlkmP4vZMBtJnRibNOQ1oJsTUdB/1V9YwuWIzmdAw
twaFuGM+ELzDN9zep+hd5wir+6hthhhlPxvPmuc1ijbShi/KA1OEU9R5pWuhEphTTXeQ0jCaB+g7
O5x3ZcFOyWmm1tx2aHIkikzXdaaN7MWh/cE/quNisD39sbN3kNBWahNyt3XnMqeII+aSJwJ1CcTR
+VR4eSgKWnjlV1EuSTb4EMewoq2pccdgVcZjhf5ePQAb4SCH/t1Of7axTd+x0ByOALA+Nf/KomHz
W1FXLqCakPqiFzhfdIH1C3y8lAdrtZ1Isp6RbBH2PwDPbB12hVk1ooEg9gH2rp2lV/i1/TFN+i0x
k6ne9aYTqkc40U5AuZohaWigAS6Vvpw47gpazhCYogLcy7g9bCdkcdWM1Te7oWCG7H0qqfXiT4l0
VNveaQYrJwBNtDZoNnS4mQ8Ek94fJBuGcC+xINPwcui8/+wSiuANGaqgg39BIfyacJUjuUitEfRm
szTGC9fhBJ+ZazqkLkfuN+GTidvmL4tUK2bz0Qs1j8Rh02/InNwN+YdZ9JNxZmZOsbRAJu4BtYJR
qH9WIiZvyX2fylUANKZFtl5pY1mDYJzMSZ6nW9Jp1ScNc4XaPFj+pfOh2Vo4NgXqAJc0YDYCYBZd
E8FQmLvScpndC8hYHvZYHBoUvZF9UNwQOlApJFkTlzb2HpB7hqFR/VLnZlMso2r78It2fFKQDJis
hogZ8DHuupZg8PhPA4sOu4P5OFDNIIi/+tGaiZ6i0uKLtrbxJ2M+9O83BpU9xQaMHIw9zSsNfSWT
tkXO75UgpubABa3QjFu9eli8hBM2IKXcyxicgB9POj/tm3ToBXHTwR3tEPYkZRm6/jGqrdTVmOHN
6f34OhsmW7X8yTzCKACYrMM2SQ+hApIdZi2Du1dxPpRhdRYy6i4kS6Pu3ra8JMva2p1cRd/30+Tr
j73ultILxzdaJW9CdPMdsdD30T9mMLdrBl4sMtVMrVx6dQbu/XYoXtCMCqHe41tFcoGHCsR3Km6T
mqdQKFNhJINfaKg8tW4j+UZti0WeMqTwGDLZ7+v1WzEOa0uyWKTTBxOcb8C8KuzvTT6cddhhsTU1
3f4XPkKNsFCpMgmeg2IWYlU3cyTJjuhfyxkFfuZYaUfWEYFkA4Emldkqwr05Aeqp2zasPAJVS+D6
y6wE6PdTNrx8iOObgiQ/II8kIoUbIMyRnZsS9W2JrxJ9yn9eSmKyXdCRQa+75l3x6IvqRTAmER+/
Y8IcCZL9nEaPJppoAPcjbJg4rB2WtuR0k7gLUZKVQn6uTU6hCyYtBo5375RDcGSwCauZZvcUAWYr
myizCoFle1iafOC0t8ZZAqT+cGRnUhAKUgO5Xn2KD3dTT7qILKb7xqwQVUlg1YtRIgKUdCWtiH2W
PvpXKWJ56Ip5j+669xq3loaMai50dDFoSsXrlxejA3yx9lgB3e0VpZARj81ffNGs8nG62RLIgzsq
uGS3WDXVwBb3jDDiZIMa77bNJKVaYTyoP8RxHTRje/z9gL7VeIt6JvWdm5K+w7GL4cLxXN02yiS8
lGt7G7YDbfbohcTgEAigWHiiZksb4qQis03omZO8py8O2CLONaO/M3bp0ihcA1y0htHdKUHtTN9+
Qe9V6q9wIFdxEveiQ1JEII/41JB6m3QKmXbQJXolSGGGAEu3c6ju1XFGXhsaJCzLTIuCLl4Cjb9i
lMQxLDQ5fXQXo3gScNLfWT4S+AsGG/tttWj9plajQFUlzjTX2KYdLDQKFjRYakOnysP2Wun9V6/m
yISfTIZyRyjwVnyhGnGUB4nFxe4uNMb1LCodtbmulvZu7/88TpMEiRxtQBR5jKPHwMHdl0S5FIB1
Q4m4Hv+z2ukSjOo5FTCzrpo3LszzKJUTe3wZtTdZflztgLD6QjpXjICEQBde4PEXYagCHl3tUrEH
YrO8x+9hDh4bGSeI3KN9vz0+D+uCWM2IDNT7biv3gUe4+yUYRniJRDorQkhjtRApDmBiS+W1oRtE
KVhjRzzk//7tDXmiqD9mswxeKrepfzPQIz4LXF8IHfyIoZBBCFnsKHg7ml70xiH/1vs8pq8m5pYz
4y5e74SjUQbnRua+Vipv0qz0Giq+elXhIZYB2CtsFHNaem5C/fPMqff7+Hdi6B3JI8hIOysShPLi
h/eT3n21MrjIJzhG53MpiR7FlzFBbixxEA6PVPfOnxq5LCjdwIVRbgGpg5VsyHLxBgNUe9sRFEln
nN7LGKLFtZ1M67VmYRiF7CNUdGPFmEhnXKB74wUjlIapPi1vkO26vSTHIjaKgKCepA++FqCJvr0b
xe8FO4OHOpL/kZyqvkUj/Uz0HLN++eLGhoMMX1VJEKJwWraKrJyurcoC5UDqlXf4R5Ot03N3uEVK
s2UgqsCIwB58vkKO6hDHZbcAsfuYg1CeBOieXMEZ3fzEcG9UqRl7A3Zxzj972bV1K3mKAMRs1Qe/
DuxhQPpkBBnLFkq36AC/7tnZZk2kFJKQokqw5YXYPf+KodkKsu3A/Ve/Zx903POkGIAwZ/gqc6ar
aEnFg5pJqSH32ab11eaWF8jxZxnfuNUuhsO8wlpWkGdejopZIkqCkcAJbla02BoMmRbhV/r9uH+h
st03Iok9P2MbaIXjRd0m6jdwRpHzKTaLesxSf+JfAUuSmQfXDr3/lqUfSfLZa9R4Ts54v0+sussB
SaiZb4CfRTVohguUlJ01KdlMmSYPrJnzBSFjQKb3+9znv8EwkzpJi8FHZaOR7Q7huz3dfELOv6Od
KboRX4vhuVWRMd/UjYtzaGHuhqwGAzStjQ571I1UUcztKaRGWBary+rFHA3GlBhtvCVD4vV+EIWm
dlIh/VkIvobpjRV0rX8j5cmCJEdf5/XLvRytBOM7C0loYiHsZEgwF2mYD8cPBuuc3Tuf2XAvdXkl
dnz6H776XGnCLNPltJOJlk0hCyLnm0gBY/xFEiJhONxaIs5BE9OkatL7ynA88MwKzqAzumfXxYn5
bwzuEhd33vnaIdqB+M6gz+YjWH+1DrTR21VKbRK8w3rUgcjekfzYPQtJqiHcGnTYQkjQgop4DczW
59vj6OhX3trO7Asl8l/K0taZFDKiQsOEd3WZjwsXGmkLywfJ2IMStmiALkl7oLu5KN4XPEMxfL5e
8Amd6cDqkTcLFX3j5x8KxsBprLpufQvs6lDc+bmXg/cpTrAjz+gZSjOAuRoEZExUVhltjvEGnpuN
ZTt38btIEpctYqoR3kIvpp8HPhknzdc8NYysXoRJnPtA5wSCUOvLTr5uQOFMRuQpBLBCQXrvzu3S
KOBl/tEf20X8jZ/xae8DJ1/WEyaGez91G1q1NSm0bHEe/2CQZDWBsaQGU1d1ssGrQ4NHgdKeCf2V
ZB8PAtVw2UTIDcqgzyburklWA2040bCp/MdbbPfQ85T3o5xQ1SGX/BhvmlcbCUfwQp7nzjlCAayn
2uzYHubiftDrYmtjr1bQUH8tKcXeSPhkaGEISv9JqsqKNHXEs5dHdJDSlEo+/isk1BoYtU+NwQ9A
RnCnytPZm/XlSMq5XEiWb8e6bz+VkM5H4uBU55D3ttPO7vBAchI1kfol1cQrf+ZGx0hFGNV5DO1U
FDCZ5CEKh+k3iAlXHgzsbntQJ/CbVq26c6b+lb09gI0jUJm6w9YNGj9Bj46S1IYUYGHSDIWPcL95
YF7fUCcEBDTefPdPslwUgVlmB42HW2Iy8E1bMz55MMOnvAmMc9WhCvglEawReSu4RX1lMnzN0uv4
hTmACTtJMXtLakgDnkUhMT45unJ2Ht0gUrgAgWr165+6mNavX7gSS3OVswPtg9QiHyVUTAhzzFfy
qQsyDASCFRM2r9Wr7G401a0gzSCpjvcjqcTdb8IeU7UOY35CkzZOl7VWbNi6j4oz28U7FUEMy235
QEgPhxx09D3pg04HyI5shlbi4IjVKMzcGIbp2FbNVGU6gtk9p96xmRdgthliplM3jZMvvEE8z61e
Y0QCM5/jIwwus71FVWQncBmoeKAu9jLRaOHHTej98z+wboftZKdjX4JGPb8fsAuHVnwewKS2JBp7
fNpEUtBZZF7luWgS0ho7umf/1bee/4kmk+5n92znnwFBIzLMCyK/hHuWPRW+TOITgIc8qyOwDubW
oAwdqNk4t06KD11oZVFqJxX/hKHRcwdJ/a5ZCU93/yVYBT0SN+avFEDlUGpiIwouqrhEvM0E6JjM
TV/oF8TuEWy886lzoyshfamBbhK+rMfQLiaqLTfGJGeeOLFB0WknAPAZoUvtPgIj7VUGfA7URTfs
vn13KOJKmq/AfBhvmomPyxBxvFudvMxl0xKkNp21M3vgsUh73/joBf7jDgblpLNduWKzSxx7GX7E
OSXmpyHmJnQLEYFswaL2uH4PWe4tGrvy3pjSCgPmjeGQ/tmLmS0IC/5pf65mjhsUIfJkGxvXOCYF
ScY+l1TqPIpxD6PsQU4BEmzFVM2XZz6rzzDNS710CA5N3PjXggzcnvnQUeNvSzoWd+0DAOeUklhN
/5zga++WB32SMp1GMEwFfPJPqbVLeZYKGZLIfVF3OnpWaPxnuxqFApTHqFSyRQMIKZGLd7uNU4se
91gn9jIx9DopkIltUsmXnIGxrwXTfAUrTJd6+75G+w+Wg+x49a8Bnz9p9rvSaLI46O1ZkSrZFrKQ
/c8ozVdY+v8MfYbDSyJhCI4A/bOTK93V+rasHfxHooJNcDSUZohXG3N+9Zwcb+wl0A+wkUBOU1LA
jrjwvAwcgNQUKsX2J6dXsOH602m+0hJUoi4z9eSRaM+p5eGi7Bnt+aWg31V1KrnNFX+TS033xClh
dWaiRtV0KeZ0C31OL8p/FsGWO+W0/gLxLnpeC2lF7Tdfq/nq6oGWCZLvy4LCUO3KE52Q87Lu8Q1k
E44wl2Ypwcq56KTHsGmT6sguq/0cag0lfanoCCfQ/7qES7uLIru9HfkcextNhh11eT59CaNBExrb
QK20hmOu7amnh/xUPBqvM4sKLQk8PLZEU+mCb96WSN3ucPNYKP5/idu/3c53HLaZ3+KktMdGkNE+
Pf1keZdp6y002aug3aV2k23SMqZBxyIXN4FGK4HWwou1QHiSlQXmPzQ5ESmiS3dkJxW0E3CLazSW
PKviELFZD62NPwbjs0gcWhIgeAHJTFvfu9jiZHRrbH7zCcEBfD2GXmQglEl/MWBiEG0QigVMZgoa
/prDilcQe4K6jIltBRhwhkpVbXPt66HLE048Q76IblNh0DO6MyqPz4fhBQk5Paquo3O0UoDfDAi8
gdN9wVVE6wou+QPczXUq8fwMV6JMjtZ3Qz7lO1ckszJOU+VepF0XQro5u28ScC3eIRd+Kt2g9P1I
yFNM4hRouYIv3tvOazQli8oTOjF6kjCR5oL5GUemCPbFVcsE2YDfvEkOmQ7hbLMOa+22Xc2Jg3A6
TwdkcMrSJO83GiKmoTe1qIyrplgKQTwhFqae+UuuBt8ziPN4xA2MHCREKySyRWYGOBvB/8nQrQkp
qCiaUBQg2Ig9Y5Ue4mtRdG5+R2iNZrLVB9jJ6Lylokn7ecQlzTkG+n/gysl9ob2PkValNe46dJzi
b4pM2X7MHm//FgiatcOIK7EMheVSK0vhjj/BW1TrFe2+Ldes5crF4MIjFPsEu/m8qNUGLn37DNCe
eDYu3XBF6uJAEYqWvkCvnrctUi+xUWZFXX4gJX7t5KUI+9AIIHbqVkNayiBebdH4IWmhwkXT030p
U+563hnx8TuMO6MIyRINVGtwIdsvIdmvT6hwJE4iNgEsrTeYoPaPw+HRryysWz8fwI5/mP7Wq6+9
2egV0bbfrpqdgKfLbcOMDamzj6cSjTPRbTkFsJNtnWCFf9PCJV6maQ2UQcA+8Tl5HsEu7Zz4NSZm
/BD4sFpMqaFx19NeP2BfIV0Whd8N/KU4sUXZ7FIG+5lpee+TLuSqyI8zLmaTtnszA7qdqzN12S8s
JwudfY4QDujyn4UQ2YUWga9+MmwUR+48EaMCs9nEdtHLhR+Ww/g8svFktuZ8anx44dpG9b7wop4Z
6WdqdPOG43slbMTIBtcANEJ/SjLyIqRPyps/IJP/h/j1hXLidQbWof8TJVHaBTi1OtXpz/QBStK0
7XdoxKvFfy+FpuWN12M/m5roLMjjOY3QgKCRFTxn/KpuedCbvNT1QO/YckRpROh2eptywreWSfIr
+7oEow5/xjyLpCyVYRuvhpdO9L5ptiS2HRp9c3hDzn+OxfnbNxtdzJjshku2cXs+ZqcvhGKaGCVV
olpQna2TiKzAjXIV1zwZIEHZ3u7sjl+5x77kW1Jq0y4VTGIzbsnMdzl2wXEUXEei7+Q5ME8PpEBm
Ny87HacEXLzON7GOhx9O7Pg5qwzyO3j02qotCMz88RQIkcGEJG/eoKaztQkJzHqMcSMgyAcZo5W2
N/B7/WgY9fG74Ob5wBuszElXA0jvBRUOh/BqbkG0kQ9dF4L7VM+t2qs9fZUDCEEDZ1Dk0XZDpmf9
OjZ8eZVe/TVslNaKcWoi/7cdURcrp+T7qxk0pNufUgXnhPLFVqZZzd1NI5okYaR7nstnzdnTbp4i
zR/g34fnqN3M58Ifh/URKbIjCksI0WmYSDEBgOU8aM3+lFV+T+jrhnW6F8PPp4CngiykgTF7iVem
2Om52W5kgM+OrFUzfB4cs9xp4Yj3oTCvC+ENj0uRS914EPzSrPhzjsCMTSTRvRZ6zH9RxBpbd1hn
FyiqsugnG1UDVBn0xZHGPhH/3svuNPEQ0sQv7tjYoUx6LmRrA1ruwtKOwxi8XYz1+gzIbtMXMKmX
Mc9RugfmWRTdjtUh45Wrfr7RFr2Ee396Rm0eX+w5QnhC9To2wJVkwiSOgTGmiocO8jl85w5/yMcH
ziA0kkjDfwpc+Z+C1x4go/CsDf/mfqSL6JXUBmC95FWqNftBC4QelUN4CGYvf9nzIMxqHu33S60s
EudJWwbBeUmevQxy9VCpjpxQ5dyAnRSnpNrudYYNOkmU1bgmrrFTAfovrlY5tA5hGajVuZ48JbfG
tECfJ0Cy33KcS9ld8Fhnov8uYAZbF42TU4jPY6qBSOFJzfONtaw49C6TVZ9fF1roN4qqnPoitAf+
61S5aBGl3P2LNGFihk3gsbTGk+OQyr0OAn8ZazrX/M9wx3QBFNbkosr63CtN3GP9E0VmIYQzUADr
Bx+QLBnv3cUmtVpdsVIRVuTQQoYQv0qUAxfXbTwCyPMZGdCE88UToIFuAxljMJz0ofMd80AOChjI
ctDkhNJ65oQj4o2hscUFVGqaP7iJv/onQ31lErxTpZxSvsu+szBrBrINYYJ3g9JtLJJxuaxT2+kj
9nwtp360cBCPrlBmliAwcWhv+kqbMloV3vHjQqV743IcqUuVm20nrEdQoYMSsNpjlLzxi3hg9eru
Q4TkJPb2nNjwGcHx82EORk3GOwiqTG8DUcokqtDXYE+kCi+TSTJ+O96GU7AIY8+ly/mFoM2zQtFl
mJ5Z0pnKLslOnt6Por8VmW19zY5V7At94qcULeTsmdJtJHGcg/hKfj7fx93/TBkUkyy9vxL36Enw
Df+DwNIXgKgEwOhdN+4/B75qZhLYlzV7t78eEYm3DrNkfk/7LQPT+wG7r6IGatC1zfxFT/uo6jeh
MF19ANLziofkn7ezYju3Ajph277PsaoGdij1c7dlZm4oWPNCyn7i5vZr9DSo1srYzzJTrW4y6K6Q
xAFHlp1te9kLpyRiyddNp0gch25G4Y9KuXLZDO97nFoMMxSvTIGkH5mtTKSnG2x7ba0mQAk84hrO
81UW3svTOeo9c3KVqgzp3IEUsltCWkhjEFDAu2wQvEP9r7dV7mrzLMR+uAJTMqP4YY/hhfOqBewc
77w2PY2Y0NNFavNiHEVIpNrnepko/9qyD9cWk6y5gWNgvDp1lXYjse33wbs9VHEmQ6QzlZKEHzim
xQ6IaRwK3FvjRIOzS9yLxKKerI6IEN4bgaSWTqQM57OZRWgpwzxCGiGHaFhpoWT3cD+hWvjC7N6N
aefdJ7vggcSUwxB8sLhPijQk51ov2LkZ22vVOJXbvaFCX5BBTrR547+ZH5RDladFINKNT59iwA+T
M17aCeBJqYybKZc87752vzyi8xn3ktS2qBN5CE1/cOBps+GjDtli9OKCWaRzUBcYo3sc9LDacFAh
dS/7QvnXLVftXUn2seaXyc4xB426RwGcB2Ir/5FYM49wbuZwD96fEpTo+ysyUjeTHiF5yTUxbdGP
k+CntnEoq87bxPvb2n/xV/2CYV83pRg8TzZ9yaaGzV68M7EqItGEvZGaV2TSh7uXaqMWIAeFuSMp
vi0YxKNd0WSbnyJ8JvqV9hUxKNRUtexfiCLn/FfaLfZIG6goGM4ucbstVuf953Nt066el3ND10fd
KAMdIotWNsL7H9hheD1ybDBvEsALK8Z/lJ/8Onq6ngRYv2jckjKCJiqp6EzQDvctYgTb3D2+UVge
NNiG+rSIv8PHST3EgAzlFC1ayGPPif6xRfYkywRZYsXKzK9VQZoNhqCrw/XQrIlPPxbgEEusxo0b
75eFhUMqaom6Vr01CzspK9NXoMe6i2ILNJm4if5kN66Sod3ZAfbg9NxDBTCNjaua08oJ72DVyiwO
QUP6U/D0ltOXDuTrdKBpnQIIIHFPj77HiK/E4X1SwmQDtbs5DYCGMZTXalqdVb7inc57WNFHeth7
gQg5bk+x3iXJTv39Ygtkuiy4xbpZ5CtlLgyjGAZVIHozi2iYQhynLT/N+g7ujcnw5pKqz1s2qOxk
71mJAIvyr4OKBtH1yO3yRCIs2Y8CRJDtwYPu9BB5RlH+t5LbU8gFKvi6GSbqmDdEZVLyNB7qiUZI
yH+zqQEnpL9t+3owTKnboHdamfNhwlfw5+dbCx81i+G/wlzqU92Ch01Cg0GKutrpygSKX2A2ZpQi
pFJ6Y4pBjj65UbPUWNYlo6zBMFb0bv77vvrZhIHdrD3P9YWL8G4VglAch3zAlbqwb7kPc0SPo9Zp
Pw2VmXQGrytFKPT3dmUckrvALmgusO8I6zeJDEUawZvGxOv3s9pPIEggFIfdKmKwVBU9OMu0Nvx7
JhzAY0LM/iUJF3MZlkrDDiAxmb52AJH/eAdLiObYgk6RybF6cNEZR7dt3ArjuQMHOy8qg7fucmhT
JvCTcC5JgnHpIjjArdSMeP9xzVXTCSC5w3jdaxxqKt16/Z61Aci+k6huxgGW6JXX6RuenFv4xpYD
h4DnPKf3jYfut9uT3tFcJxRqoh4G9HqbKjsUiBvCG6tSyWb8hvsrJHEzb+pXS9qdITfJ/RUmG6k4
/JWtPTNwkQ/W7Y3LQeI3sTfhkoti2FHV2O+mMRrCCFA3etg/O+9f3KESI9+24Cx1pcZYy7q2stvb
ZaxHCeFLRGaiBaI36I9j075gOf+YLKFIAa1/ItYK9o+EDO6Qjfmgleko4vy4VSS+IjLfG2tsyxHi
9ovaZxbJmpGnMPwU0rrbEqvLSVrx2QA8hzCj1MSuou0aIhtmjeZK4u29O1v9iAUo/INB0vnabgG4
vH6X7thOz0MfRRAm40cZ6yJExvWHybBlxEtFPrDlgEr7H+d/5yyskuIwyD7AaWpbOnpQFkHMeTWT
SpYXTY5sMrPLR32D0e5o7ShEs0qpUASMClH82Uxn8jQp/K9bVjiZ/p+bGKOMfsmbCDy/SOHCZHNq
nDj461VuDeGPDpD+75cwu5iT+soo8SzFlFS/tmCUmiK/+La0PxwSUyyo+d0lHGIfsdTuysYzFt+o
Xk2dVrMa+9fomx23h/PllbZ/RBXa1PqivQ/HL3Yc4pjH6wmzqNiBqx/fGL3KKmsrh0s14T1nCHO9
KmvVtDAp6Q6JO/k531Rbgr/DzzoyjEWCrIFVtw8gcWWmBDm45Sv7QRcW7bxaUnB2F+kEtEp7l/Qu
JiOXeCy9idlzfKhr7OW9j0aJyQf4BgdTrdII11ADcl8rB14gLFnS8c/2LWdNNya/eRujsJhAVtup
0/amnxDeqJFEzXZ7rjcLswVzFZnp/LejcdY3Un2prwR60d8tg+IbBfux1u0WIDeCfzowvIO2i/0K
slM8v2aDq/3P9Q2j6qLaHIbjve/Bo1IYv/UU0xIW35EiduwtjkAGrDFuIU3x2FfZ6H5QdCzCFpZS
KUBWZ2yY/lY4fG5s3Fc/LteBJ9ZPzMOgB8MBwLk42QWhrvXC9qxlO402RGyQG6IdkEaJTzT3jk/i
OK4eIXEE6PxuQz9/S3+oUU2MDLFRVGpaa92ZkCnTr5S/ml1SpdtBA9BvZVQELz5qiSROkBGGqsV5
1XBmEv/lxcIUezBh7E4prVmklEnH0iHlS0tfgWgTc9fBUNxCpBDAid3xB/oVtyzvqXc8zZnU1U1J
oLnvyZncFc5ZMjBJV3w+NK8pwk+27SoLmrj9pZWqhzJC7i6wBgbYIGVfBwjV0mDhNIFbt0Bw19+y
SNTc7k/1qPmNm7hfUIifkHll8sAdiBSs2wfn4YKkfJ6lhT9aDcJN69myzbH3n7mtlN70XorjFAte
gAuCBLjSVHh4RAVncXojDt3NTWB0Pr8qFTOCgGuo5qmI3q/BrkVxxrUSu1Eouw6hstV3G8FtVLS1
BZXVAcMsEARV+FVlum/K6EBOQBJ2YWN3ZTUbMGW6z9rsBKTB6JqL5Adl0/aUH/CnvT381XunclK9
RgXeHQsX/EnoThYJ+0FgQ77Ru/pf/cvvqKDoUsCRlpnmjUXwHiUmzQPijS8RFfcOTR5Z58MO1z8i
rY2wXBdnoSxjOJ6iGlv4tBPcwC6Oy2aKQ30x3aCGIgBKY8ub4ALedX+sSBWIFZFw87A1veiCeAsc
KbnRDLGNcaZNGQAio6EOUbAdehJHU4Mde3Lb37LTnmpcqkUcjmU/ulHX5SKlN/I4P8a8a1lkbSJE
E3GkOFm5M0O1MWvwpku2VIDVwa2KNOd4xq0IwIjX7DzzEGG5S0fPT3GXAABvvjtgOmDo+7x14WMG
Q5mRDhEnCE1xjgOHwJNy9x0uw5G3qpwTRF0H53yAYBNjCzNVF/3vUTEbG+nkUPqxA5e1Iuc3hrQR
Brz3v5/2evrE8foIN4n9ilxv0Zy1Ew6dpADBlYZzn31n+ZGzsYk1hzvN32CRjFETvQCKZQpR1yeg
rqWyAamNnO2KslTjXoMfauW4af+Qa4zp1d8/UAhNG9OaZfmWqPSifzMg27+UN02jFg316UB9vImE
/ESHgkopwURwpCpbYfdNJWwaVwV+VbnaM0tfmPL4X4CBoH8t4XIngcemv1fLSCEmnX54hHk7qQYN
BfB5NyDfziAo6ibtrQh2/W+It85g6YgwGqPU0jm9HDfYE8Crdc/2WfG6qU4Kj3lRHROezl5EfWg8
8d54Vh5e5ATaPP97Fp+mUqVUz6l0B2+46f141gPzO5DrPq2n5GWcobCc9qUzdmmFEkz3XncAVWUd
OXvNw92203VI2M6TmB95TOpKaTTLw+PQH2hc8RHAsv+KKgIysgcBGI5nnIXdvHqGP3XCTnbxiS7Y
Godhip/nP/EdEb4mJe2+aUndc0SrG/OwGjERB/+e3MT2wP2z6qV5P52wJHJhzsHW07KeaC/yeYpx
Nw40TCiMkWBIFHx20lljj0/ju+6FDQHBFEPd1xYiATCleV3X5y4rA4M5LJpKvVRz96xYN2JzVysk
f/kHEdqhLaHyXmNIx5s5epsY9B6djEceJL8YLj9TFbDqJMzu6elpAQ1RvCQRY/ii4Hgoi5TOYOwF
wZaCIJAKxDJG+EUCz3puENYy90HzGyXM1cwSSltVOedXc0eHyTCi2edngoWeNnD9J/jQzhtCfM8w
DfISKzliala3Mr+xPreO8x1Ma+C7Lnp2gbHjw7JUmq8ElF/H5pywRC2echAs4ceKopb3c5PHK21R
KqqCeIZBITymr20mP4HCfwrxGPs5Jc3Q0ha4aVPB0bgQKfPcirFvGWnhiAPjxZXb9AvsooBvi2QM
bUR3rHuJuqloPV5ieUmB+h95AL8zdNNjAntwim4XeBOLIhT1nw6CrwRERMQfZibOVn+WGadcVypZ
8kcZewjcQn6t/zWGrHYYC5NrnpXrAzl/VSaOHeJ1IZn9r9usJu0y2NXlW5729eXvPt0zCqSI4lxG
BF19/T77fM1aZwvE5QShsW3pFYVxNi8nOAek+1ME1QUVYlIePKdoLPNaQ9hRvzXY0MU7acR7XsJu
cmgptjavog8SMRUmAaObygklfEuKit7ITh21BnUrZjrtXwFk4QT8jbdYdIBo9pMOw+Zq3U8yIrUz
cv1brKv0dhck1idy2dH8oNE3YHK0rr/f1KwRlvuT0U0Tp5PJw9RVTJWdWxWSgvvKZ3fKlfiA6PZZ
tC+6fc5PqBVNt/CPNe4NxZaOF6+Mx6hXH/gfYa8CiipzHA3ZaLxnFFu5SaGfC93SST+u1/FD/XGz
pg5Y545+NZMYNnYNIEDER1gH4jzV7DFu5VBHw/7diGbVi1sPty7zUJQzwNtQRs+0aIFR9fGoXko+
jgKRF2sV/w7S4dVJipRswa4Gz5YXQhJsTPQcc9mQFG2ZqJQ5sz7dLgMk9dDkeoxGD77bTwDtNqgi
Izg393Xu6dbzI61Hhiz0p+j5IPORes+7PLpFQMs6Tocx5LH0d1UsM4CQHpWWlwMO7BpWWsSE63QI
yMGtIXgTH701SlqkCRwDCFQOWDkSu2+X0Z1Aq8Edm6oaeHZvkMhJ/NMDb2S2fr1AZqm4KVLG0hG7
P/MFwQ+U6N5Vt9kDR77yIDX/yBrD3HsNv7QGHYbewfDFe6HW4UhPmVaCD1e6Ebk6wTb6rvrU2IEm
Wl3cNS1j9V6yzuEQDPX1ws6UwRsesEzGEAiURzZwPp0ut1+HW6ua3l5Kn+4SSZwA/GgQv7gKj3hT
mQV+WKV1jOS/RSpR483g9r2OISPdnSyQGQbHtHk2c1872IvgucWOKOVmd6RWLFYc1MzmE91cCa2W
hW6JbwKWMeXUoSuJM7djgDOpbyXUX4stfbSyV8rKsdaPCBMFFojwxUIYS9tlTbFe3vP2FyL0Lxcr
UqkZo1gAPsrGKynWQeodztiaYeIJIRVIHiDUzmwXkVtV1OpqdJGKifTSmEPuRs4TrBOl28LuCUhW
x8j0Q7kipm3kpzdkgFE2zICdEoXtv90DjUAl7KlNrFUDNAjjoITu392v+eRWzfW3sh90/8C6+UOM
9GnAQXDMblJrQr6/oamyX7zaLYgg/X+rzC4vOneD+ly3akAE8YsOhOwfITuin9BZPLNO8xh8ycSa
rkrUbNiUfZE578YDqo+kx0SYOGzqy35Scb9s0Ul4wyna7Axgq5dzq8pYw6Bpk33rJAsI8l9qukmj
mfLsr64LyOzY8ywvLB15M8CSwQBk50e9WM3b6QU5eb0hCyA5YJBRFZJ0BfOTjhFRi4uSN5rc9LaE
8GT0lFrmxhG5uofvDjc7j5dBJXK0lTyEbVpRYis2kcUBQ5KAvaadmwbql6r/UfMjf2/FZ/n9xpiN
VtNUKwWGIZoYEodKDe3HP7RJxjYN9XO0ET+8epWcQSj93fI903ixC+3pqJanNWzUE7KWHbkm2S7B
ibHTTHOndGBn/o/NMtmZAZw+L082qr7+JsWAcF2pKt752AMtDB7py/DYeIbhzvcVDfz9QH2ulNGN
xDYuO0PmvSTeA5LDA+xQKGVirHzEq67z3TvnEdBnIWsTtvgcGoFfmXQUzZHJiiCZXXkW0HGSwdnY
Ekhi36zVWM9Yz+CPHUzcefIMDeLSzQmWakHpTkuwJt0CUji3UMwonVI5n7dhmEZ8Lz3KLmX7dtah
+FqIffhMF8eQ3H24cMKmNJ7mTgioNsrgKng7TgR3sNlS+/gv461hp6XLh6kcMlnQgFm5j/8mUxO7
Lk2ROJDRdewgflsHChiOPUIljl3KBvzPMWJLPr6UjErgxUovD5z1UAFWvSbAx36YxUjDI2YWwoON
wGrzoqnHCAARMfMaRmE8fxQ3wYnxWV4Zv8l8vju1qwIaYH0kj/rIsfkc8UejK+s4+ITnTP4JsDt6
N7LwtZ7kKnllf3kl6O0lzjxGQi95hWDZNiZV0Ndp77o+odlNcFUxy8EnUXySS+/aNl4KupZLS0M+
2Wsv7g/jXixnSmdNjfo9pa/D9cOeork5r9HFTA3AbJuhtK2zDZzl8oDRZ9dfkBbS45PDq+2E5E2l
axi+5UNWXKWbXgnRrAGhBbYXdpVLU6r+Ra7eORVFKCVQY2ZItxM0S7jX/odx1jCXraMkqe1JInZ5
ysJq6OktvyKDFif/d5tX7xFfSbhEaQXEyECi0oGxgSLrL8Y/T2b+R122b7ZPq4xmq4+mkag6UiWP
nE72KYNrkvGAs+NdkmMXTCAVg4ogi3tadrY0BrWTsR9i9fU2WgC55f+9ziW63PuXLQPzqb9RBY+d
9gg/wrR32dVHCiBy9hegwc5y8/1FTS0HtShoUSPd49g5v16gshq7inoIU8enIGcfcW/m0INpPWyA
H4mIlj+2p6cuWoZwqshKZc7CIHHPRqhhiHvFTvgniaRsUMpeGhChYBm78IAJG+JCg4GixPS3Vpdf
fBnbl99PzKXsHPrTEzxdjMnIreevo6GoeGoao5PAyfPXqR5216xFQdtkVayMgUgMXrT+e/nM8KCc
LtEE4D9AC+ZbaaRW/OldcwnJ6VKO8N9d98A6hAK/dzfynGq+2+diF1Vv/7iKBWOG9P4oU6iWd0GT
S5gG1Bs3MR0733+TbSF9wuLSv7R3WW+hEsuX5wYoISNS6rMGnpUf8P93MeMOK44a+qji57NKsODO
ORIudx/4nrO5Q03y4k52TQvRp8KXzvTOAQ5n6umnSZdtjMhFWLckSDSQ2xI+UxOiaNOpjB68OUAI
I1o54hHnxaAZp1AWPfkQRW/sGLJWzCCahfCiWHEPgG/fGEP/eUM4loKQn9QxysAy31QiHsQa3vFa
a3tCXG0Btrkr/G0w9C4Ieu1W5h2vMMrD3rCgibezE+334fziF0C8LiL1/d8BoNq4nnVeVj/mau5i
wgEfeXtjJ7c8oLsxmAKlBIkYcqQCNb3Lvr6iEK8mIOhP3JyRY5bsaXkoFPljExLFx9fKjk1yESbw
Sqt9KPQ+bs6TCMVIhtkIWN+gkHSwe6c5Yuiy4LCzLPP7s56J5PXtfJjNASSWUfc8d2PnQKsm4BSa
1IF7tTHBYpn7zY8ncjoOwMXZUcXfjsKhky1rKpDkKWHvAWI/gXUV7XPudaFv5jfTEa20YDXNIygY
Vd6QbX+54Ntj/yJwEJua55QbyDWRpdR8C7nj3Ig3WRI/1KUgQ2J9TUn7H8ae6I7SwOvv5518fmcQ
ITOuV6uPEiaHMo20TaOVjnjE+/wl6tNS56KgCBgQL8e7ywzCb6W9hulEd9ddZ1CX3hZOJpsFFkL2
uWFe0hBQIbM3Z+h0QJRYPEsj/8vQykvzbD/dvhonWA9K9yvRxzbeacXI5XlAqmTz2T1VMMJFZHl5
+oGRWA2/QvSNcsjxZpwlUawRfp2mLj8HTIb5D5hXIMgTXG1750Cp7S3shxTyknEI2nMas7CmMu16
X8Ki5TT498VZLDNr6uA3IOSI8SXKIwwa1XqH3y9LgrQ8zq9oH4pP7epSBRNVeJ3xtSkJ1On4mgfO
5DzBLDcVifUgA4Pph7U7T2dByxJAXN6D4p6+eJh8uKmMiEU6/GWryICMJI5QTBuWwD+vScrXDS5S
izV7LfC4uP/lYk21DdxyoZ9mIJIjzJIyFB/kMihZ6uVkbNmvHWz8a/QQIgK9zXEpXMReOYoQBeex
Qc54SaKNzvwwgzGu7zXn8JMDaroyKz+IqlG1LLbCrVwQbXSpqok6hSeeG60KjqNI5Jxk4/bytTMN
16bY2AZt/PRuBIUbKP21n8UYO/DvQWiuF2p+n1cfDjk4ZPI1xctNWCTeEK3mTJtluqDhy1+tvJJa
p4J3z7cd6lyWdB00pRfJSC14OdLaEJkt+tmlyb/icCsMaClcVH8lB4zfe0F9z8/NtDEbUXarEq9v
LWBLpXn8lJyztaauqs0nff0ig0UwUC+KeaLfrPt8fca3gBThKlZW0ZdXefmXtaVaLJdto8QgEVUU
ZUMPal0m0eu7cpAfKaq2NcUqmcKpD89O3ECSXm/uSW4o/APtE0MSET2TOnZkJeECrsbvYWwAXT8L
r7ML7NHHfASflrZKe+rFFVhlSCNuQ0RVwmBfvf8t7o9OABnwYeAY+HOJhblj9FQpAEySBTbCYiwp
GrheIV2Z78uHEqL+TJEuusBm5mAlZl2/RGEneRXKwnHoW12efjhsTFh1YwR99dkkCLTFQYVXpapc
1olGRRSp7bCOki+dm9Peq6jYnnRbzKkcNIjvKl+DuklfvIsDp1eSAJhZ8SCdlP6G3RRcb8ZNGQiH
IrSnLwR7uPsTmEHj9CWJ9vdVoed4zL6Bcwvwaj3OLGhK77qSU//qz8ulTbyjcSVEifqBkP1ttxz5
5G19gQelCLCz8NkEJTSINlzo5FXReJmNgd/9ynRo/ZGv8nML4XR5TAJKqUIIgpmZ+yGEMsXtQGnT
2E0YlNI57dU5M97Yn0U5w+2codgjyxpvFqGLJ85ghrPF9v8+C1q+K2EM2oW8EJzAhDN6jZvI+zDE
6MLCYixm6KV5u0aFxylABtNiaraA/J59j6+lBbG2/kFA2SXYZ8+Obbt8ubUzH0aB5OQkct0rlxhe
YUyNe9fiOh5a7fHVXTkPS9aXOb1xBvfh613I5c/Ziq2CQpZgkJyQqobOk/9HHI5R3O472xOngoLl
stEhb9sc012fF1xk6QW7dypXNG3B7462AbgwXSItqhGnFiZpezTTP/PT51qpxv84iWZQ7mKggG56
vOO/gwY/pDQuVOxPjlfgAnugxaOR+zyMiXBOHICQn9Lg4eDrepWLd6VfiNUcwVadrE7geLtaNvig
5AKBPhK6t+EP+mZzodfAPxY68Dpaagfk+a5jwiUC62EJZOFwigyKjWNqMrX6vm67ZkyEUPDvwRY5
9q7DripAlhvohWYWcoeDo5HEfTh0Jw0cp6QAkA4YkCyQGnKqwvIBNgMv6/yjHRcPUumR5mcT8HRy
VZIh1Us+YDk7XYP/lhz7Ztn4fpjNSfynvZUv6TRhIx/J7UXA8pFq4tGlgO4J/IeB5I3vIEEAzeHt
Iq1UgllAYBsw61CENLjdPyxL0RMqvPtLD6CjlnMv/TPxUPT7NjEa3WgPteI0muHt9BlICr3f681Z
/sROSgiLMXs+kgff90URh3syyB4UgtiBEMxxZDKRQf3OevtqMOwYtRPKCPUJ5KNY+RGNpedLqlan
6LHQOn7OWb8H1O4Q4FCx10B9Kjh3lrMzcI07TtME87JRBmzx0Va7e4TCOjLkd1+ShV3pFW0au103
zsHc+3zDbTEqjlHAfZSU+z25m/SmEs2uUxyisUyHsruY7ZH7gYvvQZyjhZqT+LEivqdNwSoixN6/
mn4w3H4taSgUp1NSdXTGdIR2zNG5jj2jCSdZ4aPlKW36+xschGS95Cddci/dUuxI8oeRrZ7iwc/d
eqtDLVOxQBxkk2HEjq9MWpW18Nc121NX1q9hy2rY9JVI9zDm8K2qNFjTOuJHSswB32qi5vRvBwNs
DgVdvuPw9P3PUEgtq0hOjn/x96vDniUuG95rMhdby0/jWljYw+e/0CMud17HySPy4xBXCAp5GjHH
brLWkNzSO8mZ+chx1BQnhDc5wJBoTCifN/m6nNMvvhMzfupQnb5H9KCiU9HoxRHs+6FA6S6US8Bl
Oro/xS4u+7u2rjJi0nUnCuJa+EEfiPIyaeATM11QG8Phd5JrpRhz4uLg//NxydzEwB9HVE34Fb5E
svIXClu9iDa7mrNzro4ZCHfB6hgANnYTuTLfYQvqmsNt3eUo6p+MtbqaSLKRYW2k3YVJKfnLwmMb
fVJtsKv0JBIeZfymqQlWaYe/u4mufB9ibVZi6983atkPP4QPtGH9A4RvH8ysNninexkCkO+WbK2q
6rmJ5T1/03CY73N83koLp7FnpgZU6zskZXX2j30CwvTjtqxq//KVH4G9p34ntmSX4UxzZJdUN0RX
JPSBQuD/36lrtV3647Aq8b5a1WLaAvdWftnhwegFBHT/qgTgrIt0yKX83EIF+jUE0B+BaCpY7UzX
j8XPvzVDlfA9M8JPZuYypcp5rnWp+qrnEfxgs8t/sLBvYMtqBjrKn+Bu3cPS/TeSYJdWavsoOOZK
uKYlPXgeCTPLVcWJFpnN9bLFpjqlDeOlbvwh0oKRjJehSaYB6hwH3Jnro2pCAMu881FzHez1DcOQ
TRstI2ztFxnv2xkSWrOWEGrTSSxnsmqzwenIzHKa6BPacT7XnlNvzgCANJLjsqTXpBn/iUsOuylh
3rg0b41RPupvjNAlZPUAvHczg4DGaTfPvga+NUDZlFC3zjrRqfGmSBPOv9SwpNEuSf39FeJxO8Nx
EQKbbGNXOVTzQBIGgcJYKv2oORfrAFpNhDuQ2G6BryXQfHI4i2JBErZzXpZRsaYvHDQS8RPOCtaR
tDv3rNyq8ZTtzA1S0qq9MJ+UaiAxXFenG2A/oOvVmG8762/M+EB8fOROkaOtb1rWfPlmv/5kwmM1
bk0M7ZEtwYVyVU4fRI8agxtKEY7s6sX2AwHtleCc+uLNP8/nHSdtXkN9Ikt9uyZNPVpw/bqbCFbk
sw5iiObyyN8B08Gj3Tqkq4ekVqx+TIyxj7Q4WR5TST96sczcwWFR1lLZ2eNKnMlJmbPbf1kFD0XR
qM0xZajvD+IJ/1i2sU10npTlMvEeNuGTuaEvQDw3dyuVp5eo56PX2b8ioAhk/CNcmXLDP0Blfyx2
VsZ6E19beldWc/5sw16mR0AmpiZ3dEpf0h5HsCcvaqxORv4FOOjr1dFJDiEP5vbPd3adqbO7Mnks
hooVThuRF4W1lvUIt0LMmNFX30xr7cdt0xSgU9N2Wvh0i6znBgmmj1A5N1WiDVft1QkbCTnZYS9h
Pq/XdjavnN+xwlckC6V40wivgiIRQmY9/OkkAn3SrPQZ/KYSXn49a4CyJvW3xxf8ZVdVgAJ1Y15s
WQKgLJiqjQpJyyf3nj9iiLLMvtVboGShw2DfLmtGcBvSqy+b9E8Z9ywDEnMR4ArlXF0L9HJEi7fb
irZpbNbeTOT8RwWloBd5IhsMzXk3m4wtPAo5diEVw4dGDBNTki94iKcvCjQzzxBtmvDf9hD5nET4
Js8Mzi7I5NSh+exlwMkvKCCwyVWRbMZGsqucNYtdImJ65g9/ntaq4gmYfZmnxxA2szP1Dg8lW/Ho
E+fWrVEnUyK4BbrwHKeqjWGDmcAxgptMuzsR/BMFHnOk2R5NRDgzyzRNCX1AaJdO37/drunQrutS
Bq0U3CDsnYQELadFR4kfrobtgCAdL2BNQvtMeW2y5H+4Uo7GZpHgyUZ1IRjbXYXIjj7Cwb+kye1c
IA3Vw9cBJl+sFiegSX9E4BlpdLGwX4qJkAhqif6DNVtsm+GO8EADUyoFbJsNGQ08yuvicDC3qhdW
V7nStNaJYguBkHnqQQcIQwC6MxYH2+z/mfYD272jFT+LzAPwoCo8iiSPbm5ZP0okbdXfIhN7MOZK
NQr8NC25FDdnEgW8syXebJI9Q5CAsgQB/rJ4zOgC0/Y4BHuApWoIiNXXdewbcJcrr8oVrdq4MAJY
DLxqtrxdA87G3oLKJLY0fQToR5Xa47CK8xfkfJMLEGmH3Ilu496s10KvjVAgxvtFX7ZCIwI56P+i
bQ/yCuKgqF4YbGIZubvmHYrNvOnn4rEUobifHKdHv7vKVTsbYSzfqzbhRw+tSKq57RAtO5zwDelg
WGRCj1fgMGOqHkNDnAsqk6xkUro6sGFNsykiFpZZd2qvPc+88dns/CYec7YbRtyDOsZTBa5vtD30
oJ+Nxz5EL4Twp6tGhhY7RKE2wUh/7nUx8+Uc4KSqxhdo0b1QefNPNWzy/qnT+BNPhxFL/PsGzlnf
L3Khj5kI8lQDdo8ceLPb4l1q6BxgHxv17Mc/LLBNai2pMUW5YSVc1FDTgr1fdDB9acmCVtz66i9G
D98aRy6CqvnmXmBUZSpNgr3zHI4yUvDfsJ9UdDhSwhi94UqIaEFiYw/SZWY05H80BhjNlbzTYOew
89vihX68GdbQqtYrq0mHLqbu5cefZ2hatW9Q/cRPpxCkgIpsWc9SryAqkj/slkCSqKivXowDl7ye
bwIB0CcgDF4VKvHu3/nRoMCTMIz8nSubCQZD+5doxyj0K0t21lQoO47BEXdzCOZSfOxP2V7QUiKn
yaRBci+zDS23LBTRih1wTTVVlY6Z2ZBB9qdppsRuczx8fQrj/+c6GJh9jq4gDMCiIvsMcxeoiNOD
LoH7gbBxv2y/XeAuMqNFhG1t2mNm9lU605C8B2N4SzySSPICUfjzQRAzDsMsiaJ5htrcrtjrfXqP
I6KDUd60Sn9sT/sO9cPSxoNphQQPte9iV02BF8k4mXItwQGe15bPMil5DA5W5qPH4N8RCom7kyzC
oxoRRbakTbZOl5L40UDd+RTZSUCXdQUzLroR9RrAUpDqWvQIImaoWAQXzjFZPqtlGK8Syz77YXPb
OxCaVYJQIrEX0VZfErcAHG2AVm5zBbgrpSNEhYqS3pWPnkXLoQ9U5xwpp75fzMmSH0kbW5acn/F4
b8lZpND5jFZTIv21/CwWKgr+ATNBqFtZNREdCswoUA9vZFNMTUxvZv9rSs0/iF2us9FV8G3g+WOK
H8zdM8Dwt5TzDodnEZo7BYXU0357g1kCC9KISf5RdvrpOO9h1FQB6y1KKFwzF446IsaIAvZgZIqI
0gMXO1doY06TgzrrLcn1+XQPvahd+RDRO/Zjfto7S6l408+eXDftKqAEQuAg18ZdmoVBBlr0qYTD
t6ZzewLc1n6VCB6d3ds9kix3KABxOF9wOCHQJjCeejk1DN9Em4SmqRO+ThPYs4Ist/6Kq9egrbAx
4JgzahJgTdJLWrCef4elYSl0qN/Ieiwc7ZCLEYYL8oVvaGOim/FBjD06VP5Al4PeytUf0u/yFng/
liPv3ihjiI+hOCBJkOnIKsb4JwqtX1QJZFW/dPV3hQJDS7POxwZwwyPUDHKFUD4ktkhENiLD2oft
T5E2/1SuZJt0iuFS8m7TKBE6gIPlbrqWTIe9WvmJ0h/2toJXKTHYUU9F/3jfzIiFhLKIYyHuVwqR
OUgmVxm/3eRsNbmI8XvNRu0wB88ZBZBaAaRS2pPnvMW3lKpWPM4OP5SbrjzlNWE6Qh9zAS3PZZ1j
e2EwCchYezDmm7aoMIkDQdHBG0GMWknwMDLy/iWjMXBujJtaYm5gtQt5LxJvbsjBQS/G3nHwwCBL
/uFenGfJq6n406XHF5iZiQ0F8FmbIA+mbisR+Z8K2Zgn07Dhx9+kk9b1xQd1GJnrwmlrwS+SDMVq
ObB9ekag8spMH/5ZT5sULRlKhBxlxYK8suk2KkWxf8We1ugR7J8U7wBOEFZ0f0XhBLfCBySqvAI2
PFtV2vpRYwP13+rQEJiBq+JDJVceFsiLMn9606+GPleDJvOiN6BsnhRnXRakppErynCW8Zfbc7pv
6KqUNjzL2ZsCUkdJz6HHEEsLb0GfkKQxbt5YSXvnT6gOkTp+f3uEZQx3O4CrrqQUaEeizn7h5j0i
QReS2G5Xum212loHGLlQjPGoLBT8uO+qe2NEtYKmNAR6KfbYxKVJsbOfU9XPhQVujlB3Ev6uuuHq
Lbj26A8ICxRhv3b+LDAvFOIc2c9mXSK4b5oKW7gfrd5VHhxuSpxXsQjWChmJigReiA5TTaQODDCP
rnLfFUXLFZtXm1zmOhdLEawIZau2FmSB7saOJ5Vbj5tsu5LIVWhx1PQ/qBtI5xttIWC4S6DVFw18
+oo82b2fToYTct5p0l7qG3qxPrp1VJZP9WLtG97m7KWFe/UqrAfVqD8bjdOSn49dFdMIkI5JSi/H
lGFmDytqnQhBip5qEnEQN1/5t91EvXJC+cVQzUprubYqEHTLarxR8hqqXY/PccOwAXTvPjIMdACg
6M50wEelQ1uhb+ljqPME1DLfdat5tOT6vSGPzMlXSicsMgxx5+vJlAXK2uZ0/DTBC47GuSoLuair
Z7gsRRf32IonaZBkLxVTy+Uhw6x52P8UBCrKZVTQJwba426RYxZDi8YqA1D/Jh9i/Up/MDEBjrI+
qv0SgFOnU80KaaygC+lYJRVtPT9UkGVo082GKBuFRVtp34zUoMxeGZS54ozb3VsmkpvdId3hvFtf
S3yLpuoqRTW5uj4O1nVn62VxxTzwbhyrpSf0rrshMnYgPfdl4h4eObikmb7DwL4Juv5IVZPjx2Lu
f04UaqNh/mVNNFaFuJaSnM4ddrvdmNX3614+191zLZO/AwcgeU4w+JO3AD9xbpQcaiEh72THT11S
h0M0bINc+zb9bH/tm05CJlw5v8S05IEPI9cZRvTIFoHshEubRzh1NIjp4Pxobka6EZRvasG3OcVz
47O/lK27biKqObn1O3r8thexmMduc/COItJoBA0x7+AHS/HoLHIDQ5dq0Rw0JFp3GfdTU+L8ki1C
qStLz75R25QpIkPvicca6KkIe6y9J4tWcyTBZfJ+eEjqYpW8CBeH6tmJ2D+cCWH44IROJvdufxD4
+v4ZFqj9KcPuwBSJC6zLXToV7gVMyLNZ7alXtpKkTgyPKWS0PcVoeGjoznmOcE2en6iJYrXL+ePn
XUJDZEZMfuXLN9TE22Wa3Y2Ig+ryP3mTM+jBV4pdi126CLPGUnES6D2SvunBM6V/beLST07czRDf
lkDI3qBJUdjBmMdMIQ5BFWXQriylgaIyWL7/WBxADXU5ITa01zwpnUKxK5fz3gXbMXqctAdpEWW/
YaYh61T4hQIYUR/+c+FoRwF17doMuLRbWFYzM5S1Cdyyse0++GT7v8aOjPKlsIz3gtBie7EQQNM/
K9oDUrUMBKoqZEX9GpYTEsPVr4MFAFH7HRUMCfhRiKH+mIBLa9zRlCPPGu7+Aooprn8gWedyzdWr
Umw6a1ZZI6mnptY4/zCaXNub8BtQTnsmMnys0baMkAd7KWZH/y0eXlR0ZZNfmJqI1UHZrL8/UQJq
gu2CAI1iWfJxq6R0ewXyQfPiEuHTIJRQwNCG4TQI+Vw1pd7gmR2H2bHOLVe2EEzO3bYxuL/Dq6oJ
HQoUVKv0foYPL0QUrOAnZbgRD2rmQVZ9/lOPNW+k9X4P4K23dNJ2xkwSWQw0lGqjTaXxrEk05NyA
b5RaGkkR+MUr6gcjXTPSrv3ndpsJa2M8vBdnOL6/J7+59XnzgVS5IRYmrgbaxrm4na2DUP7/tkCu
ellm5sK3ThnMnHQZSh87PJOFmU9owtiqOT4wv8mbucsxSQMQ9PxD9l1imlUWDVLUbNyUl1TcBGB/
rDDu02ScKaSyi456rb4jXYXfTRscX20wLZh1zbsJX5KchR4iRT1AMbe9JQCL5OGtludspC7Hr67X
WfcTA8Mhi3Vn1F5Q0GTBSWzJg9W1zox+tZJX4zkqnupKqlWItE+KRrietZkSikmBHpIYttZobvkw
QQvHjcbTtw0hIotixcyjAxDg2mCpeMkQzN8i0OA9YFKVSreiZmKf6ECKbATVIkEVirtzUBh3xs93
aSUx+Vnpop2HV4dj/9oy7j3WzfX+KkKpUSlmoH1HsW4bUQ9qujEVR9n6sSp7lJJFF1k/bravDMun
rsHghtY0UrKgLoaPhH+RvyOAQA0T/THOtQ1h/QIoeyPrDK9PZUPqCHxWcwivSgez+w0Y/j6u25He
c9CvQBU+JWNYcrD3JeTQxIuQ/Qyt0gmVRpNpixcH18lFCmhBjXFdlhuft6uMaK4lATjhyaZiccgQ
uIdekB8veUr6VqsM+d/1wdxtP4+g5CuZyRZ/HsF8tkZeHY4H19VktXk5B5rsrQxa2P3J2t0982yb
pk9Dx+eK3IchLu1CXgrpwjI3MM6ZQj+IGfdrBqIvB+Uma+6hDEdvs2BIqiaW+pxK9H7UCz3UB1iK
z14iXpKcoyYoQ9rS8jeG3pZVL8VfErDiq4LhfHRR6k6QyEJRbUxOZpfv5wSrzxZfXsrI8PAiCNIr
XoQzECCCTCGuYdJ5BesuMLYaD2i9LfNQS6oQAa2n/Ndj7XfHDDUSqG/ubpnkczIWXhQtAuE2AXiF
HYpfCGW57fLRVzBnAQLGqo6m4aCXiU/HFq1IsY0wqwgdP0FaTtCRxNCgw3XejuBYt8v8J7eNM7f5
07WuHoicScuULs9L3BDznbunaeE3lLd3fV5rC6a2NTq0+tX3kogs6SklmCMBDSji32Tj71yeSHks
5jlnWggQWSDvFoO3KO6mDXhx1xgyucYg/1IqooB4o/CTaIIOazS1AhNr3io9hzjXq9ypNa1m1lrk
ognn/S4tTpq70IOITauzjVZQQ0UjxNXWsJkskNLR+NEFH11UmJs/UxvvXh6df2VAAyAR75JHkefE
A7qAFvWL+CGHOmXUukJOPITm2508hpkcg1pcHed8htLwzSn5SQ/5z70z9GVbxnqrGxoK9FOCz8e5
ijSjluskPqkJNV7hkGLvXqpYv7gz0llIeMjCFnv2fn8gEd+m1N4Kjk4+4tKzQtsOiY2KQBckNk37
wPHnC4bWT0zWaRS63UcxFB/1h4Bc6i+qjERR+j38H5wZSaZaCPc+QiPqHuh7fpjkeKa0Jva3DiO5
x6/It5bjNLZntSQG2j7g3uGqLeOOSvYJ3b7T1fa9rOFWHwfTPo1bJj4hCAcqvDzkuL+WETbvpqr3
R/A0YLYmz0uaAtRClGcfrYpi22f0JB5d+yyc5HuegNwuOa2Tisp5PA3doBxOoxeCpqqaZY98zdD8
m5x7zSSX60UzZ1JKDfMMI/0GuA6C665mGAdMl6Eggv/t6zs0bPpuSBbt4RfA7JmN3b95iafTb68X
uny89ckqDnjwDnNyU+95/Q21XooaMdHe+bHE/XpGgAqCzwzVZwlxRHIchS2kLCe1aYxkxr0a5p4v
/cFYHcB99iU3vkjXZcaSAfUUErn9WeFCw3vMW81qjygrriUHkEyBuhj04fWjXstOqkyatH7EMdoF
3oVaYEXczqDUT5NJBuloDaJ8jPPVm4rRhvo6czXbNXyM/jqz7VhemhuN1jVBNqFnQxb+Q2bBdOOI
nwCC2d6k4QPbFs9lAx5HmufCeLxBzGnHL70+5r2JVC3M3kf7GF7brLK6AKamRVxh7bZPhp5kbMpk
nbR6MZ0J2Hhz7j+GM7k2W7d/Am+tqVubTsiZ9Jh0gViHr5w/5GM6rRAwIU+ofAXDHovATp/SiI8D
jksLD3tkYpvAdUbsoYSmubsP2Okr9VZHGonpo/fH/hb2uy077gKRFz4ZrIA9LFJJeTebpJGN7G+K
JugWIDZIR7qct+IYl5gk2V+DSnkGipPjS5/MbumvHvu9qb2vBZ46SfKQgHThFQWKpYWho1GP/hZt
CdfJxOrCv/3ZBqpN4zkpF/n6U3sxiRXyZUQO5LUAEfEKsRyRkDYEeCAr3W1CmvWFbI5cRQSrv18r
VznzTBDm+pClgpSVwkyJCkBGNR7tOKBmPgQbq4tKY+Btf1JVrjvhAc3v4jhRKqlIfIeHk4GGalBO
sSGnAs12Gg+7jtXfzwJ+T7macY3ONz7+OJ3C+JrK60KgGU42G10IzEKo4ytJQCFUEI0DOZ2yv4f3
aF1Cbe5SV4IW1x3akvtFm9ei1jyldHUz+3aV6/LDuhB3C+wvSz6zOwRXWUkicgTp1OXiefUVKu0L
roobQLragXTf/+DrQez7fPPX03cX7LhIPtz/66rS5SE7ko869KydHOocXnQkyA1M4a2OsC2H12Ml
cF+MxQHtE9VrF/loXjXmhqcd2K0lVDUhGK5dnQXvBuoztwzRx+3y0PlU2cpi5Lrrp9Z87mKzPIB5
eHdVpjmD/SyRj79uJrNbN8126su24mwR14FFhtzqk/HwJ8MaRPtUABeyHcB0GVM09lRxN3gltWBA
YaUMv96Xz3pcYTOMqPxacglHPxvbZMT6NIMDc1D9MmIpEt+y1bB3yWynnEAxdvLrl36cJyFQNQX6
FeOHfthwCmbZe4K16XwJY2VGJcnwltuxVuJNpCri72fOfQgM5AaO6PsNlCXi4rDtcxs7X1YNX4Km
b3YTHOop2SDSqCu5Z8fcu+E0p4ktXNwjp91F0vdK3HyTy1kUrAVxcXKNyVAdxqT1sLWNhe4L7AIn
e68R5UahABQmIpPo4fYSxIj4vdnsCJIaUCbcvFYnJUtKS3oqHo0d4TxOdjh/VGkDLfrG31nkjn3Y
KsHUSSiEMfwz6tWwnTk2EYnJtOKn2X0kqvg00NgLsw5lWLWNs75n1mUk9f/SdBblM+XAGt+vOQCq
qoF6VGgwqrK7CTpaElydKNjM+LCps2zMsIocCdszx7eSFpWU18ksfla5VKkQUwG7o3ed9/kIYs4h
Um3yjAElg6LsEyW6APP/mWxR+PbR94N3bqSA/CLLCMdc4/2dOY+efXbBAZ+mJ8Z2LwPJS+wxc4Zp
ohJrSQhmDLelK9GQ21RXzVt2ZhlMHDap2XwB5SsHhZPKFJa22Wu2xQHueOSm/4nFlWsGqfMWxGmu
RXkanzFSP6emiSE1y10hVDeQasEI0UEL/jQa+TlDOo4zHCH//YSNsh3+R8JUFgFu7LJbzumN5siE
mp/h+ixzi1VY9VJ/DHoS0iY2nWMXEnWjlk0tq87LP64X+kNWULXQOny3pdP7bDGVY4pRsU8uc9kZ
lmC7lO1ynGREBgzPIkFZ66EtxndXXx2NLx5UA9TTnYH6fImAVnOUq8bfpkQ4C6rby9zYNP1scfJV
XMzNklxHrnxGj70zcn/hBhjdOL2CR4IKJBSIVaATbkwdTROmCZUFwPbQ47kV3H8b4RHQjYwrjA3T
f0aNP+sT3QwYW4NDtFNl6r0l9UyVRhdcvXSXSOYdIGOJiy4HJRqQquyxk3oit8t/MULaKqq5/PBV
Zed+h89hJ3c/fqVaFTdxRyUAG2m5ZIFh0P23slgjCq75VKXgdU3xIQwHGyZVk/BBjzC5hSTZCvX9
rpUjz/v0NUhWMOU35hO9cvhJ0joXZAGdk6AGWoyJAs2Rjff58MAymo5uzmFzYCAj85D5VRu0/fJg
YA2zwRkaBNr0dQvDuYvhEeTYNWX5Dl0sHyeQ06W+3gWlyaAq4NSMRxwrDNbAM9Ic+D/cgmU9e1hG
c2dPIKM+UceWNlRY7oqxLxQIMALmBZDcSlx6CvrulFwoxFvzsqX7veS2XMQSPT259TVsAI6AcOY4
FOhiO/N10Qd6ihPliZxfNTZChE06hwzV2algF/9z2n1wE9VshjNgBc3XopTdjFrsvzO+qBGH6A6d
gNW8m9lZyde+rCNAVCe+7Dxlf064hPgaF6iV3Ba7d9uf2up5ipFPd8dfw/XrM250lRj7+tE47awy
mHLgrJO+z19QdYXpgpIL3XxWaW8y7LBn52a/wS47iLTBeLnnNRpytbbgts4GNAROjpskozi2MH4P
jFVQAUkQtToSP3UwwuTyDIbX47QmEfQNZNpBxLqqIKvuOXk4zwUXelNouBUUY1bXaYtwNiXtxc/3
Ys6He0gGaTUTVi+41kt4Tv8woFKojW2WQcEH0g9atcDdem//rEG1iMSw0QB97sMOow2PUYjgtgb8
Q3ADb33+mWZjGs3ndRRfezaVhKz6wPsm+NL8FBuEAAQFhCqDUYJs7kjvUqWDR6iUjnGsyzjLj6tn
sduhkEcMq5qCa4QOQhptVI7D5zwZpT+AUr8n0bFaGTWAo+83DAfSiUru99a0WZSevc+F6ZFF/KN8
fvOQ6RlhbIbwPtjBqpiR53UJDCbwlACRG7uF+YLxKWm1JZP6QSFjv5Tpo/BOmiERxHSkBCbDHVYx
wh17BUKp8a986N6O0zUQpRmdEU75RLW+A2+deUEB27OTiGzW6g9POJdkdpWyq7bk4SCHyL1x+GON
cnBwFskBZGbRo0PnqAAawnfsINFFAgG2+1jT8xK82xNAQ2TclmU7nyHzdOqltkiOJOtoK8nI6t3p
jYfA3qQYqjYG6PTIRSu5jp/e+DFRlSAxa/Y8SOzgNrXk6Cby0EuRu8nafOxg005jWM5olrxUO3wk
flQLyO5VZ7Kjy6fSYRPbzjyao+bIEkrXxy5YUV7h3I46xuE+iACiZi+/tNOprwTcoA7QSVN/mc4/
liTa/Kf9LdkP/5BaI5Pqhen52Y5uYkem1Ap8y7V8HDZYnX7TYPVnxAjJCKAQdT5r3n9hEEIbCsWu
BFYYs25G0T4eMZsq47BQ4eTaEQLgBZ/u9X0rrI9yJ1JtdhEZRGZm3WdsyNClgw9Uh4CPKwQKuh8G
U4pfweX2hpmYQ0rbTKNFijvAOcTu8uVQI/mOpKrqJKePZuGqiJ2wWNjrkcCJobSD301Na/8D4BBi
4jX9dH2SM8POs1dfKymoEqkW9IuxCQI+FOOFslmYV6aZLmfmQweeWkscgrg2UWWDA+psUUQRDXJA
bfQ0/IyojEtd1kB426w516an5AOuUjils+NG0jODXcC/swuf64itoO9UnT4f8p1qHV7jtPtnVM6f
dyKeWpGu/KNAU7cPJPIG38yfBLMJpoO0ygfr3zkMR/wiggnqXqrHCKnXemJyZbtx7A7FfKbjHHyO
i1psuGXSLPoeQWCewN382gdxHup6R90aX3spHA0KH+hf/fmBqrRhLswVyfK5wli8UTl7cPSg5tzq
3kQfaMRTyCcWp5ZwuhEgrjVIoEHxI5xpzWJ80If2w5VaWVAIa1Xv3T89whjtaNek1zMTekpbqcA9
cc/30hmORRSxlr1cOUafpZ0vUy5TNfMrK+Qd0Xgc81iZkj41pnZEzXJdV39eSxE8dT7X+YB0ZGMC
I/vCdPDbYM/ugqsdfBOeBZUXh2rCeHj6x+7YeZ8lHYlIwjArgTy3LkDmt5sAbe0m/kShsPfcM9oG
CX/Iwq3nRQsN+qnjXSxYYZ0p2XKoVToSq0yprrpuoZnqsZZtHbar5xLi/UTkHmITf1s8eOkGcXfR
GkZmvDN7CDUHjAW49fl/vmMPu2hskYABDGD5XOZprS1oeWWnkkHvCqx9Tbgg0cn6TQgf3izF5b9G
anEBkcEN1UPWoJD26G4fkUVPqooszVUm+uU+nev5zNb9YyQJ0IIfyyp3NDvdgnEx7gU1dihSXGa6
lAIM7buZLKVhVkNfXC/pJuZj8YihT2bN23QKp3Msgaz+guwC+USNgycaO2LFWEw+3OW50LkOHfhX
SI3DF3OPhEt8yAFJtUHhcqmHEjzcMDtCNLvZ/35bBoJeox+/O4FxSuOJYFtKLavwJrMqgKV2gyrz
VqMtYIqMnI+HXAJV/VhwnpVbmKd/0VMQl/+EthShOufh+3LeSn0Sesu82dW3Ose2Puo49PxgoEx8
FpHP4wVwYo+gGVXvMLGds9h68N5byDS/hjgksCBzjw6MCrP2a6lIy7P0ObUYp4NIYnJcIPPupG0e
CBlXRZgbMpNEp5bhrylm3dSDZdTU5k+ZAvHWilqKEFtw7AoVA25tsl2rjftlmF4Cakw9Eg9u3PRX
8GAMgfYK0m5vKOIAN9ptXK0r4taEgfuH41ozlt3c6djCqpS9ZqwpWSv1SoX3S+/O7S1FXOxMKZGt
yDyOLO7mWsdItKYl03abHQYCUujyI5BrR4ecP5bmPTH3WNwEojsxx3c9uoXHLDHWHQYZwGQAYEEw
FiyVGbClFuU0VW9jQQEHrLcZx1nx/z5FBx19Jjbk5hBm1H/WGbXENOHgmHuUjIUPxbhVAj8PhE/s
E61VRtoGrO1Yzh1ZncZj8OpazdzKh1WDsie1/JPbgvt19OBKtb2xXy50ZeFI9CDVhbb9g4exwWDi
T8zuLBHatXCPFprx6xvSGfNqC1q7sSBn/bUicl7lpF7KuKAoUa2f12GL9hOcN7f5Tr74ISLKRO6w
h45i4noDuvlpS6J4MoPNYZ6Tk4f9XAcYVsvgd1hFXV6XYWNK4+Q5YZS0NaYqiGnx88UZPt/QYKFb
SlcrTGmzMPPdspDvlyk3J/WWnivqMLaBlUsVIUp/lzg/Y5XvPDMI3eBl7Axf+j/1e39JeSIpCace
YcqnYUojVLfcxdZ5jMPCj6sPDvBVkUSUPRwB+bjLfQsNm/pyIhVKcOn1D8RAenEawRiQaDyoNQD0
p7W59s0Kc/4loXEBtUArW4KSYi0IqFFd1t5HNcYzOWEU2wh+bqMILbMa0NjaZnvKrsjBpvYuumRb
AkpY0YgNS6EG0YUaGa4MdK4g7r7i/dXBMlp/k6wGB12C0YaM2trrGWDx3U8T3oJRj62I9nV7/ZQC
GHWmYEu4KQbgipYr1w1eJAn92HPD+GBJz7s2Js2t7MW9xpwB175J8qONCDVIK++NFxrlbXA9MyLt
iEhaLObDdmx4XrQ2ruamkHTjlRlnwzrrKSubrPxQngzduBMYi6h8vijahN7X+yU7HKXCJTWi8P+K
wokkWeDKN4wTfyaHOVv0vxj00YIodPR1y+DTV+MHExtqnv2M3luXj/ME9wlCYite4dan5yv/pfFT
NJ8nkYUDC2FZWYNJH0OqvyTuAzgRj1AEk3e/tbftKyftV8aPcNIzxneOxs8VEC5pRuIkyRLgiSpJ
hy/Xdg4l+d16zCgfDdBSDDdKkPoHA7tPp3eyuocD72OeJjVeS5PbGc5BI5Q3KiMOfcy2YYMSz+Al
cz3OJqVl9Wufr+RRBelF87/d3Zh2x0k7f6lZkryvtPqGJzm2oB+/e10GX+NJRQZA88wk/gT0+W1G
1WXVIyxti871U4QYwI4z16n9eXmxO/QDrZ6nYMBm/Po23Ypee6ybooXT86c/rTY4vZDdlpR8u8YV
3OeSPevRjzw0U2GgaslLO8JProl3XPjph2vdvg05nBbIYnplptTktoPf+UsqThJ98ibimsOnMoij
hc+YdFr2PmFIXqmVEtJkUltEc1DcYVJDYfn+678Dfno555/IgF5vQfMM4cyO038fDFTQOg6G3xK4
PZHgnCdJlwq5cmXZxmSHpIeWyJdV+gu3P6Cyg9xVymaHNkZLqbd0LsJiHZ4TizadBgU31wvrF5mj
lV0WIvXWCkd4TknlFi2civrI5cTQMIe3YmRaev2GbscSR2ZEjgaGmsWgy9e3E9diODIOX4q8Ql2c
1fNIIlJxRWGKts33/zXwNSS2mcWwTDW0UZ+9XmZLMNupLXNHtiYPVwnklJqpvYZidig1Z4sEk+3Q
JwFfxvlpWtkccT/Kbn+fAamzeYITuPdsYmg3EHXu6M9Lfmer5p4/k9AjwVetWKap1Sx7vkg0LV4i
KD+Hs0c9yPpoOabZmkrJ/c4GyXnZthQAEKZhigLVgkg3EL/xQ8BMZvUykJLJOLk/INytpsSyIq7P
oieW8zZRCsOjF6gY0DRQ16cKuxNZ6tkFkzAnyTZrnGSI4Wp1uP5Y1S2pcoHGZ1++KCK7tEd9klfa
fXzmX1Hh2i3G/TNsdtDErDT8qASLrNIfi4Fo8lc1Cb/QbgkS6Rj0czTLbhMfSFJnkhCqJak0Wn9a
hxGog4R2ve9i2E43FEKtWZjRK+QVktH71S4XmzZZ/Y12mE54mBoEgHxCWbjv91vzR/5wegyNjdzf
IurS2OmsUSgI0ENZDe9RSiEn08J+SMdxwKMNEOBvoLzgvxoqWFvch1Zmm8gpUN02oH7K+AxfXVql
uMpXqufUIZzU79eCxF+KXiAC1Fj9swTk6YLF/B+T7jmXgYJvvkUBgQ6IUGSQNQk35FCI1XISQUlP
wpV0+R5esKH0jJBrrZG+X8bg76hDZiLtyjbJ5mx3yZZR4PQzSV8VuPTyt6Pc8LeQw6i2z0CGA98N
yu7kJ5cjC1dERZWT60CL6wHvCxqbxb6hBkdJMaE13odxMFbz8aX3iYepMGg5BziKswBNMjfN9kyN
fEHUTtjLcmq8FDjcNvy0AnW8dTRtkTg7vNOwmdQq+hdchXzX++WbGLylb+IaNrE8gX9XOVjNUZem
GzcQpdSzJgUT0VQ7rLqU2MZzy0MGxuPdyg0HXfa8leitf58sob+DN1RrYTYHOAWMDdp3yiylMuUL
F22pX9MMtp2aFx6CcYl68gL2Mt6CfTPVDs9gNm3T+annvcKgq6fUinhtqLdbSib94tgvBIGBT3AI
a9feynlmz3lA8W0HB6CABdxCzIAE1oVgQEdBeiQDPzm8u6hfjNEDXHhV8DwwIGCS2xUYGKndF3Kq
ID4aWtxMTunYvzXwtuE7eQ7W0tRF2oB9ox0zzMKOmAO54NBiYkW5EiKOhndMlY7oR0Rjt8pceQtg
yXku6yh6wA11GrdVFteK3xFyUyiJdDvmigGw4ZjjhT38MeQmePoczfpwIcILrsbLJtLoyAIh/APt
qva6KwsyslUzv5Ud8LDoqrDtj5iR++NjoD9/z9uTp7W4bGlDjGinz3VPFtKSzJR34iIWQyPGzAOA
bp3dqzWxcmdpXP0LRt5VyC38XjfahmONNCxmDZVnAom9alD9j5tTG62xCOjgayraJWhYXLYrN2uF
q1Bdt0vh47IsjBmGME3pFhS3gXMovPXy6RlaCssSCPkt9FPAoHVN8f0H1ixJ31+XKjvwixFzMTq4
WrHIFtFtA5J7mjGR7fCyiH+/R2Nv0FlNAlYyUKdPfmeurFbfkGzxFEoC5CUkCowpuboSanvSx2Te
DnD8w/orfT45Ivjq1GIaJXOhSHve9clhyIVumKgKx07ajndrNpVi5HpP+ratx+LxCguThXf/5Nz9
E9FZYj+LdhJpig61oFLk+xOGydniTfbhCke9SQlbyMHAfeNYBFZOhQZq72ELHghlU2ex6XpHnAi8
ChuwFOlcIViIhjtRQvyaGufKpaNsQBOB301LmBubXuCcxt936Mg4jRDs4qrQHvpRcQsTXyXq/JDb
lGaMUBtI13U/WR73XOhJ3+YAPkkLMC7K67JFvQa5GmGfcD2kXEQ0Z7+/WvQtL8uAYxonVIcaEXTR
KBkGXC0vZMahie+f/V2yQ5TuxfwY50p7yM016G3oIISDmruLvyDu+cSvyCaw1ZwzJKb6+RRs7+fO
bBtf+j3e6GdaTAHEvhmj1wNnP8je0F8228CvE2ZJMcKLPJavA9JROAXm0nMFgQwULNmf6QTc+EL4
gBdT6ycgN7+kndhh6DGTeuy7CE8hE30vnFmVMHbegFAfM2ShowCjwenEzLOgBirdShUKCfwpCkwJ
gMv5XC4/qLzLtCGdbc69XFRd3gOZNlVJUOteOgDlo5WFq4etX94E0IzS4zdWgU2x3rzfXo3EtvTi
e8yw49d3z+etUAEVdGtLgBr6FRX5bAOYCBGlF6qdg/8Y19kyFHkv0nAHhm0E1gGWL7Tjb97g4Rsh
y/l6aU73QiocHjN4Eea/PXXhQxi+w/+SZ4DaJEZ61V1c1k719hAgjLE7t8LT+tkVWxGp05khBdqB
tKDeOhTQswzhYFsFfVw/il1nuackYY0meScixtGMHG2ny6ttq/2CzHYInE5u9Dein4tfr6h5mrvZ
eG49q7Fbtcc5iQeVFJZNx8fbeu4cWvdnDkzAqZTIdQGLOhaWVLmPlGbzY4tzMDYndoFhuVYfXVG3
3WfM9DyMkWxxTaSb3yMrwmuOcllB0vv4tlK61Esvj0mKTV6s+g4UvxX9xwIe3r+8kNAWyYEGApX/
T3lx56POmHeakIbTre7F0NrOYSI5dfv9WfkjwydzHTNNMrzb+8TrWfXN3NVPxeXNby042HWD1PGO
1MhkAS644zwhzYZ8KihXDqiiUDjLHsoF3Dnj6leSiekNY22YBiz5dPN0qyAtcPtxGORU2hewIxEi
OLGZx9Qhq1n7aF6qxBrYiuBmBfvv05FkOTsjbcjYmZTV3L1Oil4v5rXZEiLbpc9r6LPRLqzIclUT
gt7uk/XYMkknMRbDBTVUQdWJER79EhXwc2dnRs9J2nXiPG2js/xaqYP9kD1Nb8+WeurOq7Ry11t4
9M2AXOUskhRvlpP+Rla9fo1Zkr6Ldt5z8LH55yFObfSd/evcoDXXbm5CxiWT4IhTi7535aY/v7a5
djWyUzBkiWfJpcGzPJVbyw6geG4/zElVnsB90seqcldJGBKfSXH5IQurAq0+f/YqSmDnpedHpJiP
fT3CRnB2aTlGH8z9yvT/1CkLZiJt23B05LDzMYvmPwXH5/MsK/lSNajUKk3t4qy3T0yFIROLEphq
Igja4qDVVViVkMZMRKgYa9Lt8H40exkBR4KuFt6lHmy5WAM/CYfCK/bsCNxW4vAuViEjzVIdYuw1
DZGvpLfRT4pdyMv03K6EOcMIrqo3fzHgSiZztWAT8nAktgJWiFgXBbzXy8r5yNXySi8GVyjtgZLJ
18xbnGXWeU0kfyIBzQRaSf04w/0n1kB/ziXIToN1XeGD75l+UJFQ/Zjx+y6TtKRV0NO9h4ZtF4Zk
TVt0XjU6N5rzJHVQBck3Syz+D/B7DCT4WH/GZPQl+2BFTcWoQ6hcFBXhoms6pMnHb0BQ65rrxcWd
r0AjQeXnb8osaR2tP0fKydAyiWhkG/gGZKwx4uC42SbXtlYy6rvDEJpmTAP3HDG13D63SDjaakTR
llQzOg86pvNrzUYn3jf+DlQDUocNhA6FhvMTSlpTHbajiXY7IwEoInBFVypstYOLarpKc6Bmy3pf
iNP4cb3rjPAuzW+cWbypGRf5lIW5g/MJSQOuSmeFA2EW9wZvWZovxFy9N7WPHM68AqV29WZmz+lN
QLxQiLYizLo7HIQRaVWPnGDgzGhDe5Go+n0p8BSJmWLeubLdPldeWNG1Kw6uSfQQ8tGtkayugDyI
Z1lD6qQRrYdNYDBWK/q9njyEbpiQdkmQCtt1QkZIsBLuFbeQWqgn0zjohS+DufHgxPblzHxA6WXR
B1zoLXb09L92NIuypsbeHjCjfkcwt1A1lTjGgtowin1xLqYEa2ITK2SD7QeX7U8tRiEFi2y9nqOq
ik5u9GfkB6SXGJSHs7Vk3Puqsjj1XlNH2iXunwFKHPwGFa5r94B9a0efQmopVOtsq8mN6X0tPNRS
yHUAhIT+cK5WSr3Ja87i5cB7XC4FrQj3GQKWknc3JOb0NWvxWerWaSPe176rxz5+E8DBme8ViW7l
4dBURKFFFgHtlu5tg9NKGGfstRglhFzfh4y1Jyof7uVGZj0kwhpZ9dSn5cvw8WfH1H02+Mn3FtOf
OExDDqjyzHMn301nPEvKukjE6y0d6WEzmUDfpTsaS+JelAe0wgXtYf41nN1pTKfpXUY+zrqoLYwc
zciJydJVEChImKyJ2V/2rCzGtJz2mdjXffIWCbNQVyFDzd8aJHYClKUmaXIaipUqJc6x/WV5B06r
4aCHgyPl4aFWNh0QJLKTh+9FoievxVbQO1gSC0crEsZTDHFIxO89RRPstbq5pY87q/g8Cd5ZH39E
+9qXcrxE9ty57X5mREMp6m7XEcmSzDTkZimNa5w4sNqa6hn3uA4d6FgbO0BkCwLrCMhQHnpuZav/
mpQzdX6uYynBlGCJtDcon5WIGxyr3xVpWtka+lxwNV6nLd00TvuxOcVROVfS+HkVItopj57PT0kq
ia5t0vEXEaMf/l+x5tJa5hpcNBoza7W4/6HVkfonWshD8Kkxt/wI4lFyft3IRm3mtRUbck/XS7LW
m6r6JxbeDoaGtf2Na9oXEGclm0CI4NGkYUPWfd594X6KhWQU+i6Aiod8CmIteYHl/+KxqN/L4Ezd
wiLBHI8oCyF8YfAmy9nrC1uj7Y8Tdu1eox/xf3t3yMuvh4pULWqYFlaHV0VtEsYQ/muW0TRCpgJ2
1lmKuk8JC9g+TO2kJEFk02pTBIumedGhIXR64EozVW9GjwcTmTaZQE3ieG4fH7+riUXcLhxRpmjv
RRBwYiuCPGlZIqwf+so44qskSpR49ta1qMqGr/PA5IcnDlxPSNoPuw4k1kxUdHFbLNVtMNQ4ppPf
zfjPshw49S3kJXpHdIXMh3LINCDza5YxAS8wmVtlxz6FqkoErv/rndPwPTFqhTBRjOcdDW2WYsvY
RFq1qKgoM+acHnKV/VLd+5AbAOCTvuufu0+fEpt5cjnWeBeaxyOKf7RHdDwESDwk5yQgexJtHbTx
uLeI3sK9CzIKvxd1fBGuTePuF8rGwRwz5kZt3Gyy23ZZkVqmvAY8ZQHZTNiyV0vxX+6n4LFCFTe6
iyLNBldZ6BgoVUu26RgZspTm/SXGh+o5YiRP43CMTv336fIBWqclk6g1SrIfSB9xyh8QsjW1MVpQ
a4N+Hv34ZNeuvNSPrG7u3N2FiCWz0TXG/PKLeozeEaJVGVdE68C+EukK67lttkUd1KwnikJCp1Vc
5An0cAHAV5Z8+bsqXBB1OlhYPd7EGZFUuIV800GO+c9DfFMFydUdhS8+m6TaX/jTEAMV/wig08iY
ifLb0W6VM0xGCdoisERq7YCgI6fd2ST/ocSE4TCoCElD44PuOiOsWEknjuAIlnvJZ/uze6gSEsbF
0ZFus7zON3pCIxRMoQ0GbKI/afzgdIhoQaJ5B8XpvyizlXJu+yrRPMy4bx/oyNITo41NFkcAOwnI
0gm7NNo1R4Kt25uYmX0bzU5n+BUKkS/BwRswAmTKT6AQvxnsWKt0oEElKlBnpHNTu7VpXPc/j1Yb
l26qa3qj00Fv0bAQPuIvvDI8eVY2g7tnNgviMvCb3gBCIbxBJrIlG0ztR/4EDtfRYxxsYueJaVhw
o7seq2gMfKIU4tEWNosoTaKNjx5zLZrs3LZOTnCElNogBgX/CH9E1Lm7JOdpU7EkzxDcMrQBsiuy
y4ZMkn0ZBM+nhONXkndvPILhVgRe4dKblk3kcIHm/+KQnE51i6K0B0E5j4aHMVoYGSlePUQyvt46
sNkHXkejrxsquOrd2err/mDVEj97rapAzC8wsXwKRRmvxc0JaPfer0I5d0qhRxnz+0VEhwfi1dOL
Whrt4QnZ6nwO5YS2PJtiERW6vLwn3D6Ai/CEy4B2JQ3xH8wT56dS+/W8lYWpCRBf34AKnW/2k5Tu
rrF2dFozQya5EJ7ItsHi24VrApPke1MitR5gwd6OnJ8pKyGBAYgZ5MhKewqSted9LYrv2f1ozJVI
CMmO2EccoX3+omAU14Pg6s5zREk+igAl6drSUT7jVLBLhWPbrSxsVv/EnWjvfrpaKdSJiwmW6Aay
FT7qMa0r9GhDfWu646HNoXylefRJDy3KjSCNRnAfoLMvhi+pUqv0t3CNHAFQSLAniXW8/8rpVQjz
NlrSrrZOasST89t6QfzaMAstqWmEMlBjlNneMoXUqR2kxgpTjy4FCLekxDCcFL5vn0p15bV+3Md2
W3nkt9IZTbpwwW9O0hh+caUGgcVpqwGEHfqQob8tX0KeG+VKnJYaQ7c54+bBzhV+RE4uZjOn943I
xIhRTnm69bQtPvQLn8LpN80VBE7Dsjc+8MVH6D5C3NGGhhBe1+H7hCw5mQF/f22LbGr0K2kn9mZ9
h29zLkGq09EITBMrNozhP7VtjKQqVHRqst6gxdCkQIy0vJU2jmkFp0mNUKWDNpyTf4ZV7rbPHqJ3
YeMpr0VCJKSlc1MThH7+vJLwuVktNzqQDmhcyuR+C1Ns3hjNCVHFZXi3EspFf+RptBP9kZaad5Yz
XOizA3WFaeH0feu0o2xwqJEOmyyAo3FsSmrh6cm6DhpzIDaEOT/dnASB8vj2omCLEtVuCb8CVvYs
OOK0lKc22JOFx/xYRea3YlASfEUuaYgKXO4NzQoV4G8PF/0s5iehJkuHWtK3ugtz3DutuyHg0YIg
if5xKMyEf8VYElM+npDRArN6Cn6miFsPPJDFKUxdT8FLH0TK56kU0fcg9WHymx5L6fNQrCBwNxhR
X5VqVMfcC8e4lD0KI7mxenUfYkCudonqwaKA8SpYljazNZbpSa/oKeuaxMKSsa+LtNwTx9tIpjui
evB+XAA87VCzDtCziB650JrBrAy8pC9yvHeb7GleDl++yxNCTCBkIHoppTfM77e6i6e9EGJY0KJp
ZyiJVfoRRDe32VzDi3AtvSTO02Rjs/rRMLEv5at/rikFz78Bm/w4oHk9sajoZaVvQnCwYPvGkfl6
8tHeKWHq/3ROuDjO4xn0+iYhHHbv+Fss9mAnyklzs9Z4+4R2MTedQb+mwyzkxQuJoa6jKn/84It8
Qjml1YB179wMBbMK7awCA07+xu0JwSi9GydKg8Qi93fpj07UyUDh7WdSKoIvIS9/yIOHqFzD985d
UQr3fa6+pQDVEWWvgNlggzQ4GmBV+dqBaAgeqOEN4hdiJRp2O1sp2YpVahJv4X8l/OdsuwnfnjjN
QJ/lGEZAGAzLArVeJBVWU/VwDj4H1GuWryoJzGEt8xyBnyLydziCq/31xCALQAjPNXvXwsssv+r0
ZQVlxdKQKiXiickkzVCLD87mCj0MysfjL+UobVFJcbTaM2kKsPmAsqyxdagnTPgbReQytIQwqA2h
9F+n5nimLBt7MG6B3mHjAvqUhs99BoGHKzz8LcMVEbnF7Nq8ws766iuA8f1xp4DV7UyrcClH+GSG
gObdWc/QjXj2CzZLEK9jem1mqS0fYSnZciiIsKKO6aseXeWwpiDnt9o1LzGkYwyuosh8eGHj6yZS
LLI0wb77lcTUZsn1YsndSC/+d3vCoKsJH6S8EpwtsFKrr6DM0mFQ7Y1oMar4u37HIS5OiW7d3tmW
Ql7nhnVSPTc1MzDc9XrS/30dY2NAl4RIQk5bW37EuY/ZCElJczla9SRaN6KF7Y6XKXJUN/NMzsGU
KF0s2EPVGi7zfVmF5E4xTxLBMiHjRu5oJOU6tOlYaDxNdNdRxVBNg+lhuPh1sgNCoCcWPt9ezyjt
+Zrho9/CHyDO0XKiWpGWzuOyxpJM9uBtWRbjQ0NxloVJDj/wx22zdqXUDoLKCSG2k0lr1zwXuDD8
WRwtap5asR7dADfBaB5ToFCPM1krpxs/BZ1kBm2gjlzczPlNXE0c+w4CvHWVem+TF6oRkv5vq0Gc
w1Iz1LaDO9fGwWsvsrz6jABZYXiNn15OBZC+uTqKfE0aMesmJDiaTqsvZ7SOMjaNM6r5Ncz7ulWp
CpmyfjLpsigi0W4ijVY3eH+zxRNs5ql01mWy9094i/xMJwSK9AEYnhrzdleOrd3K7zEu1u0xcuGK
08k2MAQROl9V03UMMH3A5hKDynFThp0yXTh26Rl9KA2YJQgrKK6ryYcQ9B8wZfq/CsP3MoF725Mi
dUs9/Mz1ecUfv+sguY0DfTRDZ4yaWgcokEcfNUmqnk+QlsoA06drX6OXCrYhKKS/budJhcwWJjW4
Fwz+th+aSrsOnHtDZcYXtsanzR/AybgmLWOAACt/ScjrRSIS/0tAcVDyzOH2Ow5ITmA+D6Z18SRm
HooXLFhmJa7C0U/BcK37jcG7ODPvEQHZL29gxsO1XUHEpjBOI/oXaVz1PHi3tWd9u68yFar34qPu
1BdNlcc7EukjWFmhzYBAdkvqmV+gDzDVdg+G2JK+RWS+V09HylZPpdoKPFPS928zVD7RplU9b+P7
alsc3G3NNdrOpPW07S6v/i6lxXj5Yqcsi199vw0s1c/9HLa1IMVLpbA8jTJxivcXzjZQO2GFAUj2
R/uWsvOqOOnrbsw5+sT4dMmAseJYej0pLzbx8rst6HqSGYJHDLz/MZyOfv+dHBcxTybE2yj8/E10
8uXdru/TLexnkqIpzdkYBmwz1dhZ57eTL0hp9jG/HebOCUSDVFwqvyFUfhf9+jnviwMVXsLOksSM
0ICOySQwecZEznWxvUpW6QvpNdAogh9mLQJwmQDvabz7bje9CBE3ZPKXCT8YQRz5QoNWFaFdx/LL
mZ2lYbNewAgmcIFu16NJu2capq6ya1Gvhh5KnE45CPSVX2oJrpA7nLX7mzL88KUfPDsAenE/J3Xj
m8n7HlJ8P9XyvNed0oyHfV4gLrWYimKw+YfQjHa276DxCyFE5aWxVMAalYk+1X3/OqbQlhwcR1z9
i6eSZ/FXazd1v4P+X3w5xtuHYxCDRrZpvtd843lY+ZK4ahIFJuMCW4F1oYgEsijQiLebj9tdeH/B
B+zyb8FwXKIDMJMTn0tthVY0hjpY4TXBmsx8RNeJguvMhbwX74N72eVdJGRAM2dba6/zE2Mx5OOh
DJYvComij322/mst/eXrRJVijVPoYZIA5/INecmmQqvrZUh1MZnhPDQztYEqW5DOQ13pcapIqU0q
rcfjFkI/prFrWb0kML9qit3aH4Tv1Ju8aWXCZZJfXe+zY4rsDug7Hb/z09W0Rs6W5tffPwmw61mZ
Q2Uk2oZ0lFx19gMY5M/VES15DXxwSoylHDLqEezJx/N0opS/F/We0xoM1o+Lkw/Dh/7HPuRW8u5P
gJGewpBqESgcXmJcfdFL1U6ijtLwWZk9v9a7ZhdMC/QNJD6g68kbo65g/Sf9uVYbKzEfD9IR6bkd
ZPYCbzVJIe76mPQTH7vsdgZ9nOOT56mPMCThw5ywcjK5/aRguSKatW+zO0LaLwoOUGfLmeSy/ke6
EwOQXB77u2QDtQnRoGAjTPEqK+uTuHbr/rrpOqrSFXaLhFvx2Ehk/q7+TEepU7KAPK/5r3RJi3EE
TbqFPtJYSYUgPb7lRgGpdYHTwwZuayPViLHSHQKCgZIEy5+Z/jj9UyUlVfFMAdVwKlrl3RV8e+6f
68DqqiUZtRWLSqpa6KM5eDthwDffE9JfMLAtv/SVn3hxzFnRFXvyCh6v6C4wSRd+4hR3on0jpZus
c14UyYgHcwI3ajgFJdlDMh1rwR0EgoN9uvNXrEuBqbV0g4FOFwh3DeZJmqaWHMBKsECa4so43bea
rfSsIEJ1dIHELKlUBWXftsSB8kJgpxipj7yJBNHWjXbLCdShRPBxZVmqULav1IIAfFScplLegmBt
yCae/ggjJVp+Fz9dgu3lA7sVxmwNNjcLl1jtLJP2T2tk0pE9yyp6Atls6bHad/S5JC6xFTBaXLpZ
yrDEWZZm+w0mD7W/YLydbKTA5a+J6LqOA1S7KswrE2nKziqiPLZ8TVvh9vBD0OWlh5JR+8WiASDS
9B3zcpWBJc6AmAVDqk81NxYZ+XYneO/oXuelgh9TsgJKGMCZ5/PhNv1UpPfIRGWXFklNOeWvq2jD
OVehhED/Mqostk9sNZQZaRizyk521doZ6FGwum7N31bALG5/UxQEmPSlhUoFwbUaTzYJLjU3D+78
r7H2sDT5dxTUrqn6I/3gWN5CZ0heyRjbNCs/8maXrmf/Zp4NEAOERG/kjVtv4a08qgpTqf8rH310
4A++uvGPsisw4ifxv+VFTWngnzON9wkw9GbvyhwUR6vKds1shf2otPHiN/JhUsSBgMk2YiYCc/Hw
BNdTgbl7ar/YNp3aGbYr7CV+T0/96F2+nFD/HOrPI4RBVbYrbBBzcw2wwyYgs8H3RIzGBcTNQEen
BUjghpAk2SnN1Qz1/f6crMQuzWtUD9AVlUKEL0sYa3+FFYHcTverYnMv0IoWImzO79cpw1Kps4gw
Kp6IIstrjUJHyEyAFWCj4w4PB235qhkKIMFFvgchHgfx8Vd0GUtr8uwLFu0kwz+GJZqoeOAT/2Bg
c7DkRltOVJOm/dhgbhBGRY73Gl30UuYHa9BkhT11R1ds2l6ylHr/UHno/hdhto33zJfeSgAYVQNn
1VtoeUpddc/QtBDl4XIl5H5fLHMNiANn1CGuQq+S3nEBWVVT29aKGNUN2afEDUDV565vpFQb3pfx
03woHdahfXDEwH5D4BWF9+6+1oO/RlEGNyjqECTQNq0P19bR0GvCNpArAQDcN0PAckwLAgW6QaSr
nWALRAhxnn8sgHJGkBthDXIuwjKiuIh6FiTLGU1uHeLucvCUx28DpsOZbXxpItW7zRiczHGSjFFR
qbmYX+oPE4coP1HbcjIViAOsYJiahWm4fDzKi1opA4zNhHj2As9gVBt56yWqyMpRzB6Hilm0B9rw
Eid1qvMIRBZyx/92n4pSdLLwjGf5FIKl8lESJFOhxxtxJOItyDrN0f5wgwpOtg2pskKfAzt1H9yo
F5JlZiyTb57nlOyCuyH5oqO/89pxunMPTFowvvs35PdKhdUQ+TGRScFFFXCe7iYPg9tNcx3aVj3/
y3DEhOrzZALgx/T7EuUBUrwrTMl2laXfWEMWs5FI6UNRrXlkyRB+NTB9ztcr3qjVbT52IYmUd2cT
6/K1CHaLLdp/u6yePlv7xAFtVxYVUXmlYBFWKuJXw6eziZjFoT3VS5PzWZR0OCjUMsRIM1QbWylh
8uR99MH4vFGwkTQv/NZn95qo4lenn2Pu2CwHngzcazkEJnifmxln1HRnF/b0bdbr1rvmGltDh0nv
0+cWVu+j+Eh9KZvCOLkW7bQbSQ2FWxrL4NFcyhqrURqaJIb60rX21bg9e+M1goZ1UiWzCsrnE96N
7iuYxJ3dFbJ9DYajWpr92vxvBub9SedBPeLDYpCjIsDn4cgkhaX7fneV9+6hHcI2jxSBbZJ/uUs+
nkqN6rC7B1tQLxIC0v5kxaWAXlshE/YJ6zXCoEuFd1DDbecvFLMJW80NoEdjknjimXa7ygu8rTVS
oHe/92m6I9aRkOapOvYYe0UU5jnGvBm2FdL5WWlbYC0hdfCE6UILcGvWqgmFROB/G4vXjdBoG8uU
Oqq4ZgOhafzohUXDvRPjbw7CVoNDtLK30anWu+Linp/ZPHHsG13eI1/9EmEbLGx7c37HnNVzFHZv
6K0eDfiOfPgQO6/RHn5Nc14XjFKLlNko6Y3ArISlp2kcejEByeWnZAlG0GaGgW6FsD/QSrXdVKpA
dryiDC9p7vc1jgfLMC7+N7DXFdzn8rkcjLtqybYx0Boe8Aqu/5uvI4hQmZw+RQHbrXxN9lrMiMrB
EsfRzDc7DJ23NUeRr32niYkuY07QCV+/HB1q8d0EEvbwBwcEdRZmooTs8JKAxIcQHEWDn1Cwk51s
uXOsGv55rrexCdpaD6t6d4OQ1gPu+3y9Qsto8UQE/vWOMbTfsi/PlUbb5ginRUsYRjeDIKyHp/gO
lvo+n8dZhFNL17j+NPmuhnenqAQLHElvivCWl0rqXQD7h4yQ6oh6oe20lsZoAQ/1weTwheHUf7OF
ISuygzuzuriUv9PBcAVRGbaRkwCJzS9JzaVK+QpdYMSMiaOIV3uCARkr98vqdcn+PrE4j1F27yAX
6LbvIfkDjSMv6wUbmZdx9fGkG3xdoIMXrs4041nnKPGTrFfezzhBSxP7rlbP3iV87dXGtwVYySM4
ixDx/g+oSdETXeWlAXLd2tbvyT6JduFYaJc6VlGAAHMYX3AxEpotBtL8R+JT0IbUQm9Nx0lT7r2o
9E+TIbbH17Dr4vgoOW9mWyrSbpgpfBAiCSLfbpC2GEPLOXLmRuvFS9pCHwnBK0aOKfmmUY6Kyw55
bI9GWQ/WXwt8P9nDn3rEMKfaXg/NfLNKgVut0yk0qR5ttc7QJEV0fGuOy8X+Gg6CyLg5U90fvcBe
C2ZcQ/QXsELfbnPsMHi4LcKT3PdD/HC58gpyjyA+LYFPdujxWHyQsrDOQXUX6lTy+iniCpJBycCo
ys/q77A4eLMYav6r6hYt8R8IlpgC0Ea38Gwpsk5cRX4CdWGS4jeVA+2jJEexXUOKDlPfSuB5ah+c
dID5SG6ninEXvNcRbK/kl7A6Bmyexo0c8nsM6xSOEsjNYDwXx6Q2m1KnXDGZEqccncU9INsXlmXo
GHxhX43vmQrc17OQcrstfCwo9MgbmvltkTcU22CQwMe4LkzuQj292eQ6ApRktFbXk8wD6SH8rTPc
mpNiuVBBPW067CmgiEvfKR8tOLG4m1tAaXf4nWB1EfM6eklS+Jbhwd4nZIt/BzxJ89yIOV2+m0+B
Ti1GvuhNKl+Vxq5Rq18GIutJLAjIqBpXVqv+eNXQLgEMAv1OU8ELR5c+5lHhw8a5ZdSrJW7kjyLt
Tyq/RHLE7ZobaYgiwVB57Wel5cfsRF6xZ49ebCPVMRVRJpbVBoLpHl+t27OYHxsd1fCumqKlLNqs
wLIV2UeOfCXEFsG3GPugXO+Z7anmF+I5P4RdY1RZfy7IwEgxwL5vAUixpWQUFNABAAnt6KjZ5d7X
rj2a+0euhkn3a1nuVpR2RVQr8keXm5WvJFvHQbin/VvBtcdX4MRpx1+8+oWhX8yi/Zn/8y1usGZ6
Y2ucOq30t1vG0yhLqhulj/RIh488I1MP8mWXMZBtcnF/KOoc5l/oJrwZ+WNn89fQK6HvcXA1MfGf
DYFXAyDHT4tEbZg5YxwUxS5GPiqIXhi9f+xBQrtCDoonlkbJ9ikOfJDrezLgAbzf+GytK0MugnBE
NlWbP28j2VnsEGVDIKNCmB0VmmABSLkArI6NJeZKFmSxqskJyRqd8M863O2m/Z3FOf5KXTljKioY
clnEUBQ6CZIbgHUPqdHuaI1PWUlEnpgG6ejMJ0evB+OkY47OpyyYiz0Af+yd8DzzwHY7c/l1Meaz
PmxJzC+S1hBzTFO6fFb2Vfcisb6HCmrS73KKGyMxBLpApyCDMp6TnPer3iExxwDZ80gD/FAg/0Fa
282twDOJe3lPGtIu9ynSaC9oew00CnFZFMqmMrdkA8Y+3jzBWvG+wv+f0Guorbmbhiw3wkan8Yef
HhcCbz3ObWSjVMQ2C9HJjQlA2ca27RggTU486B3x7axxXUuc0i4T2JKUo44vuTaMLrb+mo2XhVQL
+M9SYq+On0wB1x8MtIyG6GmbWlHl/6xUZYwhseKsQ8XAJ5irj/75UZGemcF8BWRCNw7WMlpc/8IE
9hrP8/+oci4CoGu7dl+zE3Kov+SIn7I0xAkZHf2X+rG5MXm7moP53BizuB5Fl9tlbFCEmMcNQEHI
BPP1aPqipbEYQJR+1i7MD4W66HyHRml+v9B1EdJsrxqlcNcQCuweCBK0Jl7GGeJ81eS+Ku2y1HgC
WUUhnRfuGPSi6iSo9aJF90khs5muK7kBqWLKNl3lIsbZxJNMuJYo4c5XCKalxrCPR1TXbwYRYFui
z6P+XZSoYYgR/T72b+C5TqULnlWTZiTEDSCwKxdC0NFx20Z9ADOTwNfssi4SMq2TGhI8EkG0k5v4
czw4R1yMHZv29WUT3C9mjlsP/5R44LvTdEIxjW5g8Hv5w1FMYr9KhSTcQ/DzIEMIkRxaWQvZnEJb
xjqVHuXcUrB+/f3PiItcGb9GnUf2aTGIaEfwsv6TcMJiiTVMyjXW9U7yfS+S1f6oX1YJ7ky/oNrQ
lgS8Gw8n7lvrHsgq5q5kbrx5qub7op0mQ/EydKT8wQXicyR0+qXt+HMvq5S+4eDaa23VI95sTiIb
T9Tiau2g0JiGqnaOmxBPOnB/g6H4UDV4t2E/YkHN9gTgw6gRV+naa10OvektcU9kIw9tji9pCs6v
fuu0xid5+MC2bcS7rzQVenx3S3YrOtSX73VegmLE0TdPuY59tEAiXn8qNG4bcWDpMXY1/1/++/o+
zHCtzz4IdvucYbG7BdnHzY7O4gRCpvIG/Bq2BzcO53NRSmVTNpDtRBJLKBsrOmdJ6oQJX890BQvt
aMj4M2J7wI+qPz4Ax2ywY4gUFIyETIM/JTSbiY83Msw7C0Fg80n/L1Xyn1U/t2rEST35ykHqInBs
uakX2/gZB2GPn7G0SRX5PIggmwwTyrAnDqP2yye4S8/J1IU6xu4f51HDSD3g+LWEyOIk9DdruYlx
qfcBbyWlciS3sXd6TzW7sDSSowxa+VhNy8RI8jFjDzlWI8qNV9khZADVqtFJ1DmkqRo2HilBM6RQ
1wte77lbfJwSKQQWK1lWjMTlFOAREobvogo+2bGei5OMqyIjsq0LCjysVWIX98moQB9tmx41S4aW
NaaZkq/wqK9J76MeWdjh301KvhWd5z8ZThd7Nuzd/bCl7X8pGPllA6s/BVlAEqoGRNkFG5yymrJ+
vnTLE88+a0g0IqVrIezKnk4B7W6K5gQu6ptB6T5HX6dTum18JEqxUm2t6qQqwQ6Rv35XviHUcY1S
dWrCE0x3E8G08y45Wh+bLfcoM9/MKXWPy9wsfHJGCthbaqTpHa4cn39+t8O8xtGeqsvunR1bdb1g
/Zy1PjsiSWLncR6I4ABm7ECjRznJ/PfV/aKAtXRjDkNGyFw0tgPW3hwGMPXnvNT70H2AL4Uo723j
9ZM8JNjOS0hI9BkXjho9/GibC9IpEr1pF+4QSgXeprTYZ3zQPvxUB3jTRoN1yqhmjFLzBFewqkOk
p0HDnMrGKnQ+2drcgzCSPhdl5eFnoFSXQaj1cGUXbkp2+iBZfbX1jNFmkbVH4bJV0Qp1LOvosR3x
/76bzx46maxGq4teiwu9Z5AlU3js8tp9f8gEFGptOyiYMiYpf3FbqFM4uJfCeMh6soYfaFmb0+Xi
S4tDsYHqzMPKFpOYUEoxitVyP9rbJeQXSHJK6E504wIXgUaU/rX/Z6VPnubCx8RHUT/cOY40boh4
hu5s9suVuds4R21AB93wNkZElebH+S+vCkhBbxOhug2viiDtZlANSOTeEn6jyzlft7i7E3nIFBAb
s1Kp8JyKcWpY3pm2Mtd5LNbfaSmU0iSZvoUSaCAdVPJaZyNHlAED7ZL3AC3aeBqo9VY+7F46PA64
EqMuJG4vwYi+WEIoF+fY4grzYPl6tpZAf3EkEoNvW/JtGCAktCdVSaXQVhuj8Wx3IpmQ1fof4OqT
If4i5wex7VSltFLnh7GoRIuahB+FzwA/S+VGnBzcXwlNXJuJClNUrtmjKFnddaQwW/xUJPLO/Qkw
Y62tzouSFnV9q9VLnwBSLFbUOTkfy7D+e3+x6jx+A1Gmus6m0LzJ1oGVEm4uYW5Jeu1WA2BWSNZE
ruKpuiJeJXdSVHv8rguk9QkRD1fyYgwJvsWRiWEyWMqiDtzd6RU6jsnJr/QHGYrdYsAUc8GtLn9Q
Im2OkMEdIIhcuzMkyoX7rzthSdsw+TnhkZDPK033U74NOymmTflq7DLoC9CcpzJmB4+kUrEyWLlI
TMkWIVUe2DvV3LVVa3+lFicRa4xkXHDwR9FzbeazY7jKMfjJtAYKzHglsfCYSd73uAaogz23mt4q
MdhgiUOc+wmEDSZ2z3wnfpL7X6InfFcmjUJ6Txqvjsj8mTBpN7NuOO5yW68KEPT1wZCQvByvAnhn
ufhbxfV6oLp/YrSpL3zHvUgpruaOGoguoZ8ukRdq+HzdqTAvO8TipkgKRb1Cpu4e9yfFULV1VRpq
sNF2Vd8UTTXEg1FHlD2awhG0z57L0uTRH3eEvrNUbnB51IycdNYT1fB7yQQv+//4GCSM3ZDRH1BC
UF+UxT3+2yXZFdyfPUCZ0CAe5R1sMpDeZC5ZabsO4/KFRdg7RtBOd8UG6BH2g0MZSe5sLD7Bjn1L
yQF6qfx59im5TkX4r3nX3KORdprHN68R9Ag/Aa8rPr94mk6VXPj4vyXs+JR3TCsfz3n1QtoX3r3r
f0t/DAelRy1HmA+3vrEko2pI5kVoLgXXp0gfq7g3Nzc3wBcrsi6lp/SqDd2cx3Jdxo7spz8Sf1nq
dHovttr9X3XzgotDJJ8oWCDh30mASuZhUdZay4ZUf9/hbvymfCkUPbJ6PY6PYPhrvZCky1/pEFcg
hC9Z47g/BR+N5HX4oIEKNgblI82Og0ksvVpV7c5l2SO3scTe5X3V9Sx/C0ZcZMw/BUr+hXj4tXeP
4WGkLPuguIv8i113J8p+4Jq0QP1Pq1eSmUVRf67KUkQiSD9D+ep1BSi4ddVbRe0nFbtTm3yQrQsh
kHfA48eZJdIrl2W/tsCVYpnNKHIhEDcLXTf8XuyE5lWMV4L+tWov70TibZVtqSQxXCqctj/mSQ8W
cDf1P49qXYa9ehkyuKv9kYAGwmsEkfPcE5YIu63yPe22l6DDNmcDyOCR8jnJmod36EE3F1T1IKJt
NQ2cNm9M+WZmGzWTtdfqU/SuQjGwF1VVeTO9wUgrEtgIV/HlP1VRLCzMInxIXPlmtDudPZCgdM5H
JSjnWqkHDoKs86kUUu56zQdj/cfHOZCR4Qm4NBCfYNYHHag+z15m2eGTUPkeEyyC46ff1StnhYMM
WfYkN3FCtGocQKPvvRkds/2yXRT73cQAxuSx6oUz9Mp9Re2v23nWRcc9JeYXCf7fukqv1c8iFZvn
Pxa6rfJZ+BJRuAUBr4t0rB2H+L8XPTiUX10oFeetjiD5fW1RKF09MXAndxEpw0T7A4bEP+pxo4Ik
qDqYOHm8WKL61F6BZ01xWrgosphtupZWEH3lIhtTKfROScKR6BASm6c8EcaMdmfrpU2JTPMTi7bw
ic3nOQ0dw+3S5bR31Xb06VejfOuZboLKlnGQVFpMt7c31fPsS9mu3zaoYGfyEkiqtJAga/1gnEL2
VqP4+5toKXEnYfwbyCeRltYUKSM+IrBIyz9/OICEIjx5fNRcUyeFJeTcxmlRZ0+DHZM55lQGpYKR
ETFWQ7g+3nOIO6Kj13GdZ9Im+ZEs+WfrlSIaRH0IGaTstgk113rp7roKLKu+OC0xFruVwNeox0hq
b1Vu1qB4vfYQ4wbT9o1jBvJbAOyRPreKviXkOQsXKUmouO4DdIWG6kYxGHa7yIRXR3omnBcNaV48
ytyZG0bWt6B1JN66PaEdgPjceSHxnHGUYwXkiqSmVs6RJhEg2uKLMSTvx7NUQNIejHQJFerNY0T9
Ot8gOUKsuFYRMDt+yvedWevvS1jFkGz2CfaA5WU6C4Beb/2LsUZS529jE1fAlchy/9X0f6dVgDaH
0C9dTQOI/yZZtAKzqjOhEf0lRZgJN4/r1tRFtRZGmJe8jK0/n2wxQG5SHKBjWYzkaEjZfiuK+jXE
kxQBameqbsQqrBeyexF1D2Pn9OZKzZ2Aa6jRA53rQgAA5lYfw6EwPP+PLJhofeMAk2saFsXl95Rb
6l2Nc1RKc38HMSECCCZIPJ9XPq9frQiINzypotTGtp6N1IkfOfG4He1vNCxs5I87tzNpWdrEyxvd
aMZuQ6H/rRuqRVw+D+W4Qzqig6u+wNfT+XM2uTUX6V1cOZKYA959jAdPkrL/OwLThWyoKFb6UkLQ
jOY11IrWgRNU42Kq+RExNtNQPVqiM164El5a7MCz6oljMeQvkXsW/+Z2bJc/ACG/LId9bzzy41GA
EC/oekWZrqzfTUvz4IZ5tl8rrIX7QM/MPRELZwOqRQ6s/968y7mwU/M5RK0qYsG+pgPYrIgYii36
yv1cR+/uF+eG/4KejYJ33GWNK3cQwttFl9t8Aq+yop6vXDRAU9xcYEMLWBlaYcNf6pTOWTY4nrgY
zceUcM+EZL0giBlZIjGk42+Fo/6YjKNIprDYu6VCSte85RhouBdJMqE2DaRJM8hvE+m7uNRQPmK6
hAlwxcAHPCX5g98krsirgAiwJlyWduzZYoLmg92TFy5bS9zxkIMCcRZHA135h8xNAUcJLSr39HWK
siDc5zoGxI3aOk1v57buSNMRI3igJGvm4bdN3+IUAuHL47w13/hRYNnMl6LPmS48/RRM9BFjkVlW
6F2pIXYFl5HUzhxtfr59jHjM6vqOi4Zr28zuuPAcsXL1bqv4L8Eu2cA7AAAvpvTuJ+vaopkQo8EU
5EjzjMKH7KOkk5PP+YrXiqifh3nmur+S4TKJ3AV7cXSNHPwvL5PZk5437WOjBP8r9ODtEbLkXLlH
hkQirKsJz2Iecp8zl+pp/SklvTq8JSSVJ73AbEQkeplSKA/q/wYNJs5rTjZA+XtwpCLoKt8PGpWQ
GnDyGSuuDZmMo5gB3fs5eT/5rmVmoJHcuU6WBRarHgdd/XcPiMBynD5eyL1mEBRVoXpjRatsC1si
K4lxlBosbaLJ/YcrpXfOrUfuwVrEO+vT5ly6CQEsERzyqOXuFoFDV1g3DM7tkLGum/b5CPfgitq1
VHzXtxLtihlFOgvW2JPLn949vqG2Dh1p+epFHbJMX0A3Muw018SOLpgR2XcYT5cS86S/55Ja0XEr
bIve+QadYIYZRoX6S8laRESQ8ZH81yZdSb62INTaqBu0+5Brj1MJwHfbW0fid468EA2/40ZJsm0Y
fBI4YDbsG1pTRALRIE6HBN6X0KacP1o9R/qBshfiWUCZAkFw/xQSKDIcTaBqAaZxQDi+/6TNrEsk
lMJx2rnlbfAjMPi9ETTi3AZ9C73fmaoxhgeXdf2Qe8/fD/MEhQxzeFeu+HtbVEK/lci/8evOyhar
/qsF4HgZlgRymJAgISZ4Tvp2CKcwOkV9UoGt0XinKEdPwHqtkl26us0VW6RAbj4+2tCRe3zbwWdm
nhVIzJtuHOeBOjnehSNrHuZXuAhe9V7M8I/XULwVhfsfJDNGZ448/Df65g2+M+O/qsI8TLCqbcxi
GZYFXg1OtB37uU0GuHS2fSGrF1efjFgN6McpQbn57Zr1f9Bz/Dr169QHETxnvHaiUAHMoXbhoiFO
FmOE0SxkkAmNLVilSCFtIKwrq8FsJ2C45cH+TtQDQsQ3qNVS1+Bd5f8RBEghaQPLUAMqwYtS7iro
Uy2A7lqMoX6wJxXz+WfSclXSCbAR1nTbhXTvGZKE6i6jEpVbp4hsZRDBsPD5SY9q/h3ICXuKOhPl
W56C8MVLojqxzVA9DBzFzzJJJm0kRaAnRdhnFjCqKEsraevrXYVP9hzIFfwzVVvwnzinxHLq6gBt
atwo5J1LMWU7rQisIlJDB40LdoYhSfNcHFFEkan4Hd/MhKj1EKJJAB+kfmUWbcR5QVwlSL/a4rpE
1Qg08HsK2xWkxD0Qq2WabjmdHCa2ZJSV1CMZdargg3KuFLWxipBwo8gZMHuzhNqIQwbQ9Dkzehox
AkBAOA22W6Ru3rAyLMBtwI+2Ccul2t5pa8XrFFesPfjHFdapaD0+HZ39Y28hdSlsIOAYPfuyTSWd
zxaWdnUmArm99Lxk5UBybHPT+EFKYA9+BrKUQZGHsiYD1zlvqk/eHcYgHXN3oeslEVBzuVJiy3j9
5PhFG1TbowvhULtMSDBw2E5dStdJTWCK4W+JkLLqv6pYV2rBZWSP4QaLDYIsyhucNnhQukug/nSU
rcdLoB8ypgSCxSAy/Gdfn8M5LSyBFzLDW+5XZnHHrZja7+u2//GKNzQVORjSLG9rAMAlGDo+IcY2
VCqJZBQftws6HY6AzdXZwjvDYSJNl0G45UVHkqBFfjsd4OSwEqlJ0KxbRdCyIK+l/2i+qqevWL2D
wEHBAewxNntC+xAWLqOKZirPfeu92lVGHAmw+iI45qCV9OB+fU38zUXLQK6qBVFBhnJWi2JwkQf9
CNjqdnYHTjD5V02rd1L+0IKAxE8LRTHLdj0LYCC4AOqhmA7bhG3U/ksXwcQ2MSv4UPdvXGivVMLg
/NK/B+vWWh6Par5+I/LVLlp5MRf9Y2cIYLDtzYqEBEM6agAdTfPe2zsVQDgZ89ZrBYldb4tz5Qq8
DcgM0RM9/yR4xRZbB+in7ABs7UMpvjMuGi4/QyqkiicKhFwAQzt8G2329dflphww3PYYkSdciK5A
cT7eUQVCsgk0XKAp7v71HiAsdBXiD21GzSDD+KMG4/kXZy0FL85LPTTSvlxk9bttHjtJW5MCMOsV
CvE+iDCoD00cuktO0d/rhifxadwPiXVkPxg3cct4ktyy7TY4KGBm7+apLHrEjWW1C1tUnDJJW+po
SDraPyQEZvpRIIlvdrArUBqOViklCuPUCjR27+PQs442FoKkw4iA66+TdLq/Y8kDanRnTNDy4qpZ
OvVyXSw/Y7x3vxtOyHivsnDU2qgAafCt1/cH7xtXXHaBzlz+qs5wJawxsZFCIsr/2r36z6M1RTWS
J7fkeJdHnnxTHiUWxq1U5XZ95Wk20TzS5ly/yYej0iX70V4DccG5/ecSpR6wZO79u6CFzRjiHDiT
8qBv847MqlyQbZ9T0YdkRi7KL7abcoA7IVDxWTZhA1ek+ZyvrfJl2Og7uB6pk2DOOZ/OsdSAi5uC
29NfhnXgKqe0TzkVzfXAMkiRuyDp74u+TB28NHDct1tZXqD3dXeqmZ3khlShnXHvlJM9Settl5tE
9P36RL5wpTL+0o7UHQ4gzDHkwj0IQuFZiwoECLKbSGqQp8zxuWcEtCodbMFANvsQMR/WitgxwMpa
uWsUH1RkjR2hJQ2ErIgsvdl2lJa6yQAVOianPrkIEPOAXhcnTrK7oIyTHlQZqrmLMyabvLSBNv8f
HSPrLoOx90PQHK7QLMXMYsD7yjCin2Mkb8FV5mAH9s5H2LHQlEq8cNUsY5jNBa3YOrlMsYi5SKkK
g601fsY3sF3vmCT1xwGDH2kcdAdwUwyDZZufkA/wT6JxlSagHMfuWSTtMovG54OMXz4gf3Yc1c59
hmF++FINvJDkXfJ7px7GYDuTstPJce+j9bogWmUjXrTamvy3aQdmeqgeaMfZVPPQ7zBs7dfTUkj5
mDjBCGXJRIIUlap6m34y6dCiJ1a0QQOGpAFrUp9xdsbCFF7cMhc0ymK+grCPrtRu/u2nhEPBU+Hb
huO2RBDf51+tRdz2mVc1WxeAxF0LBlz0JCBinW14hGh6SPf2J4uswM6mFSQOjJkppcind5clEQfa
ZehKSYivPs0p2MYH4XMAA7dMGS6GV1NmjEzpJvmgtKPNaaNiYTE68GSpsNhu17UCZnizK6jE2nGm
x0MM7DmvA/OeMRnGmDwS6Ye8TtsfxydDkk244uxatMcFCfTZW7nW1DNE/M4MD6nQdDZR8chRf26c
ivCoWtHezxcQ9RAPPDnpGwaZ5VIFjhFu2MHwVrg6nB7lij+omRkhn2/CfcA7s44tPIlg10JrfKxl
xe80uNmAYutEakrZCyowQfqyprI5+pPG+PNtbUnJesZzFwP+keWOWPMM1vFskzflpnNUs8x/mAc7
//E1Okcv4/v1HRKymJKKaeHXzzZT7iK5NKyv8LzwEb8jjNIGyJmmEMjfIFfvTO6712wRlRsrmo94
UDtwmpbnAFGFGqDnvgeV+5bZ2Sneo/lxxIbIuZ6V7G+djpYp3FLxd7usTJiCSJngTXizDXI9cjGy
CNPBTtKTECUqtDG6LpYRQoRvkKa+YPL4F3lvg8z2uZGS/l+QyA3JRLp1Fd3t3QeK5hBzoDSMIuEE
4jwtDUtyZmsXXTeZHl+FucdSWmYWY9pW2f64QfpsFqcRjOFW0FxkRgLJ6oADhTRSvITwVApRhfbd
eEowyQqpuiA40pLcUtuq6ljDwu3wr7J3YCvI6YJpbgGHA3Ukn6eIeFn1ToWGFbDrJBDVcPR0/tVa
bH5de362HsVhnnUCJ4uWkQWPixwuDqbU4gxbMaDAFQhMK2jFLtRwuMwiBWsIjoCuWboh3t9eYPka
oz8pGC+/KE6d4j/xwciCwayMbba0ZigYWNZY0mSye0OstQcZhXX9C1eJNchQjLkkzobZN/BcESNe
CflQlmD47qre5aHpTlHlNqVVFfvqKRKR/sbsWbguovQYobe21cbmxezpPqO0zqbCcjE44Cqe+Sau
xq3oWDYoSCNePu6lLTXxDXw3VjTgCG9j1+mHzGrNcXIYRDZERFgdTUHoknoengjdBxgT4IoRhhid
9OwVbnkl6gxjkcDSMuoqlZR9M5kVHrOMPZGywuiq6qXgW18Oey1Vr/tJ+JCBjmop76kzZrkNnxd7
6lqyVNp2rDhHjQYDGUSAuXko3O5yfj9tE0AcTOV5grQALdNV/8w2XuDY3AupM+dSZo/nbzH5icmK
liA5rhI6khfQ42YmNY42UmdOJLfNOpgow4WuBwdYXtzZdv3KX/ASZFcvOvt+mo0UOjSQijRTKj04
BDYo9Q7ykUuJ+k1eViDrKlV4CDEn9VqNN5X6KunnYUcXFQNWzZM3dRz8qGHexA02ndNYQiNRSzxg
c2YOcrWVnSKbU3mIR7aXEW1DU4Q+OkyiMnVb2dX4cMmiAliJgGpOuGWNtqF8im046kXii+l5fKgC
Qde2sEq3G/QZPdSCSfdSQ2lBYhkPv8xEJkNmxuAtDbhFi61av59WT2nqgAqOBnf1OeQNRqzDQ+jk
kPgmF8Uq0uykJNz1CujQg1ib6cuchxU7n4P4mj6kWfaHP3iaIwZp96Sa23N40lM7PvYQ9/GlmXkQ
uY3obL6LuFkEe2UrDaI65wDz0dVogDSCmlNuuiTnPEUtgncyFRJVEECOKFFuGONyRwsJb5Uc4rbz
sVkZsgxgc2UuvkT8KNigq2fNjMRNcMNTVVn4Ru3A2jgy0dAgxfb3dWJewTgr4lZU2T2xopzh3hFV
gAzdv8Cr/B6tL2W6gYRZDQj1I9xc2piOB+1ChE24OJf1K6OSjk0ROob7yaawgvEL2IMuocqhQUil
9wTZmoFPd6zGSd+cibpjqoJLzUQ+KsDOjVLK2o7SLdlGsMVBqI8ZrC4f2Ws0FiXyIPlJuc4pPpR7
1gIzMm8xLNLCwmzx0ftSROgFK1iSbLKrGfAT/OYw5bu6Pb8brH3ohHsCb4cLy5yMB53DhOuPD5Vb
sHrxhQJOrrP/HHdTTKCG/XQsch/0OjyKXIdXsWDAYQHZM2KaJueiiybeuqInU8AkN2yBJ6tFnPex
4dj90Otvy1QlTuX/g2tOM3J8T082PFOl/4PoHtDDskdQxYSfwf9g1kDxajkBy7oWz2q1XGck1X86
6EW5EcTEcLZzXtyokR8eDGH6L5SuoP6n/0DOff/q3yQW6p4/TGAvwFfnxGRH4hi9zsnsqrV+rcDN
tCqR7AVUWG8CquSlRkhQ0fJ8XoS3dstmfgCDVqhx+O+fF2Jn8ZNugDjTezETsfxxXtgIw4nfv4Qf
hlp889Qu8rKhmJg8/9bT+tk+mj0ByqCkkBjLukczAObau9887MTBeEZ1AXyB+dWixZY6Oa4eCA+j
6FRga2bc7fZ8uo3Hgya8qDwN7ed9ccb+beajbTqgxFWPMD3xJbH7WXqRQHF9VuD9IgTDk2yrZE3h
t8pmo5lk0A8xtt/fUdM2Fjij/RzfrtdpWKe+XE3uPNTPSr2lg91PclYBZJCv3r8hLVANoVgNGABN
hVD45fzUzV4a8rbM8ul7/ymxLY6grDDSlN3oJpSm69wOCuOEOiXtwsvIgdTc0l42cUqP1YTokqf6
YXot0nYAye6G5yhxkKg+ukNBSOW9ksca9au6WKKDTg9/mfIR0KKpgUhsf5TtkrlGDofhyTrkN8Su
t8P0/wrzEWfFESa5UFfSi4b/STI2IRLaTmDtK3XMYd5YsDHgJwQ2u5WzJ+SycZ4Omwb1V5BIjKov
8WiLEP7mPed5wEiwIB/cRDp0UJWN540IPTlml8gybNRIBFKarOlYz61bbSDAvW30j4hNzJkQRCuP
hbPLHSEEncraDlBlmEx2z/0FKmz4XEZBg5Ddqx4aQzP9Y+KI2/dDXtlM0L9rdD6AACeJUkF1rTBv
5n1igIRxjUQWUNJa7GPgqg4MP7CJoZezsvPcOLjkSRTPcRCeGTMkVnnRtXhJv0NmWOQZvg1+ZZk2
WILedGaePdU5EiOtLeyBQhM/3vcLh0FC/yfCD/f4RIgCe5LJudtMxxsHQBE4fOEygZ0RlEFnEOcG
YuqLv3G1DUQ7bQ0Vi8iMni8RnSIIu4JBhZlOc5AThRmYHIu7EB9YIazpr+X+AM0CnIWF51C2xs7p
XXd8K7SDE/TSKiggQLvD1yB3g3/WnmjqJsm9vLZdmDnqlrI3srA4o8PdZYzEmY3CwCSYZE7Sjlp+
gK9i6nJpbw6L6IVQIosN7wWmGl1SSq1HA3HLva9sVBY4z2+nHN3/FKCVuxWP06wNJEdd0zGGBdip
OsNs6/vDK/n2T2Sf5f9tTNZYUvq39NdCe1AYnqKuRRJ5X7tHQJ1x/na92bZY9HJU57zxb5lmcn4Q
SDcamDjnMC9HnbwPRq1fqVO0IAqidblptqtwNFzR42ciPqpK1djc8V9aqHLCu9oGBZQGbVAcIwnR
8aW//EgL9bnOvcXjPVe8c6wjw+/QODaGylyg9Sv6hvb+Is9oH871AwPGqeap599y96I3qAwAMO+g
uSeoDfhLK1dRx/W9JtyHTiuzaOQXc/nLh7a8w9sFYQypcOkSmKZlmwYIfqox7ma3J3eIiFMNfq+m
Yoh2tZF2XduZdVrbEVg45dr7I4C8s1RgyHP2xoz9uKFoN3azojXfRuHjAoe+ugtvDCEFXC7+byGU
jvNBg9319phjkemzv7x0d1iul9KNxS1hYs8QhRkq8zQX3I1gptPqETt9ofloUkBnpmlwAiHsYiE7
IH9oKcx4mO9XcamBL5f8IHxAu27xVGCS+hDwe/JRE4XV+QbeFNXlh9sdpR48ePjAUOJugkBnugPo
zFtosi5qKeGTWEbUiHsbo2QAIREQ1jii2jzYdILjeZOKORNF07bK0zxBhHuHdyl0uTQ2MLLKE8aR
t8oCIXsne0VqT/2enK/qIpQQ8rhOKhA/cId8mKfBdp72MQdsfn2tm7aVQ+3gfB25UV2Eh0uIrt5S
Slhhzt7C1hCBWlT12YIGRa0Qn8X1HYGz9GSrgDfmpdU3YdwNsipqFfJ6vnd46SGckkJSg11toE7y
SeVjf1Nb/+/tOBQSSR4LLfUCRCspf1GdDqPe/GpgmX1K1WsbOG8rXV1/wculPhD9P/Pz8PmauUrV
PgT7ahTgZVY+IxJcLWGro4H5Hy5OfNEACQ9LZxj9jdx7erAd5aVcN5uT6gFf3cHC4qdIPT0uTzdR
KTMqt7k37Ou85vW2aBtrgrzTkuU/IRXhQU6hdjoAn8B1c5y4qHyJE4Csie4D6fCf16mOZfkCE1EH
TYvvKhWEWW0hqA4dKlEBN8L0dCOFQW2osb+kiXFIukBA6MCAx7h719Qm/b8i39p3Ek1Pa2fXvVI5
BVICxAzUKEQw4gftUQ18j7mLc8kbEa+Mr9Qwo8NPv3C7ISGI9LMrNT+dav3MQlV2ds6f21SQrN10
DGst/6BrZ2gf/Kn8i0A51t5jbYTChD3xYam1m7qisLbIGptSSly5DEHsqDcq6/JI5wiG0vShxLHC
I+PGhzn6z4IRfQ2SyRVQG9WlFGNNCrAUqU/a9eI4dF6ZUF20o//1uhLWcI78Vm1AiE8IYYjaRTfD
i0lwqAWsXbtUyZMwuEGnsTaXywQ8RjBtS4urdL9iGkMlHy2Nu95wXHEvYp9IVCq0n/fXg38f1KY0
NG9tZpAfkB7JsJDxpu91YCXE4S1OzZ5cR4jmaRFFbVWxtDers7eY0jl1/uDacCtMHUap1VmDOkRC
HL9ayeQusVHoMn72Iqd5YvXjoKoVv1D8fHJJBfAUkfkqUO7w6zOXmetJ0LqTfVS2Rc5AqOTRqFEw
Se9ly7Od0p+J7kYVelCRhED99dLE6h0c9ovP6HJjoskX0Ts61hkEbPHQX/PO6RdFH8Njw/rfZ1AW
nXsmJ7PC69TdgbegiNMuS8580raA+Q4vhGb6SzrWOknwnIB1LaNp+PyqbF41c22ZCa1GVQbvd6Fm
XBxn5gRw817jypT52ITh66KX06dHkweCsBJ09vi4z5yBSqdMAgvkpsa6hYP7ezJp/dyvMYUVtnyZ
V1VmiiHJgrjkWBUZDBvzh4Cd0bCegsIPIfgfAXn9dLrha9hFKzYw98EU9pO+ihM4e3S6C/9WHXXX
vzeVA5CTja9d66Re/z1E22h1Bmk/YjPNO9sCOAcGVE9OrELDE2rLK+f1ezggw6fPRlT02j8scYZY
2PqaVeXvUfJYLQXy25zC95Q0o7tmRWh0ufzb5riLIvLXGMS9UnUh12T0J7bHLK59k/AyUC8xWDr5
t5dbW6hkf/Eunb7YXRljiGrgCRmuJq0LnBZxms3J4fcViSISztvJkT62j6z4kaJjEHqRmpDrcMt9
9YbFHZHyOttdlA+mx5iEzI/S2iL5RLOjw60wN5LPQrZWZFr5b6iMCsmH1rp9lgb3IhU/H37PuELD
RgFLqQ5diXcyghMnmWI/gWNkCnmipxpPvK2EFebNBUbLx/oB4r92Kh8P3QxZ1GE12Pm4pgtj7b/j
iBhbZAB5D+5l8teesU8K+PjGcLIkG/FZwE7x5lR7iX9DOTi6Eu8hP+Yx42gy9m/zMd+84mKxzBPA
I9keyHqZDEhfg5+1y3minDT5EEl28MMjeMje9teIyuCblOwqfJTprqLPg17GXLV9TK/QVc6hb8bQ
8IjqFLWaomVGRGoaxLWuDerKnm3mc1XwZTzrBWoQ2CYwfIm5YrYzG1axL0igKMJWUnUn5LZAGfsu
bb0RLqCqglpA6i8Vz+69dkDd6dkpO1jssPfBMSFTveteKx4bWKXcXD1M8hmpKqbl4iV3niEZsQze
AYenPTmFEYDI4J4gOHB1hXqY66f2gz1I+JQJZdz1GcRUM67iIazt6X73HFR77ROu64q6HVub+MWf
G6iubcIQh+xQ6rvWHXvvVHiuBJaOvEkKVDiEFcwe7/FhoADgP0Ncy9XwkRR9WfMUTpG8vFUgT1B8
PUd4+Ab8IiCVMv2i7gXIPjVPiUXhl1ChNmSG+v7fqAmnND4bt4x1YM+udli2Y4se2UA0tcLkIMvc
MtVIuDYGhI0qbCLkG8gEhWUDdxbdTWPyQkY+qy/Jbs/Y26r0StKW1RJtPTyteSz1xlLVfm4uktwZ
L7Pv0uFudFD11WEg+otNrqKOSnAoj5vB2PnVU6LcoviMX/3Rw0uAxKd2EzWcYIsPfXF6/FWEpOO0
JEjFMD/wPlGsjs8g1K5dGjdrMZTN8GGHZiUusgQQu/sgaNNzeItH6PPYcdERtHeIajXhvai82UA3
x7wc31ovKl9D/DPVgY/h86x40Rd/eXYIBCfiV2rixfHTMAeTPMg06wjTL5wimyIjMCLNLKDpoWtV
mLLakFN6hTX9WVGO+8OT+4Dl0GZ6vR/B5kt6CKw/inLvQV3MH1Azs0wbYaprBvRdn3tLIkxbt5mx
iZokJK8+l9ijV8qmEru/Y0GCoUtFedzxAy44+CbewZZ73l54eWCZQX+IM/gGqwKExGpyyJ9wODho
C//+IN7uzoFU0G+4SYlXSmmz9q80LBBiulOmZy308GefqvRDhCX0fJw7ZxnjAQ1JHAR7okum0MSt
EF8wELvjyERB9l55WBfxF389aIEQs9FgLv9Nk4XAD3gN01ojIklBohd3+fsG4+N8x6bQMpmdy7q/
4aSrVPfyHTEakjZCZi1n2RX/t6dcj3PNbaml8VQm/iKik9p+M6GfzstWyqCuN0c2xGCUocZgiPZT
8bWsnKwYlX2FIpNW4KLD+g/URafBdLwAZbsVIgPthqHXVsMe74R+Jn4TBvqzNO68omWA5yRa/ZLr
8lIRw2KXEsqHhBabwv3PC2YTlV9XRu4TCV+Yp3z6A8wBtnmL7VCBZyqpqWzrP/fh+qOaTcL2buFo
A46Ny81QWbvrqB4D5fVbQZjz9/NHAOUYtYIZn3LYqZoRdZw9w4x+wQu2CTIqZh5GDcU69X5AcACm
UHvNxrmMq6arYjvTHkDDhR8+m+j8KaEj3ySyTOAFAuWIy+eUYlEEIg+IPoh3sw5aQTJiBJg7ipjD
Y1rPCApsAPnNjGWlrzt81DZc7LrmHyX9YRcte0clv2r2/NOE+d2/v0vBoZ1j9EsZaRyiowv6e9uN
BurFLFa06yes/8QOOe87ycgR4Na90NEHvZwtkHWb451b0EcAMOpkhMqVV9BDsB/5Mrh1EBWbC76v
+UXJwgm4K5Mihp2eHeNVBmXlPyOy1z/4xZ84dIYd99rUomvaS+9ilRljlTHMBW/kMyx/nNBgA+UL
fveUTIU3QO8aIYwYbSY8JJpq4izWjXf3Z+X0LSvsWpDdh7G1jpOJpWEenvDOLrSJCTJXtF/bQ/uD
IpDFPf1XayT2+B6/L6vxtrtpSU8anbqRSzpPuU2zJb2DTzCrvYTMi0DdpDP3Ing/F7C7V0iZuUvV
jxprfZe+ySP8ILKVXBweSj40M2CwfzsUUI8HlIlyFQSU00MhfiP1DTG0SEinF+djPq63a8mzgSvR
5PY2squ6tJd+yt5DZ81Z42aFmP3OtOjVhMeFilW69sxP8PfZBEcyIDugAdILE+V3fLNLKkMyiFo6
XyGvzGfNMALCN2Yvwo93OHLhXxg5Y9b8DkPk1UYER4NNx7pxfgzUu6GLv+bLYc5mPnvYfmzISjm5
EwguZ63q4UJ5I1lzVdMuxCqil3B/ZB7fKmKHOpLALw6BI7+Qb0B+heGe7RKqCB5SJhJeBx44SByW
JVMSJt8irtiDu64cNKxR+BDRpH2MzFY+jKxYwQe/qOPxyTKHz+Cu5q3Yd9+5Olg7jKhc5bo5SAYj
LBZs+ydtFzEKMuPiTHWaOc0bvSW1vbXTJd7HDhU8lr4SWukRYnfKFj3teWFDXxN7fgO5rtRWWzI6
/OAEVJiyC5YJMV7dS8WuYr3gJjcl5b787D3w7Ukmq1ieZGna59B0PL2gei1rd/6hGb5XUBO3ovv3
hldQofpTYWV4kGXnscTomcE2UcySQQ4n9XPvX1t68wUdek4qwY8+3MbYvaa67BUJ8f1ItQHhO3gO
NML6vcWRm9S+iYDsm7s21ucRb++jWOSHaDsmW3p7zEWwW7EM/zqy2miqsftdy8WIaT0/YETlgONu
bClfXvm2k6hTKRUy4FUl5gE4oz8QZ3X3Xb4mp9cMCMQPKVh28KU6Djc7Xg5E5PzxgDvWPoGZjQgZ
jhyI6g55wyQqaJNjM7Md1BGbTq8zLb8iDFLP1BUeUMs+eTbCW3+zDOlHRfqEQlltNIxORVbutb/r
aCXiTatYp4r88lQPFOmYjNl51tb/gZScqQ9Dl9nE2OggbqmBh5Ksg4miaKNrzj7vE5QIr2bezo5X
UAfVlPchphzqwzzp8g6Gxu474zrf2/pA7BL0T6X7y6P3JfEADkS8VCUUvoksrny02gLmauTYz3AW
13YIRFxj1/g4kFZpJhf4svFGwnH+7n6WWkLFVcweNxqR8SWcIZzAPebUfO/wgiPrG2vsVkif7Ds2
JgyO3DgsB9bpUNXW1NAHMwR1mlw9prp1hUdW1Rx/hnmE/8bzFe9GHyISeoc1OgrZlMtW7KVgnSQX
5rV6maCV5yynqbk2giAAO+oJQbBjgU3y09ENPQQGBEEzVlJRudWaPzgdOfq3noUDhhYD+aAtXAvx
EI0qvZUbEN7TrKZbJKJzQAPijpskApwX00puBH5/2byZY5QPzllgOConMoqKEBAlOXQRUIaVS30g
Web4snCU3ghbjIPjF+qUP1D8YMvTWAyplYMwjung1ulCdgs66t7Lztk5+OVyIkkOIw7yAIJqBB1C
qo6IehBNe46iDMdjNnDIs22ykf2zxg2b0e63EJPMojB2iSD2+FguBZVMmtDPt0pBUS2yf3j6UHpU
V0aek+KFwYTfRw3XEWzgCjyfPjpGQatf1ZLn2GycTH6N88T6l3Qp+Lp8KYiMGdOlgXherhE5ZGzS
Tkm4S/ajjx1Wqziw/UAFjrX05Hlng3XCBHQfkmMB2OqtDIUa0YsSPmy/Lh9QlZ83IwsBeU5STzw5
u6kdw5paIoprqB0TjgDxsEUPYGICbYS26cwx7Li8MeKjyl0yAZWd/Er5w+Eb0BykeWYjdJGZD6Oc
HPjzd8juBkaZ34ebWeCzyZcRxFcDlkzAsYji8i6SJ+H+oIyP1+4NX4GfdMWpxaUcWxH5+8fkNTdC
IgI96q+g/xnXvHnOLIr3irj3WQq1r5LVDIlhn4kHZPNXS+K/oLHYmBjXXBmIJBhjQ0mvLVWCdPsP
m8WRB306iwsoMqRTcytBhdLWTy06gU3B94SNii5kdY+BizaTomh0X+3wpO0MtY1zgUHZrjii6cT0
5E76sVn8CU2UFcYsZfgpCpSJUVTKG+F4GrAK6qnHhHzWNze6kLcdiN7HRpCMY9Mu5SFcCfLkJvkw
2v5NgEMlKN4UVj+EUcT6Jws/YOhhMrno6PsGJEnWsrysAErN/psmvvkKUWzWXOnVmeqCW7LEFEY8
ID3HsMc1O2JBaeSc4tILY3l9LgQsM1MJGQqtrXyBkAocqa5z7tNTe7184smEDFInhHCJCVih9xml
+x4wzzUL2IwveAlsbCe42dz+Y3jU51KxJ3170MeNQHKRG4Iqr9C/KQUQbrsUbp524Wdc4zbgQnlM
BrbyJ15luNEAQQmdYXzCwnwuvAAdctmxuMTM/tNo/HWGYhBcx+4foS0CzqdRzwojFVhP43zeevg9
V92J2msLKrMXiRGVdmPsMkI3fFxeEZISXaXd4YyaCno5kTX5CiEReG9tvF7702IWE9koBdFOBZcR
2qbX2CYDeZ3DHEYu/aIEaDdeCRcJ4VocoFyvWNahbaAm+hKL4mzPQm9kClLxyc7Kj+FvJ99a/XS7
3+Rm5ppYjMYEBZoXfVgdQrzqorLl8YAjx4gfwoJIW7z7hh9akww+uhbSZTwgNkw0DgzL9UMJsjMA
a5F+HoXziH3wVm5TohsEiw5ODErkTdg7/VNLic/55W+mAwKKIWVIuZa7N4ozMuFJS56dyEmlVlxU
yhd388FuX9eXp9PUXPlCWHoYG8r3xnQiqq47Co9b9Mm2wLDG48zYL/cFMRAs/xKXlvjpnZmoDUAp
/KICeYw2q/jrI1tof85YRvUVkd/NBAFwQYNkvL9ON8dBaVXTJ2POJBFWlHbGgbQFe8tMhW01jstq
qY2t/9tus1uvIDrbOFybFhggi2Oo3CprL7czhOhgyJ2ENV1SUQ0Yi7XFqaamymYQlWkTscQhNZPS
KSzDVTz41SOsoIclCySoDwrQroSchazeHq3UXym9KYMkM/fO2k0rq2QAfWOtm2nQYWYrQfGlVGGx
bgrBGqiQORZdoVHh5B5fZTHY0jmK7Hqo5abR8si0F5GlbE5mRqiXXXTzcwxHzySYytlD2JgndYi8
hkHuKiyyzm7bqLNvvc9sihjAihLUsHV2QIKiECpSWEqi4DmrSasv7W+05CzNM1+cPBTRWxdFV5hn
EywDCMMb1CkwiXMxHIbnI92QHPcK6/ZayKSCT2orLRgrqTYmDmRXFls9fN95RC0ZKGzPSKYJ+KSp
v3qCk2niZoDvi01TgBE/8R9QAnliGlUQSWqc6Dh+0dUc88HafUCjfe0MF9iWTt2fuQsrnZBk8i4T
/jC9v9TKoXyl9DZnRVCrH2blEOiywWRQAnnwdLp+Bk9G1iOdiO/UkSOqH+zg5ORekvpNX/UHmvC3
wa+EEOtkDvQvxtFxxU9/9cPWZfbo6UdOmoLO7VW9Lv186iQirXL5WtyWig0NeYzcPL3uK6S2EPcb
dCXX8YummivrT6GydhATWB5Pnwoq7f0NwmHWo2vuC9GvpIROsGpsrK9ItM0azw408TssBY7Irgj4
JymR461WqjwHTEQOLxUAP2T9gTI1a/XQRoGFzgiFgp7F4WpotK+CfIF40sX2ALejUa7HsYOK/VBk
3ZYkNlB8o5zOc8omNQHZ6CKRRl0a8/4uVX39cyuTPZZMNAnWnrKya88dLJl50ZuFo4GawtYgjfpi
3Wlxo6GYZOjZajIvymi8i9J9T0OOihQ170HhECudOFNDXCnV+W9n5kZYfxfe27GQoww2l2MMukBp
XMF0QSjdtMcw61uDjPOD2PXj+aoYCcg7uRoko/bsSY5hskFmWBFJk/mzxn2C+bvZXHC5e8ObfAi4
gmkmW//bJTYWiGlqwrr3CPvpJS6jKMDRHcv/donMxT7iQeVBSOATLROjp6spXIRaOVkRBvS7pYnM
6CsQya8HEqJPLQK3A+azdtJplS8KE+yfcKYUGBoEJQlN/+X25NCCxttXAyFlNnsVa0zbVaJ/rxZT
XZpe6AsH05wJ3xPh6wXud3Cr9wnrB5JwG9igTx/4jUyzWN9BYPu5oR4antRRV7lwfV52oJ7e0ZEi
u0mbkD6FDwCGYbK5C0/0zdL2MEXtrsD7CTzjbjE2HTkXXK0EEcHmW7u1IAbp+yr4YRQwTMiw7qjO
FBPcuBiV65eOiyYLgsDVdzx6+m9ItaqgGU2TjKk3X3s9t6P+s0j4qGTJUWmBSrHB6Y+l+N61cR+Z
09//zJSygnDbD+fiZDBjMpvv5WbqRLChq4wB/HE69AGjJMZbIa1VuqFK0Ztgipe1UAu8S8waxY4H
gReRsiMJ+Brik2dviBLFpH8gQHeGTh9dPMxK4HWipSbSaMt4qmsZzsrLQEEe6Cc08VT496Fmtsvf
njB/e2Q7/+uXla4JIFUBiG7xgJnkPNVz9WTYsaM/uYKHw9osxo3rxnVdtjPCLxDgRAvcaBhBsi/f
bVg0z+2EmsoPMJLHKHVBXUEwF22cUgp0hcDTp5OuTSMmwKoxXVZ5FkJmmDLoAk2sUCjL7jHcCfvq
iuQ3eMz1UIV3v0we6hRc+IcDLPQzoqZCGjcbVa/2jA2bya6N8ohC6Ka2wHC52D2lIJYIc0N8spxN
CPIcA3qey6fW5YR23+NZFL1sLUxWZpEwmbzdYPHWZFg7UF8BDDiyhNrfdOS20hkCX/QahfjSlM5+
YhLW/x1QdtB4DTPCjM2PsIs5yMREbDGhE1N/w9GEdsGMhaeLfqJedytUg6wFp08xNiX2z4kgAB5f
MdoAHckhmBzQ98Yk4We7C4ITTTZkS6iMn6Oz9hgMunRi2Hnn1IQZbvWpWk/6WJvRYnV+PjzlPVyd
7Rhxb5r4XVsMP2qOAx6GBIZ9nS8DP1/ZEJP3/d72XGTqKkWWylh8EFb/+KfovIDFJc9BYTt+WBGk
1eGK4kIc9llVx/73HY3hVRAjKx67aS2pMgTVgHVscBlQPcGyFSyWLYj2Eg5jSHuJf7/8cS/wZDuq
RFjT/Suer8eGYjN18o09RhsaCKra2zwJIMq9/oh+Wp3jA+Ls5jR2JuxXk9RBDmnIelo2XD0cGpzC
Axpq6GkT10V1wTDMlnLsT63iR0oJOd5J+QUv0bDbU5zUtx8vMkNt31efFcrC7qCYPA4UddGg9H8o
62E0njX9dZ1WPFE/J7s71hZjkfwlmsr7248loWJ5deJbUhq34PpIAthw10cpnnjILk14Z2tZHPu+
AgmQ/K2vU8nlXkrZb/O7eqI3eWqiYjLhrcc3FwvNcKQ7yX6kIWP62ozaW7qRKT0F6lxWbr0sVnBt
nagZpxU4w5cZCb6a1zC6DbU9puyXVka2iCmCF81MxFGM+sMUTtKHhqUzy9ul/MHA+KHBZ+c5twfX
bKGVDqmNlVfroqqgE6luuzv//dSqacDmq+k+jj7V/r2jd0qS5jPbMKVSqCXfezcEH7yRMyO5wOjV
z5PuIJd07tZVETAN8D6OudcarT66HzK0gGlo+WGuDf2bIev7E6FRrRWSqn0VldOeryLmuqFlj8nF
4QyH0ub6ndjzOzZME40zbRuFSF423uwfpMvN+CIijxt00EWXPyMEc+oxwjlWLpLK+L+DcmuH5VsH
0O0f1YFIpjdyS/hZUeuBbR+WgHnCnL4EvyMebF+UCIw3ZoL5arI6my6kTJVs/Jd38dDoyLyRJT6l
E4Ekz5IsKhr+kadQeWCJVwv1zwYaJ/K3YXKNx0GHjNYFalqvz8ao2LkAi0huHkGjHDxCtFo/Tdts
qtLnmJ7bZ/FkSWa74Hc7CljTlrDmixqxeyHLTiitrGEW2T3BSpcFeJ5qUh5z2mwhmQY9RIzanCQQ
5JGQDXbPDiWatEZJjEfbWf7z805VFnicCBIZFBA4LTvOP4pZ32FEeY+ZTdbi8XNolpjy6fKd+spc
OfpLmquJYjzaxAVX9LwFHli5xMaZ5bIu2Fb6q59CZQ6exQFy7uYoLtaH4qzHNYLwe3Bd5qaJcVA5
rG92uMirRe1WfHXxzUvRlOd/zm0DV+5Eeey9HZTBCHISqOgjIRFlpxqegnQxxLUkL7Ygw6F6oj5P
lQu/1VfRcFDvDr1EeFf9ZlqkQzJocXKQ5lp4ebCUh2DSpjfGrsfwqpA4KTAvml8avVVu+zgkc+Vx
HLQl33r3wGF6e1+WrNJAKnP8IAWX7Bot42deFIoSgKskSCRT218DCHo8DQy0VVEFtXaVhTcWOHtJ
Zz0FMP9gNcJKZLwBC4To32imGMHmPEOfZ3+M4TYIOIwIv4drwgZ2KFgGYhMADwMiQsuYJ2qVpYtv
dsRAMyMfFXDcyM2Ume+98cqcH0a51e5ClLPYpfiJWFz4dzEY5Su1g1NSi0lvl/VtHvgnBYw+5dAT
G+pu292jwsuI77IHATcMqdWtWV7wMlErHx6Qf233M7/Wu/H5np7i1Z5Xzkpy+azX8Xzrn93b8etz
H8+LjibYIQLd8USJYalHRfibgTyxGeI4fI/fIBeyC4BTKfq3oOFmUkOMImAIm51ta6FBY9KbMd98
aDzeFMEsv8ZoAgodG099P2HyBQdaOgkRfgSjKHgwrRanqa4UcZ5MGHZEjItkcReVvWV3vO9izQ8B
ZYOTLII5Rf0Tf6q4mdYFB576rKxc5PRr62m/5s0lPpYzri96KIcnzfnPTkuazVwphG+iEeWCWtnh
XmyZFkBUubnJWGEG1ybHHQ5L8auRHdSaYv+F/AVI4h7AeNxK95TNjR+UPcVNZvFSOibrr2xVfPYk
lTt1uiDItrkHPxDuUnbAtqDTHFciJmumM1a6r2K8potBiyHgmu+l3spBccVhXpcBHY4Uq6n5NMVj
h+Q1vqKjmVrochSew9myKT52IZY8kqIGdkG1DDp1MHsceyYg7Qc3Vk+qJwKBRP9SOISB1LyFflss
z9bIhwxRpSvXfcQaaYPAmo9ZiZJN7sZhXoq0HEQgElR4Yd6T2NstzcHB0KnkxLM3adeohlw7JntU
HOyBfEAlg3eGyEixQ9SYyjbsPCkHUXHlMqEEaQS9Weh2TwPLjfhFE6BLa6CFdC4W/RmRdxOpPHyk
m6Ii7ueCCXvWsSaDp1s0Be4rHgxX7OU18fyA2T37ey73IevKhTHr0Sdp9Jp5oGiSpVAqgFcpyw2J
ZT5S6da9T1oi1T+Zwuz95Uc4Vq+6fDxz9btINILryGLb8YmCALsDk1lF5LE+D5AHmYAB/E/5GvYj
3MuGS8VN9dObS/NXmEDR+eoTelwiXE4FAI+vlEj8PlOJggxVq+skVMtEtuKOAF9akoEwmx7gu/eB
Ks5y527Jzvv1Rbo/l66pXKYe5aFDFIkK2jNbHpF05ADNyLTmZj7cSjuyqFzRyUHXfznNOiXa6CmW
Gtjb/mJOvMpbKtII1pJpu9IIoa1aCBqpEXF3td1AMtFYo25ay14oKPL93GCB+kdzv8SSOzbJiCUu
Q8v4FFcTzwQjEHtUaOjdo27pUqBuUna/9Rnwf2DsU3owQPLfkKhwbE/jhoD3RPM+j3RZU2VVAJQj
tda3lLnGSdeoGRWmpG8GL65HPNDAPuyx7/H3ketNWU5a3ygDbH0ABtT7QZwBMj7eDW1BrU4C4BvV
g4eUHrh4DVyBmUNwvdLmzBIS8vikHeNHlDMcRALKdLuhzKPhm9fFMbNdETg8cDonQtItfV6woail
V+Ax3QlLpgPle3DNTZxnUAYzMZpkiFh/V6DhJ9+CNw06qJyZAFTXDWaI63Ui17xKD/6RuctMBXYi
BhHriwWpkTJA6ODd1Wn5vwJnnQokiSy0GZkAYhxq1e5luCqN6Euz1tWnw0tTUJDD1dsIUg2B3VjF
yFWDfoSJru6TbEWz6DOBhkTycmm/KeFqVjP6ZI2KD4uq34NgaAaoTKpjwge7q4SKQZ08mHEQJchu
UsQiZJ9Z/SE4UBFIwp5Moi8SxtN7Y3TcgVHtOPRx8CqIcZAKTQR7nu63ciZDAAxEyEAV8FLpABV8
23Omae1XseaxoptQU1c0x+a2fEMjOayONLMbUJifJUmysMeWkVMKH/nNaC0ehpxTZJUnPnsDHihN
sDT43ytS2u8Y9hDIKdmSTux1OhVUcSBruWoLvSf/2FjrOusTubgwORGlPH46dGA63/lKfy7tk6Dm
lOjW2FKlBf2zIS0sxJza0kmQ0J5503db+8lTDxYxlNN6nFssqBwGWRGcaWPWBEQeUM+n0t3HvoC2
L1KsivpY7EvI92CqR2PxCJWR21X0Wl29ugWm9HBIRMbgSDom9vVKPXock58CgbnpbCN7A7LF+0wt
HDNUzxEPtRgbNjzdMuXCW5paHDP6Aeq1YdFdg++LCSdF1EpTO47c2VcvmmWM3KzScD/S8J5Hz9f5
fjTfIpAtzgTifG+RaUBMVHc8eoeFNbTfXK9Y6Ye8A01BiEKoVACn9sgO/P6nsWhVZyhmbRi9LpVr
NwMcn5LorYv70hxdZIGjbXJ9UVTz/5V+yMbdZWDNZW5Nz/JyZ+WepJLJUpPCYloif6RkjTgI1k/X
Cj33cFeO6gZGK+1nLYuocZk9+O1yW3AEza8knOh/UcCeeJWeDREgFHFXNN+ctK0hamTSAsmV6ort
MHgqNnoMmMga89/wJEmC1XLIR4v7fZFqEkienWhcXtRmhrB6YOwyo0Mk5C1wE7fpdiFx9xkWi7V2
H7PZR5X5S2eZ4nZlKkEsYkNlYy/7UJrXX9ZLrPTyO0JQ/VvqKj0Qr1oFlK4cRhwQPGPQrOUvPob8
M3G/R9sX0M7e4RMKvHMRKhiYExB5QVCfBIfJboHt1rJSrawgwr1xCMxHQDyBupEYYRFf1kqLC2cc
V82OCuak0Qhn+5b2pSBHwMC41NOWRqDqAMtK8vVbat9Zc+WFqwfXC9XDH7WlldMOWqe2Rk4LjjTV
hm4bTiAZgiOD4trGIZ4oF6BIJuy/GBusFd0MYMYYy9zTg/hVBV9UpTKRpM7vV9CCtt0dc+mcNqz4
YdCC6kj5w1a+oBSviWdCIICoT0tU/IgXHAM5TRbSWASNoKchqwfLhb2rEbUY8usG9eOYanlDubR9
DrnVELyCmGCAMSgIEmbxgWOS1bg1roJJvayK4XWvWZjHFHxEl3gD01nN0x7q3ToVei90dC+lzE4f
3KIk1adSmNPLp5L6q0RJ18OVNi+JRfA6wX8uZ7hm6iM4HXxWzaxjLkSzQC3wIC+XIsHtXp7HcuAH
OaV0BWxiy/MSsHKm6KLIAvHQUAImJEU0W3j7Kr0k5eqGNpKtexQ/GMMQyjA0DkWPs+dO77vQDcwD
u7iH5Z8KBBisnVyGg2fzYVaTQgWWPvZlhoXboW3vSSToxzxOhhAxgSldQFbwVXG3doe8hs6sLgdS
/SBQU41ZDXtR2rweJsxCwUyHvvsA+AjDyIaJqhZmApBauOih8KqfFiOhits/tAY1BVnI9MXbOWh3
OsEamcsBEMjc5YWKYmZoqr9bp3j6WCcBguRdjXxl/5a9xPgv8lgYuQdw7ADRxf7w57h9jCkpDDQx
xvNDWgQzM987WuZcSqCHaIWHQM+KaXyzeXIV45rqbqY15FwiIoymms1YZ5cnj6qaMKaNAQhkh84y
fIC9fqhw2fD+XgXTRJe6hqsxfygJNa7k1YtbUbHj6Bc6RdsYynoykKD29eJHoAJuhf75VS2XUPFq
cqJ3MVl2exMHNPgkIOTUGJZIz6MFV8N4xMLKl6cWYLKGFV6mBLI9SGAv//U819ZsMF82/Bof8Cli
02yQ5KGLeiUsmbi63V0ac0yxuJaH6vnqb6CYDgn5jSsCDg6sFSlXVaUeiItHAcbPkQdIRIDUfCiQ
cwBfkTaviMEmlZL7DaYj7quz580TGzQXfQbVUC1Cksl++26EJc/kLkNnqFoin7l1r6g/zwVD4G5S
ZkaL9uxCIiCwqM+uoYQvmIyZas6W0g1dNpw07eJSVfVUwd/4ArnajhytZxNdkJrABw6FO0ZbFi2L
GghHVPyI2NdPl+ol/ojHFhUCKJ33vW9I+s7+9wVUFiIvDy9kDaA09eQyINy8DdcfSwuj3Brlrj90
oPT6l8EZKg362D1V5tA51XwA4e/2OetZWdTWOhO0bxzdM8zrDf95Ay6XdpVELi48fXSfsRa8VO9e
xXzVc4kjD4LRjiY9aqwa2yqf1rpIAN/+YPp4Fll+zlpPMx+bEOs7qnRs+g9r3nt9otwlw+dZpcCk
Ch4ZvfPhyS28jZEf1jKZgkzgyXDA72NxdXH55Yer1wvvzy8Evh4/6WgF36aplPahKqY1omf/6mtR
ZIw4QKietELXWBuid9+XW4ZqSj8x57vh42LPASNh9sycUmN/i3WztaFshE4fEbUQlV/MydRTygCx
NypsiGt+311zSm21Kjp4jNUmVUJSCXPLXWtPKdvi7RP0r7TrmEPmV4VrwIYifrZFx6uO9XFCqGw3
UqYG5GE0JTISCkJif4DizAQF1NvM4Dtp/WfhXpHBLWSjQHF+yjWdnR1ZbGWanExAJwKG7UTwj6f5
MGoCSrSL2rz7aTClfRhfaweaofD8eW9OslkaBv5VlPBNSgrLblpT56k++152YjIEnD8lfCbWhrGz
B3wtXvxnHkwMgKaMssstg0OtHmV49AQoapwSHLOg+V6+FDwTGLYRbT6G/Xin8kCwDAF7vVn1Tpdy
i/A1deTwFIsJawQt5oL5W6iytyO5fANW+RsKaEE3IicqCDwZoRm/nU3ahuGNxfkQeZP0bH91ry5A
Y6IMSstw2wrgaHFGO3yuhhKEVzWInyyVfSSpG0jz1schaFsUJBoXPm0ceMpWB7OOYH7mEn+cmFYn
gc5pr4PC1nWuyO2dlP8/3tHyyzZdsQ112v3/6U2Xu4z0xPWx1Kom2BitpDezy+LYNIDTIpdIJ/Sd
g7bH19VUPyqqWuPRC0eDF49IRMfBTCQnDa6n0O2KVqY2dD1T5BAar4hP0vOtpcKtJCHebv1zVG2s
rfKZfW6cJOoZo0eeH1aqTae1RPCDR5S1u3mA+6CnjDy36i4E3gYc4XelfA8o9c+eXZF8u0bWoIOi
F6/WfBgqzcNWBw31HziGYReJZ83AUTmfqZSxVGJWpEA7MpjXwOl5qwwdt0cHtiahzUPjfIhnlhuV
4GlZrckoSoawi35IjgyQM6n7kCS4sCak+5rAc3rvkhh54K33cfBRLfYEG/TUrv4kwHmSEjFvnXqK
n5iPP9JdKNBdUkMJsrQxR7QeR+udmapSaHfNTIvV0Bt/JQJFqVLPTt+Ev35UMImvqKguETcRRttY
fW+9XrZwTrbE36cxgStnzhROn7P1Tm2LgoDyEhmFq/MK9t7bd7MbY5evWDVhhThWx+IuCEdM3hmr
KRPFtSMB0pCG19bPd3fNXbtRQldt49FpWCAzRi/ncFjT1LFupp9CKMhhVUhrnoDTscsrhrVS5vrw
maNMYLHDGSWhTHGovR6OP+X9tSg5SK8ClAjhPOlE2TPtPM6CsoX4Qk+JOb++QjJ8Np08EzYjvTX4
bBl2ydRK/SRBoBKRDmjnCAk2XKZ5mD3wPV5ALpdUX/biUOTc1zsmEbWXRqAoWHRlWUPA9vjf4quK
u30pnefgA4vofU9FMiZcJ9DvEIBC2H6AXFXI7aiKwqZ79kV///X6D72Cppgw+BbxWFj/nXRAZOqz
TCpuCWnrGYGQk4ZmoIJa2WYvDMdkznPxvfIFMAOF76Ien6ZF2g8V8ccF1Jv2fNDOGslOd4mOqHIA
ghyF5kNGGr83eHXpPKwaRToojLcu0uwz7p9qjEhgai57hWHtTbSDSn1017lwi873jfvKZccF3pdi
Q4O5BIR0Lt07YNK1vYlIfmzv3aqoSQKisQ4lmlrb6kO2Wp4ecL2CKCCRZkeKyi6qWelo+njJZKCF
nMXv0GNwT3qyGPLwrgK9yTkr8cQmxJ2QCo36pqWzJTxnwNZQ+L1cM2cBOxK/kEk5pOXPJaRfK+RW
Qlfz+aSbXSDjKux6QncDUAv/S2W0eQDPiLfhU3Q8grBpcy29qzG0kFG/ysVonSoy9+BDzjDD1Jtm
+Sth32bXodJHbkYzEDO7gFPVKNfkxdmNgq5XXvWvIAV2SEJhf3h6ktaToHxE5oVs/b7RO35s9U4g
S5lIzFLl81fcczVGUxrUoydWcqhz8OMqhvdxFJD74C97rAq2PRK+nSd6rQw9+S2jhQNlGdtDM9Dt
No7Imh5al0htbd0RnAd5kprFSZvf3TVp4I/+cDDndyhcvEK1irl6zWbSJh5yOuhjS/MmWH/3hCje
UIy2c+ZNahg7AaJLR5swolVVMuk2NXN3K/VormP6S3nH0h3VS5Jxf7JcO2BLJMFEXVAhBoXLrbP3
Sz14TKXEUWNAOL07Yo8rjdRB3aFzV18MJlyPVLBv6hi8yTTza35IOOT+lp3ffm56KKDmr/cLHaF9
JloZrYnOv8sqzWPTkeBK0AO/SFdkJ4I/EzWIVe923/Y0A+vz3fmRAPlcxrM6tvL4KV7vXNcltwmO
k2+QGHH4LhB+bz9OSfc1D3ic/sG4heiKiRJxtGz57SNe4butq96FjUDoPrjpOt6Hy1FjG6oAIoKX
f8D0BuJGOjbTXVcVa2eZGggPUesNSO2hhqd6WZXQqNKcX7ETcy6sYvJNZRlaPCGlPlXiVALEndR9
C2fgKtrcNRKVusWtwArx50uuZ0hQLhtrD7Dhsq9S+UqYkJ/z2Ilw2Qufrrhdo9LO3AX7DHAK8WKT
Pyzd7B1u4WwMpn1XurJaeeZxwE22rGjsCL+diYlYnj0TIjpTGQvmDRDNeiS4fG+Hnn1RHj4pVFjp
1bNBViOLT2JQww8+pKNM2XbKIrCGaFP3+X+1oc6jOt6MEa4XehPm1hJPym/eKC798GJMSa42Fwx/
IS/OPSPEpt7znTU6FgahhSU2Sad+/nMCQpJlg/Nzjs89seAr6ONjBdQxi8fUu2rxjhUIdhUiaC+x
E4of46XjV2EG6PTNWtBjDQRStYxpQrtd/VT/O6xeIcBdIHdZp3eeKAd3CAHYfvq+LW/cHZJNfcwJ
UxZu1nHeY4DQyA2+EVKfro7OkX7lxU/nJqBMi2paDQMRfniG7062aFNN6HulRtkocc91SMI2xkGE
Ri8RGgjz+tjdrLt8SL70yqq1GAvqbQLA8dcgODI5tYePVboGTRUX6GNZkppSCYV899JtHABaMepy
MpNM6C9jxOqyfllv2STt523VK19RH7pAdsASc6RLlbFXv7pSEiYW14NxCslI2QYXcKVgmLY+o+8A
0LLT3eOmcAof6bRA54sUtev1uB8Yiji5C+BID7MKVtbrQINHMDE7MHbcTtItS5NcWLPRMG5UJLfA
PpTbgkQ8GHtFA62M+CUX2XRcThU1d105I1HjRDmaX6skSDp+aHIcYR49j4mQy4qNc1Gide+JJvFp
1yW2WJGr/QOlCEflcdjxY6WQU890aQT7KdBdxbASqnt8G7PYuwMfBifEy7JLAnsloYe08Hef27pT
UAAdLcHpQYlBpMGd7ENAfbPeov8l7aYHa1pJ3LUbe7y06QQzmQr5eZX6glWdVxUtS6nhKNHJKXst
JmwHTPP5z7hQMvCrY3PHAR7VgwhhuW1tysMZQhtMVtbAe9pkYuRzi1cWLqaq4KtVTBZUU814WiJ7
8B82/rwDIRvSZ8xVCovMMPoLHWfMSMxR6PGuN1L//9V3i/o7wsgKdXHHLb2ZHwmegeJ4EgNVGWb8
h8URMINEvjwhwG1ss1y3KTBrbHYrdmqnQQjodpEqsQXQGFe8NOv1nCwcHsv6tL/GFrd/mf2B7H8Z
9Ioj9gV+9ioQWv2D9Mrb9uIvDFA+mz05AmWxyaIl7fyrXf7g0/FxmyrfubDO4x7rumaT7xoS9nnq
dNp1biD3nfd/qgVEwR0Gl1bILPGhBahaTFWceIMCF2kJkmWD9cbyFc1ZDBcgVBFxwrYpR5+SxA+l
S0dhUL3sa0eDZTch54bJB/0AINgqUno/tmI3kuJK/LTRv0+2xiV1WMEDteXNaAZ4b2A42jn74l8e
D/KESk9uRd7ryEU3J8LIZlSyVtOBRcGfmi+55sAiSCmKcLGMf1O49ajp45kutJov09No0p8pYwQI
m2Vr+g3AGHuZTGPr9US/HXRtnHxx8YDSnVs2DCo8WB19RzYb+VRzUw7c5kZc2Kr/7YbJ48GcdQzH
UUx0csHGievblb6xsEJE1GhDcWDzb3AaGee+ITMjbQ3jlmgzJlEwIG2FEoSOEcXDDDPTXvcO1ipF
aKbsruW4Wrp3nwM2oaP6mhnh/Rn81CD4yY+8X5fInUsv3zXe7yZlnb1UuM7oDN7QH5vJ5iXiYXw8
9EdmEurO1EdEya4K0DYckuBDQtN3op5hAbESU62cKPvJVH+23RDr79LyTtpy3ey3S/6d+65xBbmZ
GraV5NBmZCu8PxB8Osy5dVecocmKFE+CvSw2PoDXJV+ZQdO38Ttc6JlfwiDzkqJpQWxazzqFJIl7
F/UIwVA/P3VkJQAsxnkKlmbfdXQll3miDQ6ysZPJCCUZB71FDzPv7cjNSOPqYll+BOzwqqDptWSN
oIB6WHeqdMtnrLg7Gvv2RAyZjbBZuso241TY5OyHqwzuNDl7gS5A6c2aUCrKndSIdEaC4ty6t2cT
GyF1DL6Sgx8iUN4q+k7XJ0UeSo++w2sUQusSs14StlcgaMhaG6SXCqF14H13oZdA2Z1m0m/W5RV5
MNkrBuFgQeLitcYMPRua0SFGB8tgiqcm0sVyLD5QOZqMSkvGSro2jaNWDm6qh6Y5WCGPJsrqYJw0
xsa/ih0yYC+nkAfBvXLa7rBGtuI+IPxzo/Sb6AOwbOw/naOHRYGbAeCyOZLVvZTSvAWXJRfaRHzS
1xOxCeGld4HiRAup+WVShjc5DDOGeDWlokqA7an1WyaV2QfDb/fhTty2a2Mw4GkMw0GTwRTerwJT
6ctm7iXaQ13zUHZkGeAjTBfa8BtAnPZ0bFK4uWqRzhLSoPUwxxSj5PC/5CNWrnoarvmHfWvmlUpB
bqShdYeHxED/xKORb+EeAvXp0qKYRpTp2VgrW8sJejQ1R0hHxx+psm7B51mEbbTFLJBtnURaEwxg
uJ3cHI5AgrZxL1Dgd2eZDOntp7Sxwa/Y60XjK//qk5N9YvtT+XlQE4CoMlw05vQyu+Raog6vlNKs
tNCTGBKLT+s1cO8JUyKltHHp6PiSeAGPJf9nAEVCXC8t7S8VI8FSi3NxXJ/ByF0QYW7K17tjHVq8
QpO2vhBtVMiVd9wqEbVcoydk7E/azKRP2TMeWLVoFLnwHQIettmocB8WnBtR/kdAlO+InZUoOkBY
Q8k5ErMvsWMoPdDHHwXIzciPLoS3uJkdomZhS4R26Jv0AmIGtu3/baovkFue/P5AqBBfg/z1c4pz
Vshwp3F/eOuV4CvhZv2VpJBq+fQw8Q8p7mY24otNvxWWEswWafJXex7Yeo+7zvB7zNVoLTWxdpSE
S/VSs9AScSNoD+e6m4R16n6HkUzk3N6Q2BApTAN781Eh7dduj0ZncoCzRBqUSzpQGvOPxcO11U4f
DsQD97iY7t2ErhvnC9pcR8Zs6J1Wjf9Folt8oWRXB2eQCX1I/s7g5P8b7/3xzNB3cO1ySgBitg4S
MxHMoJAFR1GJOKrex31PlGPmq7v17y2fW6oc6DMSlGj8daaKaJMN/o6OqpPahfRbdSxXRaz5igyH
rs90ynSK0veoQdYaQHS8WxzmxqUFUSQYpwfehIlKgiiQGBqJpKhnnwfk1b/5ZTIad57racpC0L+j
j72D8OUIR4TzkZPOcrs5WC6sWzLsR95cIh8xRuvRS2vGDULNuqScXsj9LWjkCMR8XrC3hK/rSl5N
+WPyWJ0NYzsKUPCXL23Av2oKyvj8k5gcUPAIOs00gR1Kw4uqYD8+Fq/16lTsG2IWoU9Kiha8Y7u3
TD2F64Oi4AqoG5IZbj3RdntpAO/xRG0bd8ocoO3O9CL1qIfh9MPdj5PUvV9DoU0INcwiiPslq/Yt
nwRaGL3L4abVUie4H0Lqwqq8LnQJ6Ro2A5lIGBQb/+3YCpOkHAl+aXMozh4ZdiDvKSSs/vMOeU3u
k3tVNfCDxZRyCP3gbBo9R9M6l6b/cXNyPV740M6d+ArjorhwtGmNzWMtXvKDxTnNvskPqu0N7l9i
gQk34LB1Vkw9o6rPs/3ewsFacUUWH7MsXEOhMr0Do5KV280W/YjUzLIf73UoqP+v2dqwSUG/a5tN
1oybop0I1X7vNudAYwuRn+ReCK0VBlqdNyvIPkUq3fya4clJSv6iNUc5tXMYRojoTQIZi5DBOL2Z
U7oEECW15LXvqJstoSdj02BBEQy6nUpLalYOW3mrVtDRcOMCoa17sTC4oDwThGKeLLt4n8lpUlGt
iVaCohvRavGOpAwwshRBFLajS6ZpxMteIwN3B4E3d5uIgLFdaK+KjKMa9e4V5Wlx5sss92xzEc3w
rvJSmfmu3vCE23kVB5Vb9pdPt24tLKDeu7QuonxeoXXQzLSDNTkPNbRCKXHmIKX0HMPIlpqfLIPB
3jybD4+msOHZg5pCPFaw9pSM/9SFSWeCgHx+94fNof24ZFZakDMFvZBIT7x4dDbsAU3tgqlzZFin
m0Wsf5sgwrDgmz3h2xm06OqLiQ7Og1Qmo36mgLBrTSGB0e3znLuBCVoY5/G20z26NoW2ROUYN7js
868Srl3p9ktaxEDP+9RpgMG2ud+uS079g4dNsYbJUM1M1mKKHF5ToPXFvzZmdEQ2Clexk05K/feT
MIOEsBYgMX245LkZCo0OPb/4gHHXMn8JSdgH+Sjumm8BSuAFLV7bFLVDC7Si/m9Lqkh7N7krDOre
fZYR2blSqOwup3PTTesxXt9gw/N7kIO0Me8KY9yXxNgOCnxevBmIl18cvH+LIPnHD+dkaDRbXlJW
5iSxGy3PZRL/PwDHDENFJM5fpDAlqur2v29K7VaknVpvXj2AssXzAEaMiouF7/WW9VyCVDtd7LaN
RUsURq0CkCbPnK0c9uqVam3qka3Grxu3VWhhO/zYvowafIw5FnrzlRbUT+hlXKbnt77BTxP5dZBq
h4+2YhsFFMCXx+YbKkQ3iJWI9Symjs8A7VI4Nyi/5OtdFVoiNw4fUupUfBUHbxTRbB0t0lhkwQe5
KH4Hu+nKNbBDVHl0+t76/7iZVOchgAAjj8V0+a/ef1I8HN/iQKE9sLJFu9UOYHZqv9CA9lcM/iH8
jZt1/pKYk1DV4plwmdkb2W4Lt9ZvWpvgPa/tjiqLOJjDPTG275sM+Tnko6htGWZE8ZPWoBW209tk
YIueAR2C+dff3y850dzTkJtFCx0l5bsnjX0/f5wr04lzSifmwn05vGcOinFN0acxwcmQmimiHCsh
yNOzdMHve1Nq/tZDNlrX4Pt84dl+sB1+hA77HRvFedrlTI9aHI9sDjspf1t+TbaUTUtF7p8jZU3M
nBWA3gwyIULTTy2pY8wGkutKuSnThavWEmuOqtg5UlmiV9P8xYlMVL1LKGOpdfiCkS9aar/RXbxP
zlNQvgtlnRS4+EMjAqvFwtVmJp7uYbI/++5Y+1SQ52qgc5vIsBxg5HYYoHTCH+qq7Yu7ukgE2vKQ
bDipnJNOZQpMvzUXZSpawngoy4YFIC7HQEIJuC1mBbGKRYuy0FHg8jzj9C6YTaSWQoTnMDPpzgBY
uHSqk1KTHF+QxvuPlWVu//FR5I4yVSKgpQZqODp4U1HbxdimHris4n/0pRkw1RXB/LKqA32rbc9+
YDPqyFTQ/jKe5uaUdWbQZNaiwR1tYJ/80b3k3pN58ztDpZhlTOtgZ1DHAs33EJuGJB/bWPBHOVCi
PgpWaHwZD3C/eNN7sCOw45ADn+o6Uid3c68CWyFBwZ6J99KJkUdQ7LvlfEF81FOrYJgSvph3fFf3
jHJkm87TkJMNtrEwaGnQAMFIWmYUqupX6doUxVutuKSkPKnYo2eS+EOzLdFw7H7qtF7Trm+GRqUk
iqgTdRhcK7CedMS7W+C0At/Njm80dQfbH3oN3c9X8NEr4OpAVhHGaDZ3sYFD1CTrAlr/I+v+TDi/
GecywU7NUBvg0t/OI9Rp9kcOP3bD3A7lkgR6U/M2n/j1sZusd/LSNWJz8gVa8kG4zhPi7gJe6CJN
GpErX7LU2QQxbgoMLoZKDjiZaIuqCFVg93MaTTij1yZhTVwsW3cCq7BACE+31g19Tl8Mv3BzsEyi
oWbkFbj0WbBfoe+8/qzOgpWxWhDys0Mnq45KfKZSvPwwtqRj0nZNVSqq1JmP6KQqRpZRfqqek5ei
ZbCTqBTkSdDbKgCkfjz7W0Jlebg3DJq2vrKnssiDZLEwc/Po2rUtQBSh1S96QKvtVgC8FEAUifAN
A7Zdf5Iy/yjPSziRubAbFL6dfJ2FW6hNwxexUKadNLSPnZiPEIBEW3g6DRveJhoaY5hBaVRD9x4L
qgLfGK9A8TgOdzdGDw3lrMTeolZJbo9CWdZm9PjAqs8gc9CFKcqS8ii8Z4ySe6WWlsq4SyygI2EZ
WGN+MvcJMTtxOMt8gE5OQIKQDhUek9WcKdOSBPjOVgFDSStRSOsOPMRnDJy8+hTmrn8wH3n1FBFi
mqHzKskRoK5gpPMdO4eeoq5M1aECJ9GJJwCH6JtVECut2Zc9wQeMRz341RDrtqUtHrkOS8HxlkN6
LlVPXL3+Jdv8LFxLiatpfpKAyVld79StFrZG+VCtpRc8VngGNIltaF42cZUHKhzyKsiMf+rR+xx3
1hX06I6flJjCPMs71Z8GVqXIUD1CiN3sutnHzZkX8TiLqvOTcUX16OfIV3vmft20VhB49d1jFGJk
F8f9nwLA7K0EfxJj9BWICNi8AYI40ndJ0jt0xhIwojNKwY7f07+QPzbyz5cIg5ftP33oyvKp+DjE
RxhfOTTUpwGef9hdWHt3hXXLxvohUECvY8i15m2VQOL13sK71AOlXbn9aUZtt+XebEUpiwKTSkn+
QyXHFeRflK7MUKXTmcKttFPeoaU0QtFeiVHHmYcPhl0ZsF3ymXZjKoGc3v0zHD3HKHr2eDs2Xc6y
RNG+MKGAaJTohyBNQ5TkLentazpPvhPdt5MoYjBSd4qS6F+YW4h3gZNm+qXIcxEzP6nha7gKL3u2
2QCg8t7XjvIcOt7zKHNcyCGBriq28JTURJemTqLdRLQV0yGTreXcwYB+jTOZuzkWdLjjrNcXJj0G
6hJPh4gkEZZ1UeLJUNpaYECpT5RH9QPeTwGqJDQgt1FTvUL89AdaosZEm6U4wQ9smcW3yGpNFxfX
qOfN2irtAlYuP7d4OMlzmFe3U1NDV7X699OCw4EwU7vvIyhZlELrgxwrKusnWOixT0scXID28g7G
ENv2J+uoQ10LiZh6oTw6xKUkeGQkfFlgCUvmzzhW3JGc3w3OgevjOfs0x5FePHWq1xmpZ4Wm6G17
Q9WZShy3NS5gcraQxQXsNl9Omu2LZYBx4q/XhAtmPW2rF0/TXqBMNSifs2K71N76wGi7vWVSFjxy
aF/E+qiKc6Ssf0+aHM/kwNW8apUbdzOI3pIfVZofeF0VhK71BpeZBI+agBwnva+N9lRTGGBGq6KC
P7VgQyx4n1wRncbuHkojmRSQDu8h776PJjr5pilwKyv+FcUefkO7OhkfgAyx3lecS/cFCoeyakJd
PY8BIB+SnWE4RHz8snMgbqzgGHR8+qBxZzNk1Bu2ik5PZNkoGj6TRg1z4OLBOFPWfCB45oK+fv8x
3Plb55D1ZVtaiR34vKhMTXDL4IeegTssHLhOpU+x5Yq/bG3oCkb2zElj+NQHAMEhM9adEU/ybF/D
h568RWvV8K2XwJ7XhJ1Wmw0vAwLBOiJsvA5cRtCuHernygsSLZvGIwyR0pkAZetmVv68bHpsL4/8
zD1UbJIGkGyWBXCkX3rX7rGjD+ovF8RbCqOH5lot35QQd9luAfyQhI3Qct6K737Os/2iHA6IspyJ
LvO9GAwuWcWalMEO1sPjPxSAHLgDODrHf7bF6eTnTYJXCQxtLlbO1xJ/TSjtlGXDx8p1m/VUtwWC
LXPnIk7wVcP9ztshUztMqC85ETrKGnJ/SKRe7xuyEhxJeghm5qalKd2KB+0DaawTj/nfrWMniSCB
2/0CPXqxuxwqt5sx3wFunFBd3RFKhHq+svEzBkwTCudv3y1Qz6k1QFFZWmv4hDNJfVyiLOIht8f1
cp8h9zxGijc4GmWnTqTbUdPTj83WsgJlmILSxulBihiP4YKx8mUFV+r96LoEGnjzb+iW8abC2gev
dVP3VrbnbUAo+tkKGRkGg3vw5e94ZkJv4Dv+tiF7PKMF+c+YT1s4jKh1bkXwMuZEg67yn3p8kGDM
ouholzz9GZzte7VHidrNlIvC9HvKsvcg8hE9YVoe1eEO90LKi5FlQ46nxuE1omEO7O4wo1bnb9pE
t6EpdxMIAveH7II9whM2ys5NZC3GrWG0TyROknoeT6aHYMhOifcmrwyYNkh7QjpbXCgX4UmwKn2A
BPbRE6TXxF1K3cg+s1Kj+D76UKr4bodwIZx3He5VYRg4C8XnRjCTCWQpGOy8mJli7klp/+Hm0SRS
Ci83+QcQ+W+1USveB+Ar3Ia15J3z1bBUVKYVpiT2PQ3jE+30pevDyqeZbaa8v4jNe+lWplstfwRX
uEi7nwu91z5uh5qJztPnP+bsidHlAeK7DuypMAWO4W3ylh6h8EFEQwO4vGIF1zqEceprflWvyGQ+
B1xBeQGD/bWaDojZFmvU5Y3bFE6DgAoMV3rpXECNAf2dSN4EKOIbhJ5hpkBMMwmF5weJi/2AOWr8
l5f3MCxumbQl2kT3b/RMBuEJhSOJPpAav4kCeXGpeczmmg4HejPurNMpfEpVXuMY00D3Z2EHQGPj
v1OYQHbyNgvIZUBhK2uZDHBW7514gqcyFNnkd0GJ6BXXpv1JbdOnv1eZePUf2Nis43PAdNUB4P8d
uft+AYn+HAYTYNvAcgBPv1xDiXH32hIkiKJ/KKqSrwePsymLWuytEKaNmdLmla+srTUB/oc+H94S
HXQYphADinFuNcLHmPkyOXO8i54E7BZxat0j0HMrf3+Uwll5TVTouMNk9VFQ0CVMkywx1ELIfkTr
oOL7b+ASHk9V1EiPB3cx9NEDuSIWRdvMAOvs0jPijO+c49rXiniElqyM9DiOp6etvZwwRrsUcRCF
k++c0hPsqBtPjjd1XsrIBJ7fPzP914s5YOnycUZocj1F8SnM89ylXBHDptZnbsa6coQWBXcN4rg+
YXiMvEVFBqVF6Jpi8pbIARVfYmLN5LHJFHMdmCZvdS2Imy0uIFxvP/nue6BgJehQFWwwMeaKjMEG
wGns4XiF4mU959KVUUEQ6HZyPN12JEC8R2YC2DHXU26bLXeOUd39xZzns+4YRDo1+dx9Up3H7y73
1ngPEoc5WmWJB66oR2aOVxjIOH1PqQMg8lBJNNH68RVgsnfBqnK04Vkykltyq+iqw2kADOnlELLq
YlvskYezXomyz+bKTPN8QFJ8tAZHNtt3UBc4B+XeKRfB1NLzyaU8H46q6gBZ/dJeW+vriZ2gjz9z
gfEfVoT0YH3jwHCm5fVu6hyigjbjg5pHNCT9u+m2T2aNhcsggR/Jqxdpu8vVRmKZHJhlCCML9mt5
ExYC7Jpwrii2XwFdILAFxkHm4E+YpoKiAuF/KtmH8xZGp3Uv5OafRwzY4AyagVq7fZw3r2IGngrl
fPkQsVqX7CAnC8qcJ7DKYish87S/MVXkUHx+nq2JldIWwFG5NUn4dijnguPcQc5pQBHOKtUX+y+z
Dbvv+m/zyqBONAF8KqG4T22AuMP4nSIjFOq6zwfwYYDpew4gUrd/JXNr3KHALX97N5xMC25Scgl8
i2gCExQTDCQs/MN1oppfybokHZ7tD4NK9twSJhmR09M5fKqLNnx6gAyZ+SHD8/qjLSA1YVzkSLvv
CVJ31C5ux1wa7dDXmJr9LIfeWm8ON/Ce4Vehbndd7RZhWV/TXPa/SXgevFWAEEa6zSprB4abAUwd
RNlh/RGT/lwlvyFA6+0pC2PSE8J+1E/Q5qSqp1sNENFUia6hgdr+/+oiAAJrt9/nDlwMi3XQsduQ
93oE82V0wmhHqOP3d05+EdrfZMxE872H6MYnkI10sl+SKYxO+/JYD7xc7wmeGTdon4pzRq6bE/VN
IFyYz21s0OqZKcMep1Dkmpbu14d8EeiDqNHo8v+pnwbCwc0tpuro9y4mr+J8Vom6mal2il+tZBJ2
s98G3R8sRDsrIPq2uPwkuGtZ8ZmQMpipbFk1Et6YfKdJk0ib5sm6miDxzAn22HISUeWkOLY3vv7A
dxbPPmiezxYhl63e/HmtbgO8lhDYfsL6zT1WatOxvjL0FDjeQy4PIYkmc7s6i/NV7rupEVD14VVm
027ryMDu/3uh9LbOIRYJ+MfAbuWVjIy7wunIFpUw/AdEuIaaDyuHKil8cECNNAo1LVLAUYuofiNf
ILJ7oxeE2T8qaCOGSWPLnTnLB2q/lxtj6Gddhm5GdlgBmulX7sKj7eAFQugKmMtfLMdj07ykkd5I
7APgJffKIhqmEsX/Zi3BSH7m08H/ww0iE/DfHg2dOS73ZDscp1CLUA8gWBAuQlXb1CrrJf1asCAG
ulPsVgD4L8ViPvU62ubdo7QfiiZ0TqNCyfjSmL4tDxlOn1DbkspjBO5eUzRGkkTfs1wbG93YtHiY
DYXgzIca7U4Spw4p94s9+/Kd/iy80Q4OpSbX/hFuRRzkhH3snRg7EfluLVAmssfJgmKw5t4ROU8k
3fdBUl9RncJom+DSrZFFVCYaj1gg145/OUF04rYVruJQ8/LwOcahFKIbSjcnutQyCtFPievvdIyL
byrGImH5r3Zvt8j++LIu9AaLtY//IzfNXQ7nZ1vzHToKrVpMaJuIzAxDdUXvVfeeGn2F64ZjXqiF
5hjemqBxx/bJ83qsyO11/EGjR3vm0KaGfPzDMJ3ShwtX20GE2+BFb+xp3t+Kj4jYY9ZcaPpiHi1W
cvI9LCw8ssD4qNVsrHyyzySEyosjfbhHOn1qU5x7M+cszz+8T8D8Qm775ORZz4NLpoH5hojkfsUq
rORq8lNA2tOSWoZLOdlbQWSXVRCZF8eGJOJuWSHPt2CKYTG5rPxPc5WZMLms0YpIL8m2HZMbSvr5
3Hx1ynUiJGuCsM/jwKE5c3s/ljoENeyxCxImGsEwKKOAk+6Nnr3Sn5qria7PbS1Q4xRcV7jGM3zj
CXRNA23ITIaQ/u3uFB3W4wQJNwnoqfgwxv6PzqkGB40UuH3RmncopHZsK+ovlhpFadClXNWtsTWf
HrR7qk1KR2HEC+YfBwaFVpNlYKxbfFM0DDP+Tfx4IDGpAddNkXwWuZs3HAFgipCPhlp5SwICHJ66
YjU+OvQD1J4O79Xfwlexe4EREPJUx7ctkLDBrqneTpwGTPSIEWR+EzKraJ5sx8hljqscu0dy7J75
+Swl5ZEhEl9Z2bYiRAj/xQamJKTUeEr23Jx5pPyYHr4mnjBf60/+1gz7tl1bLjcaLXFZsoqliBgS
yY5UXvhXk7+oLMO1j3pcj1xu3orlOaCXqnfyJ4X0n61JmCwKMtTo1Is5v7zOHo5JFboc/rY8wXxU
ZSjZRFxoSbdKBCsv8MuKPcvW+Gp030AFmHco15SylngQlx73740uQvnF4sNJEb9LXFk4w+6syUQp
VJPszAChsKHEv71FV4cyGzvXkQdAdRaVApAp6+KTr9RgFOnCsg9pxk+DfzVeA6YAGi4ij+UeBCSH
iddBfnujDqISdfk36kTWqAQ+roJ07Fyvo4nYJxwIwtFRJR4+qr5fXykJHHevnLh6T/avpHskGpmA
ghkkCrQsYKFiYU2mHlrg3uHR6POYAQ8e2Etl7dURu44/vdfZjt+4uTcadXH5Y5ssP39aRbWQoN8D
Bk+hNre3ZsHDjIdl17gWEOuYBUccv5VVrf6k4suYeKbeosJ3KHpcxomkz97wNW7sLCsiD8vKgP/s
VpO3++QVi5qEOZnhtQPPL10v2NQ9uwslwofDMNs3Kg9kQVDoyAwuYZHzXnKai6fxlciFCbUEyoNq
YM/d/aA42Sh20bPmh4MLSu3fB50zP4JLXMeEiv3cu2r38GZ2TmoW+C0dQUvrxpZAPZ5/nmkncG0g
sfxKHpoJm6Eo+6CxlSH+uR3+x/CYHCtssJeivZNAXrcVPd5SHDQNbsEJvMVLTOlAg6PRDu0gIc+R
XpM1FAzrT1SEFezfYktZ7byxVK5ZxxD47UpFO5/4yDxvZnPkuE1daURJskagaHcRZVTch9CzG4jL
sG0wMBfxS8ilYIvw8FwvMI1xFV1Lh00Tn43ogBXvwTxpqycCHiID/l8tKfPKrFpnC4CJoEp004dm
V87Py+NyPRHHjya5DIvNuMLCpswYdKFk5Lu09mdgqOYaLSKwdk/SzwMVN4PgboCOB2GsekL6dPre
L71gRxQIm85PjWdYjNThc0ZSDKzC86o5kSZab3lw3BxVg6OaKi4/3yuBfaz50O5yDm2ckLl9YldS
/1KciYf1vjWNsd6oOPvlUHmTvplbW/LxDf4Hj0r7KWZ3V6QtM7C+FaofjRlPdPCZ/iN9ApfM5pHg
J26CcftM77CTCBIexPX6mrk3XS8vL0t2+Guu/vJhi9sZ/Kw3z49qd4j6jyVqJ486cAJ/h8JXmuyc
DmLcrViwo4jr/+v+8gQpARLugR/ZXDjtdz3W2eB1E1APJQrLioim2y81IhvSOPtaE1eUI1of2tDr
2KH1CeqKBjeJsQ2q4tJLHeQY+3wmiLLOtgFScgEitIVJgIDC2mVgEW0S+c5IgmNwnwR6NgQV8q0a
wtEmeI/mER/RdQf7IoD6DCvfAwxGRwR+kEAVb3x74YsFgiEpZdOwvrv1WsSHKv5MSZWMSS4FXU5h
IRHaY+JP8WwWsBNbIshgplHMcYnG0khl/1U+MNzaRIeEm/5+Gdh+rIIztbeXoRKQ9KpN139Mi39C
3bBIA9kRsexhB5zSE/bM+K3uitrNP7q5I37xPW1ayNVYZzUXlHUhtyhVUfXrTNh1AIQLGfOhbQRM
3hvtNr40BYA4KnaFQ4SRIHjC7luPQlXhCJ+Gbwg8xAHDFZwBzTUbPvNXoVDFc+7b9f95tlh4eDwA
Aa0Qnk9KCQQsmdQ5emA8gjrtCvtXSMssKmu2Pdu/3jlAsAkzrTJwgBXxao3f8kF9Vlr4+uOsy4bW
ALTXbMLueT2H5b+GN/JPjRUHo7vVdT98Cdll7D+viZA3Z5umZlswQ7KJjPSsapxGuS1IbjJ3vwAu
5dAdVv/fJb2nI/XUvreeB7r7o8BPecwaVmOBqjHgr2Rrwrg1i2Kk5eIbRtW9PfozXdLLF9IXDwP2
XHmk5D2Jfl7EZQAZsPXfkdWV2Jl6gHd53Fl/7lEB0iI7ilt7+tQQCjEhqfyQk4+DfBdDqbLc3Qsv
v+xxjVfxXuvxaP6gKLwxFxqXFBzp2lVsoAlGnQH/3g0uYzAuWP2jE95lKRU7ADbvvTg4gg/yxHtM
D7scYTqb016/1HnSPnC7+JYHF9epzLZV5f2/D8v6FmE4DAKwPP6LnzFQz+X8CiB+oyb76UQhN4w+
H1SYheIGVpfhV+uQgvbq0anEqeYOUe1iHTKyznj/l9wdY+m6wevBUCJRnmZk8GKs1lxmbSPdiwWM
3Y4h3tmIdxYjIQkPcG4GHVCB8Q2XZx7dodP5BG2T46F5X8afcv20KRQf/ltJz883vzcSOnITdwfw
Matbx+KmfLrBOdrCpmipr1Ea788sf15dJ8W1EpOyARtmdJts89wrHOnTjgPBiWJeUq+VaeKOBsdc
YYmFW09uQ5y7yBs/jTOr4lxdRxU8sO71WfK/m04RmHdacN0SJZZS+X04H90+RmawYaR17pWKHtf6
8tzDMQ+2GNo5nOlwBssrI8RAjweB4OyUiAcIF6/qbHM36MSE3ARrRX4ofOT/4kHE/Lzgn3zmDon7
cJBVwyxz9OEwJQaPf8GAl1uJKuZ3jOtfRtrwh6/4A1l4lN9CfcQENR9xF0qX/dtKmUyjB0WQdUR+
3M4UyAzopROPuEnOWWVbxK6tlK8eR4bMIThmmrWRujMajr36+UzEuOBjUU3yz/+e7qoDhmH3f5mX
yxZuCPvtyWY19NiR/mnYPf9309k6S/blFbwy33CuBcphVB1XjstCQPdRSgpzsbqpJDK3/IBL3Wrq
ze8XrM+gIHPesr6Z+hwZfR7/PUb2CNa7MhahdwMPQ7k7RkQm5FXAm0LcOOhg74LmwLpXXejF9hvN
pyeOu7oSdrt0sGIzxiI/14MrKSsZ90ST90JKOIyXbc/9WTMoOuiWqLG+U965Cu8UtXlFjIhHcMck
9LJWpBh4FrL4JtmyGzJl1hDMUXgpNQ1/S4XY6liLfjMqKuf1+hmuV1chiHMP1g7hRNyRCP8HZT7x
xenhPvCM2F2AHR6t9og4ANAXTOSO+Qo/2virSdi0GKpfqFnf+7O1deBB97nDYBPT2507PGzm92V7
D8SFoBmQyV4x3T8+oaRK10uMyA2zA9TNhIYuV+Rh3al4Wo+AtMseLKXWpB0AmoV2h/D5X6SnZnnV
0Pak8gTSMTyBU2nwM1v5S43+BwKpZ3H3C4qbzC/LGITtEvAYqwgAWQpjFd48e7K5CEmbyTqoRBCN
SIijd4yAPyMqztLU3yKgbziLDDcAa6VSqkzTxBVkdtGUD6y0i1j/++MNGW/Drr6LsuAZHCT0aLDu
YYKf5J/xZkCNeaT6t13XUab1pee2Ggzhw8xWxpLGnHPRSiGWCoUKYt0mFkJ8q//VhN+Sm/aoZEh1
YAWh+OUz6mR3wzmkUPpF7NoqHh9YPl6Ymzs1cqnvTqqVpxOINv/I1/uqwuiktL7Ee9nJp9MWXnpC
IzkmhyKKoP1UrM83/Kbf1Lg+lFC74rg0o8uWg6VddVnQYvzhTSzduE+gfbfeYPWFonmzqgLhP9uL
Yqoc4O+C3NhwSOuWV4jNNi92UL//d9GdwJGWEvdAHVvB1DBF1+b+tOg0khePW30Esgo0IkLuDRD3
iIqIQ9ybT0DUS5mWAtRbqEqkV71Ru9MdHFC+Ge6bXOqY84S/YT2k1Z5Xj1uKQHd+Nt3bI2NJOe9P
8stBEKrwV1fAZZDXPZ6V+elJs41kLdg+aNsb7NrYspNBDsczW0a448aXr4Dz07Utz5GxZkuMQRAs
8F9YsK2suA6qkSdX9g2tLfZYP1UTupSQKCPDjDj3ZBYEUybSubUnyDqp6CcYEWQ5Ju2sBSG7/tDH
Xd6zBAg1vsVijJpf2RTqLNXXGbBjJi2Dy/YrEUHIcmTkK6Av52P6R4Z+ANMzo52ZWfqeWhCjXfZH
ZVG7UBB0Xof0/RoSgkLS8hMvcV+4A5QBcfiblsIFiWr/Cs142ejR6uybdwUzbZla2elS+ARFwywu
3dGSzXwlHem2RTBoibgik2bDGKvrlMWL3c8N3dwT0y59DJSQEBfctuR31eRt6kOMjxs9Rdcp4DQv
VVKSpNTdbynBrwgFm6Ted131WtnanmWpCjNymIfkdC0h0LaQQoZ0E4O4OQSKhZJc10P/jE6vDbFb
lGDTNfCQEPfrpskscAR40v3yN3GvJOYL11l8UzrW0PzhFpclGcGQVQFMqyS26V2M3+nAarol0Kjj
GgnqRJyxpov5VhgPMep3/526WcT2K8mPRwpr9nRRztfEmRsRuauw7lAqVOSnadbVVd21e/GZORSC
XO3g5dqCVdLIAk6OI1YWreQ//FurLxExRwPIqZUC9VCGwcDyJhZe7S4nQNS9lvNb1fAVKgdNSTD+
zF2/lUjjstf8zz0y+AOOrfIorENFpE8iFIOfnM9qVOpqxlKgUMdTEFTNtbHkLCkcRjbE+mBN+QPM
LqCMQwSBa+wW+kptvBL0trofFBdKQ/QWXyava5piciDweKqCSmL6XzsyteV3YtH9gY+riJ38ORLe
ZJTDY/mGtbWSBJ31ZxBRn+dabh0h1X0sTwGs23dg0+QGBilWphJ+I1sQbHbunt9b6l5a2E3rlqNq
Qoh32X1BxuE3Oe6xqbyZZc9lXVlWNOG61EDA+mueimWDDC008dO7SqFNuwaRAIiAw2FbEF/XhhNO
tuzZlptZLcc4F6FVOBXi6vm7aZWz1hZ/OhH1eZQUqTkFWFkfS3i70fiUdErGqjrkrqB2yIfhKnQq
YYlervPZcxWxMInkuj8Ef3mp1M0cq2LQcrG2L17QYCBdouUZXcB/DG9zXZWWjP5T1cHJSYhxM8gp
fhiaBIYIx03Jp4F8ZNWcaVZCVXjTtW8ebAz/Y9AhWCqPiFqZ0wiq3jlfxfmihs+yJUKrNkgVpk6C
oPp5hlT2qH33J88ciQ90R9iD0JfcW4QEjOCSM80pKT3I0k/TCjuqKMilLdrtDP8GCQB91/WFpHbS
XhsybfdWckocEBqM6NauA5akGXjMOGLy3uchaKYQx4RdbuWUXZvKM5gFM4zlR4TgQFbFLrg+nglK
KRkiEr2W8yn9NBQmhHk0iMIO4+piQpnz7GN0v9m9bSY2P7XbRkNLjFlma6hWgEhIp/FhinbWqYmT
ThGfvl0tb4tY1ETBGoAaBnUY0tt+uTYOfAeTOz1tRuDj8YONlldEFGIxLJBdkgr3na2yRBt01iW3
w9JB+d1iyvATKdtybCOWJzJUZtW10l8iQpul7I7LZluJPXTPtGygpBIHa501QU2IBBMUgPiI6ffy
zloJGQnLYJuLqhtVZv7sX4KiGFnEY+fp7HVieF6XYlBsVV0uBZd2BaDkUR7+zeM6WP/gAy8NN7Wu
FdIEJ9S7w8h+lx210LKwMJ6skzIXLDTtJpjMcfhkOXKjo3FNo/IBNybXHeS0/5c9DWunlNIJQqXf
M238pZSQJrHC19pCuIIzrMmTp1+JPm+NgA3/NYX73lcBlaWfe+Rwzx/btPcbfYUlyvXOlJkeoCD6
SCTCTNOpdTynwq2oTSTtSSrGoWS+2CMnYEuTZE4QgwAaY6DB1YSOF7idYrHS1F9Mh6wfiJxTSUkQ
dtrWZzACMcDn2LAh8RXijb91VfyIcpJhJTF22ntJoOE31i0THRtlBUBT3h/HwqsiOT8p4BQZBpGe
aV1o/L3sY9cjUvzSGuYAu2P65P/uXBKUVyy6wJTKLB4R5Uy+lqi0gzgxvyfEdNcjPxRTFx9R5w4P
/jeY+8ge2T9KHuBZ6wTkgwQcw0BhU4HP0V32omK9cmC52bm9UEGhuqE86hqFeLGlafAugneCaOA3
cl8dkFjnuQZnD87/6b6mL5WEqo33Tr9lgAjF0DMQy8YdjG7PnQZK654LOgvglltZp8h+gK+/mDmA
19uzav+EaEldRN4HbzLgt8u0FJSuhyUmdjW1dgd1sXwRfcdexckhjtBe6dJph5RbyADeV0GEoH6c
BkB1olAq8FDN1nEJsopa350aKQXjdiHlgTvL1dns/Rh9pgqkj/K+2qHPJR0yzP+7ylQkVfer1EzN
RTBSdk8Ks4h9F9siqVfHLZPLsjxcbsGx1idPCKABBkxrHxidbZCV4hMncCS9p93ITPckOaPwcXAn
P2TCgZfVctdE+0+DCqZkKrKfn1IDN/B9n57wvg7Lu5sNxtkUKVbwzGmgxY6eQRcncYrXCRCN66Aa
eCg9OPp9fKiqhcAcNGDqTHQvDfcMPDkzQJwlrw/4pe83t0tW0MunQxAtrIIqfSYoVWnNtRL0gH+J
lXeYg7Ssq1fh3rPPahse4OkM47m9EoBZB7bnC6Z3teuETicKA7n7F8pgQQWXS/1fjpdzfwRv+XWd
ktrqIr1CXAbDdgVrNqHWxf/3YnX79NHuyGonaI2yGkOmcYGrx5fuxoK+/NnMyKJOerItMRs/34O2
zZ3ddpW6KZ8kWVMFv3r6IYP1s+6mrBZmLKufVHRxHFZD75OJECecblyA7UpLGJtHJqWh/LfAMvmm
90/WxdFv4gOARGcfNM3yY2LNoe6h1JvhwzV/UXzT1Jj7gGnin/5L0FFNP/QFZsxQI/7MECVpZe6X
X0WGsP8Slup/g18vZfGjs9yzOjEtEql6KTEO4yzNv6Zt6r/DfGlRahH26Z1bdNbnGnEqT8hcz5EJ
W2wfyXtGa5y3C66luDVktxPYhZMF3ZJmYdTW0CDDo7ehaacJKHD37PZ30Hb/SuT4XBQvwBHYkYjY
PgakUJUnog5RpVqP2tB+Obl25iN2WlaXUT359FHX+eJdNqJHx7TCySfFQQncDDyXc2yddeeLvnxw
huVuURGMGrnTtg20sL1gbmAQRDJZ5XhrSIYw+hAaBXv/ogcI0k+t2D28SxWoUDAM1rSX0Wa0JkZq
kvVTD6CXX8+AOUvO+X/Mng9s5Jnw3uuU5UsrAimRCM8JbUwb5rHN+vRIYOOCyNtkqWzSxKFpWz36
scryem/f9AK87O1IrpYD6U0Pt/zS9wzi8ZdxeKtB5oI3udW9OCpSKwDcWZdtQ+yCwb7g7t9nD8zs
/ytGc8VxnolbBIg/RF07qIhoIaSXhLoOnW7odOfVxm/Sqcrsrex6is0DlfAfZo6Bu0RJm/9pAZ8q
Tr0PHdTfko/Y4Ek4f2FCwt+wDVKakEmegwzLxJKWxTkAGHf8eNKunkrxDbNjlCrTkR8U9AMJXWtf
blB6NaeW/dKGYW4RUeivXxgwjsz0vf5aJnGD/zLUYin2+a0PQr+SFfTaWd6ld1PR8Vpb6GWPK1XK
7QoaXKIc+MaT1lODO57h9vwhT6c7Q8Yb8RhVISmDzDu2BM6JXTqeA/W/byWDYYGKd4eFGtEgUy9R
IVAP5nDfIm4FuwArW253pb6MKP/4LopC+78kIl/x4hqQl2G6uxCtl1Q236L8SEZAPKrG0+3M+VUM
QSTpwr83rEQ3UplM2xAJFV8AqJKu3cTxhkOijdGRHi4J1HbZKNH3yuLrLPvwDbxrvdgPVemKbaRj
sC5EjuSQxetuS18n4nIoEtpw5Cse0QdZthpByTH6R1z+x4+NAyTExqg5bMy2DQkM8loCE+HjOag8
xjFfkPnXrjf56ZDeQRcSUZ20q84zr1GfrDvTDOnUoVa0DTmqyC1sk6cpR3vfEnc7tA9p0XrqfdXz
FF8RI8msxV8D1z5MncNKlNioBHoXecF6UDuq7CNM8oaiIm7Sh2+pvs/X5ezZFJ/p9C4cx4jCm4c2
AqxalrnXMX7aU1b0voXT2YlhWa96ErY2oC7Jfmht/4nLIuN/fmtO9zDe5528OosZLaLmG0A/jd6V
KHV51fMz6usZBnOX5WqRXwfdCG4KWD1vhZv8SiIs2DY7FVZZ2b688V+ikZr66HPyHYjhyH6gHYc9
AFelFEhzTgd4c1cZ6A5gmasxJyOLvm+ObCFrJYYG09sAmxj4Hwm9NBdmCTQr9P8HxiNBdfaFCVYg
NbPD6aCo1LGf+cKo1K6RgDflTsWqLS0GXvsFr+oIpvf9O+9gmZzwSkKDzda+dWJL+XLXnZBw+OMP
13IGXvDgTuBMBQpwDBepxThGqjmEo9Y6zbBKpZn6e976scJZLa8ZSKNyhu10quCiFumTrd34u7Tv
DPIwtJyN4u3zD1hy/4APsfrCsSGAS9b1c7SZ+ukuoqv0AvtcBoK2UMY9Ci/4HWzYv4Od1JpcOXCP
nupfjj9B96RoZhf7qjGf0IaDSKHYqQtduwNXlKfOGv5u7lAuQLQ2rbblxfBad9fAVONssBuKNzqX
FM9jxyn1zPJdPVpcE9gf/cEsGrNMbjlwallgz9751oLXxxz340T7jUZX+Oejsy/VViF0C8b0hG7Q
pEzb3eTnn2RbgP6ZQQVE41zPlu8DU+eVP9tYNY3Xmg5Rpj4f1mi0csIYw34PwEabjgQkJDy0bjC0
EuQDRVuu0sDSwMFPTucreB2dpBtSHJrGQRpDdK3W8hj7dVpglk5GCrv+Jwp7c5yvf0tIfwL6Mthx
Vq4PMkebz38sy7pGgv7GpNulJZxYzBkkeAbIxlyOgxgkSy4/Oe89uyLBQR3tpp/678OeV8EtgPBn
yjS6XMXx1I8e17Ywxhi7czRVqnZJZ73tTjWWenbM9qH7CrYR4FiaohtOTI2LXditF8nW6SHSL2JC
w1o2laOomTphD18fW4yAz5rDxzkduYlFaaQKyFzxQccgR/52BJGxWXBbtgARVZzLnubhbHk+ixwN
YPywxdlRPvkMKSDHgWNKK2TjF/nH8Oiwu7KYsXDsHXGcQBtWWLmNSAc9Oi8DpcJGMXZ1ncrv98sD
gLRnVrUJd4VDo68pefVJbiSACKJ1BWvn4M6Oy1JpYAFdH4DLk7o5xFfLaNoN82py6Ca8BBgrR7OJ
9ibg0Pjh7i21Dko7Nwy7eRut7eG0ZQBfU3Zij1QNt/b6xIPJUFwGoQc89sdIEoKFBEDbk4cshFDI
9EuZ3QnJ+gsAtbG4LocODaHhTi8c5x0Oiz9Qy3eNzEjccXaVZgiPayvcoKmwdod7fRc2BFnivSeB
kb0zi0xw/5ljjRJTTPi7zirbUkt2FU6BUIOQXE7Cncs8DzjdxRNs6TkP/quqKvzy0VYs6RAyldd8
8pfRCMaH/+uvVQJ0NZQV5Yw+fiVyg783rj6Je2bbbFvfJyXVW6ltd6+/CBGgR6qlIQYCD7PBzpib
Ts6dlBSlmO1CfmZGM6F+oACszCRyD3X4g4LqP0n6ly0x4+XZnHW2/6EpamDBS1mHtfJ73lJbF013
xCn7FQiOvrpKDnpNb0zZp2yWGjxIFprZvfM2rmcYgPmmIWSCph0Vu4Kvsg4ToJcEmVIIeMjBuo0u
rFqKWTvO6MvTxD5ynd8h4Pb3YGllXyb6iVTPJLUHYGDPHN0fgjfS5U5EQKVU6QR8NxV2wwBzldAp
uPo8pxjMLkEC9PqBl8wII4ea1f6xXhrzZZzK6LfBPLf5FpparW8pAS2uvFbag2egQRiwwd+svtJE
m7X8O1c72RzQvj/tUq99WjpTAa+evmfV5mqFNDInQKK0DJ6T4R/Ueiv7YYwm0MOc6xFEz0c2FeCH
lCFoVNtBSocqzDIziOyBqVYgBYRa0wQERqvJlEifAIEJR8gFQcGS4z783HXpki3P0KE3ZqlNYBf9
JWEdCCsi07999nb1W1SZ1aJTXb9zrDmGp7Qf75vgd5rZhcLc+7ivKNoEDUzUJF953TRSJdDoqFqb
jGPvLJ866f89tQ+TF1o3TF0+0RVL7UPw85h5d6VKeAni5B6O1b8eVRHiGyDGYzcAXqdesVyYLXpC
7pxToo+5277JlLnIobPgLb2yuo5UfgsTD4iB3iN61cM2c6jW1Hatv41E1RY67+Uu3bj4OwzaJweg
iuIzZe/S2A6r2RMnp6lHTesrcPy7aip6MeiWGY5nD1Le4kTrdGhI9VG65IbHvFWEy28jzW764fuN
rE2QOClKRmeaNPdm8kTQEMAYzQ0WWbx4vmtuCZNiXOpzZzjpML/pdZH5PJU8ma06Vv7A3z2LJwn3
PmmqOReirR5470yQpNFhGAvrWkGugNYjlrjc6usZJ25wOHi53KQg/6GxopUGt/zVdVioVp4XJ3M5
gqj+cczEO/XnT84B/3X4itwHWswb5CLWHfui34ttKcgv37bt2MG+27sq403aCmxfBjbJpWq7Xuyp
X5JLoQfjoQfhM8TeaYhHIz6nirAdrTOsLKQcHhDtTC6o7iV8C9fErSJpgJrpiI16u2/VgenhybLz
bTSnBRXOZb3rVQ9VOTeRF3gUVUgNUXcPNFkLo4HI69lopfBVpSPZTi3/7s9dOth3DQaNkNL4Ev6u
3JSblLZwWy6hmRPcqCib63ZasLnmP8UIF17RgksxAPysV6UOfpr7Ilz0Dju4goMshueQd47mGFxL
RWwJXMp8FJ3UkGqWusaHoy9B7AuYxJl85f81zEzx89XOLdgKedIsA9WMvF6TobQP+U+EGOEYiJhO
3Nhs16pSIW0A/HyhzLi4TWyH9KjJeq5Ya+w2xkY/niYdcSHkwhtQtp4BLf6HtFj60rNZbzSzk0uk
8UrEGLmydPz6pN+O1ttvXFT88sfJnCSLfmSsSlHRVw+JL6p/nw+1MagkqAjaTymIBuHYBLT6OgCg
jMhVqE+Y9Ka6OfbQXolv0AaBCxtQzlndaYeKeCZtpfUOoXB9nEE038PPc2Pq3PdWBLe3edzaM4ZK
rNnqJKjbvYmzqsmlKOtzUnst8iSIvAmRkUJQwC+sT6eAG9SbVyWGcmH5iowewxliHcQlHNQZIRxn
gs1t6bAvNr37h9UdH4cmPpmU3qOScXx7mL72ZkSo10M2lAA/jMNDCX4q9kFOxSvsFYmz9RGYDoPi
D+oJOjJGeWyuvhwO9yEKATslZjHUK9Y2NHUHfzieAJ7SJRERDfG+9tfZZ0db77Zrhj7Aod7xkzGg
XGQvrS1LEEql6xbfg9NENuQ/8SufFJXsozCFxjkR81f3dm0xY4IDA4mfhSmfN9Hey9SnwBPc9/rS
zJpZuDFpw4iIwq8yBGu1g7NEX3uQxCKaAsbJVRqVfHv79sBqyhursT1Ap0ee8uXOw6kOyAurFVWD
r9NyNEAx1Pe92oAwEbD88AXAMxoTlubR/dXivwagxcjXuxtUrGXEJ37ky65BRNh8A5oN5jsZf9ag
Q9sniq/n1Jkoi3xUDK4rzWYU1oGHQ1EbauhHNLYTumlG/BOyHRzH9ZE0/EnMI0cwpvDaGDvomD1p
gjcHv6usAZ1RDnreebKnR43vnm4/EqHT2KWId0aSjCumex0SPZmgP9Tc7Q1ZSZ+ec42W0+hkSYX2
zCVk/iZeYZpUQAunbctB4L80R9mnjdwNasHRnxDidVowSZQXDMs+5IiXjgxDTAyI87RxOIs1XzaO
eO+lHKgwgOB+TtBkDoAwfX8TQtF75I6scQDoOZkPVZ1i+8wpHbjsgxkSLATRtQEY0k5MyNkTEljn
EtcpFMDk2Ps8Hiqih8yYEEqcth0vZtibgl8Uz/+JoZ4oyNuxixH1znhDnD1wo2W9TDq4yJZqK2Xy
PoTYHoL7jgsdgfxgFkRA2Jy5rd9Tkbnv8s11TjTHL0FS/cNYEjBrve4L/6hKufHv9NIVxYLLM4Zr
e9kkQUx/vDcsvPe2SzhEhR57eWEfVG5wmTb3UnVwsUrh2pMl7BMSrWf2Anv6mtvg7u3CatnAsm7i
khkunGx67OjzSAzRruaZVgpq9WKI6sXJQWRDRT6MuiURcHgS7ctgxIoLD28gWmd+7KYtbKiISC68
N0JbvCwXo4oSVHXU4wB2trUbFFoS8hQhXcBqWDUp8wuTQhSoVbTyEBKGgQVtyjWgqq2dH/2Eua3m
MnbMl0uZAzlqI8P4t+AsSOoSMZy8lSJ8W/G0PL0U6ZK3MoRHAlOTW6/D3wVJIEDbnipIwEyuKjZm
zEXokY4ZE/dXIkm8uPVGcDNHNUBfPIhuuhteK5itHYSGcxnfjEdVsVnAfotjnGmBOgQo6V4l6RnE
Tpr6nSedmKRikrmR4BrXW71jOxS7o68KPLPdWcVnOb3ofWo4nMEt/DHHninDKg6tIgbv1F82vIe1
2C/8K0NVi8Cd10Dd886rMhY7vlnrYshj7P1MbXuowUo8+M5iMVFuawIk/m5Q3sPYlSK7cIaidoMn
Yvh1STsxpDNzFc3rgrHmNmv5xMz/Hmks+E75J3tyVH1sZyUs8/9a5hp+N6COo8TQ0JciniKukNbJ
NbzoxMP5tCvAvhoq7VZ4ATQHQrtSUmIGBIki74U5rBDCZ8+mClZz61h0fTu8mbLD3HyCk3EKM4j/
vhURgYNJI0XsbOoOGU5Fn96Crl4qi89VeG2DcFc0G16XgZ+U8L6vx+x5UE7UpY7OwcfQHsdlNJLW
6OIQQIZt25SbdKc6NSq049CX54iH9nC6p4BjUgG8kmWwfNVf36Jvi/TNtykCXNgPnEUzym1Kwa3e
hk952YXSdBB7BKhibzCQ1NwUk+l5yTEjkZ5r9SVF/4eMHvCTlarySGcL70xOQ0HpYLISFmq68PRm
FnN9jrueO/haC7b8Orry8Gv3fMgNwz5sUMqI7yq2Pr3ZWCqZg6pnBTctmAIGcARCy6O41UOJYVVu
v/8awA9m9Tzn512IeC8u8AB5tA9BpipGVzagTIBbzNjSdC/2cCitPJ3JjSPK/GufHap7e+E4yoZ8
SrmfAxTCkNVWytb+pSTOvj+FuaEeTJSNQwr3xXnwHFMxTXTNtnQl4XKKFa2PXRiAecy8v4sYXEpX
cwv2INqQ8KTRa00PPxVyMFq46vMoi0/ue02ycXYc3hgKlZT13awQho7whfmpsjK0Uh2dx3hXK14z
2r+kooyljEZ/1u7npPt+AQ5EwsmlAsbD6zAxCUYU//4EoUZFkMcgyYsXRzWRLVxcHYe9kck0kqy3
Z3PShgvZiQd72/y8sG/P8dZ4jGdKdvhKhLkbUi4Szn6BsWRLdIJkPWMrWUDBPLoF4a/Fky3eBD8W
gEF2Vjid9AicaViWGYI7Gk5teiJIr0/8NXe4bf7h0qEwIf/oD3/R5nR2CHWkKPaajZY65Vtvdl+f
k2GDuakYfYV0lLf2je2W0h9xna1nRKbNJqVd5/euDKivGopY07i8Y3CrwxMMnHTmUcCpOQjpzx4X
T+cdGczy6TbPemXGuC+L7WcohpEaukKSmVi+8kVsnnT9FANMEq585XVWD6De5/lBRXIVkS4yZCBu
feSqeRJl4BO+GcCV3HB9EN+8DP9Lm88lJhMIGqZJySZIj1QsYZNjBM4tNrXVRO2ZQzL6rTeOrsBr
RCCKLdxBxkQyq2N5DbjRe1Cy6XqIN2XfUSAdVV3oP/Sx2mPmRknCM3lDg2BHH5XBa4HgR2GZUXBc
Evqq/KDoUqpNbJ3H8nf68PoeDlTsOYssQQcmt/vlM6FW11dl8A5iDsBXNvr8JVXlqQ1XvF0IQEm3
cKBHyZ0xDX6hnvNgtLPheTfkQsLG2U/i9N/4nyGwpqTHtHGzbjvqbfKHiI0QGNf0cBAVHhBnarOu
M9EVFA5bdM+x8cmszSnaSR2JpiUNgTvzIaTIq8iaMZIdPB+hzCGIVLeSvcN9S83kFD/faKfsRWdS
1pf5sGv1F4w4NO4erKdlMdxJcY2PYOZGN+88TmrO4EjjPMXDvlyzyd9J/cC+JBW50vnE+nP1VtZT
rcvoctIk+/N7UISDxgWi73StZ7ws4V9ZFCFpaw3qBzdk1Q8H5rnNS6eHF4dgEArmp75wG7b2JkzR
TqI3fCFd9cEY1/orMD/M3qE0L55c/J+ofvYv4nAbrPwvtQb4hd6hXUiJNZTkapuVLXcdjeqhvTOT
9b0PQ4LRqt9gcpFe9kgCyVvZQbc6ivv4IxzSiaSo1apb/UFGqrb+pVLxYrBFqQ0FatUbQIMb4twR
YNfhsF2RS9y/K0h8z0+ht1B78zueGF7PuP/X9Gf0zD8gMPZGu1jCLQElCMHvXZz8maFMo4F9Qequ
0gD2QglVOpcpfgNzY31FYTTnQz6cnVfrFXWLWirqK6H8Gp+SGEusXd2zPK/9aamhbiDA5T4dRBP4
Y5tdr9+UCXOogPPiaUWRSveCI5loUn7RAQNeDl/44m9rIqyi01rnqyjlP4Ud5YuJGjl1jOW7Q9Ek
dq4pSdOeZsz0MfG0W96rNtFyqaDQCvfObl5O3c+sBseFLwG0+73KJYoDJHr0iNlk39WvBWF7541j
H7Z+Unyg3QQgMLdQivI+W+D7IaFiIav+nc/B9vVdl0Wy+w4dgYMfJq4o/5FlhBzwPm3J4eAgUagj
a9wK4sbQpP4xJ7WE2aEzCkOt0RhqvvodUSfBv3Cpz8O2KMdgpmaV9huGf7GqTh8XsaVT1aTrza1c
iwhzuE2+2tUG6zDaC0xuG7ihrfa9YT5Xj2LfVizhJFaWmmlcqX79bCwUbfCvuQ23L9rSz275lwvl
/48si84erBCl0KHUQXjSTdvVY6/ku7bWLxulb9WlhcigTDelIgCfNi0T1b7k+cpXuvSUTJdFrJvW
pJ4NXmRTMgMoPayYM0HKsPINm4AS7fFsr76yWiN5oeSjt7/D5M1/YSZnKeDFjtXs5J0m7DpoMh+o
Jt3YuQqezJtZIQSB6T+jsBmpP+45ZYDk3BbXXQZ8KBCtPjDaSpKuiOWXV9f6N0li1kxrWxkkliqx
FaoehP0uMJ1cu7m+bWMHqHP71R+N49f+dcdyjNUbYpEyafA/klk1qt2xJiC8/374SapLGkgeN2x6
6cOilfp+HP5zv2CSuIK/+VGLu3aDknYWZ8SsH4WSrP0VSJxZRq/ODyNd52niX0eGlhXWy4zGuTtc
oEmeVbagS1UTNLIBR/1vBUyMh6s2Q3ttd4re0ibhWrXjz1uOdyZ5cZsGi329ouDNpdXlzd95b5WV
LzjJi14XdTZuRgEiF9WGBjFV4/bzKA9S840eZEalOPjXMZZ6OgmFvJm6qWUT3K+MtFW0TqIdWIH7
XU5C/F0RCe6cvmreU47z1hhVmZXCsDBRXYIwvpvXr/5WDkmjRZLZ/eHfcNK5Yan6SACgAWxT0FRl
PAYd9iHrKIMj8jnW5t5WsWmuO/Ob44s8GedxfEjwhkYn96V0yx7Xd3cQ+NkMG+kJJgyKZNaW6L22
Y8PJRN/DGtfI2iQq3c/uFo48hRRT7GgaLNmpCmJ+eCKjf1MfcEtjdI0bohBvzgyAss5W2WPDVO+S
OnHmMNPD9zW8h+lhdZeEfFOf7Jq6VAoAHHmTBXWzZtyBZplvxiGd9HmQKIbtdw2pEB6nBmzydYz2
uwtk14jieckKh61QTQh0qqTFs6kDW9X0npAqld1j7HkDYI4b7EZnZX0oKlHAVx9nMhM4f3Polnj9
7LQf8SjWDxoF5OA24ItW75Sa6303aP+wPszFl28Zwz9w4MbEAK2MmnXD2kPwt6haoAyCBJbTOfvT
Qc0BZTUC0mDboPjqDT37EMDgNeP7eH2bkyZLSfSpFSRpKdN3mYg+bnL45mUQGK1klq26x9tp/sYo
qWjkndFrz2JrKl03Gsz+nvoXk9hgKykXLXWkUohtfevVyYe6yI1VcZQuBJN5Nzoo9lP8wfj2UkIU
QJBN0A8P8vXxkDAWxVw+XNR97A8336QvnywG842GTiy+U3DDXVM7X/hKcMQf9KtXJrK1fda8do/P
v+xIAmImKcDFXcZvZfKywuVznwfz1/lSY0FoLmsI2nJijgghm/kxgaVkgB2BGXjr7veGszO3iLDz
dWgYvB34GNKw6ZAS4wuHVZYNbVq4C3Pt3PXK6R7DMQJMCZutuWcQfkl9Ii7Kgs1GVgUT+zbQS7W0
JHmY5B+0fAZjekyuYiJMRdAZztnrYGtUdwN0HvGimM5Ep0tBc58mKWgIM9DUcX0WKDA2Rhm0WXYr
Rix1cz5EkWfvNuEvWnJ8UnSaYsU+QIIHfaDBfA1s21GeyXEshgVEbkJFb0+blu52qrrp4nhvCTtv
mZ7akWH9hSSxH2xJl6pbeUloX5xTyuaImqkVlaE+te3Eat57NEkCOpOmHpdIFl51wCP6xa3+HwVb
1RQrqaqtH49tNdkInfsAjs3btmcZUQSyg55TS90VV78NT9ZKj+AEQa8k+Nq51kY7+wvUhiQpOXea
c9ZtdmURIrPpJMV3RvUeld+ytRdmwp7XpnUf0jyW35Hbwz6sthRElwtgBT3UypGIobOPe5mfcQVf
vgrnPkwqEhKan4jlU6lMFZZof5FHufAcRjNvaGOmxBldudTksRWZM+IQQuGrunKD3fRTCRMovRKT
+F5eTOTvhTB1eoSzn4DNkC5v9IBpvKzVK28IaX/8v7tRL4m2GFaMu82UmpLbWxdpgVDD9T0=
`protect end_protected

